module pebbles_core
  (input wire clock,
   input wire reset,
   input wire [0:0] out_consume_en,
   input wire [7:0] in0_peek,
   input wire [0:0] in0_canPeek,
   output wire [0:0] in0_consume_en,
   output wire [0:0] out_canPeek,
   output wire [7:0] out_peek);
  // Declarations
  //////////////////////////////////////////////////////////////////////////////
  wire [0:0] v_1;
  wire [0:0] v_2;
  wire [0:0] v_3;
  wire [0:0] v_4;
  wire [0:0] v_5;
  wire [0:0] v_6;
  function [0:0] mux_6(input [0:0] sel);
    case (sel) 0: mux_6 = 1'h0; 1: mux_6 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7;
  reg [0:0] v_8 = 1'h0;
  wire [0:0] v_9;
  wire [0:0] v_10;
  wire [0:0] v_11;
  wire [0:0] v_12;
  reg [0:0] v_13 = 1'h0;
  wire [0:0] v_14;
  wire [0:0] v_15;
  wire [0:0] v_16;
  wire [0:0] v_17;
  wire [0:0] v_18;
  wire [0:0] v_19;
  function [0:0] mux_19(input [0:0] sel);
    case (sel) 0: mux_19 = 1'h0; 1: mux_19 = v_20;
    endcase
  endfunction
  wire [0:0] v_20;
  reg [0:0] v_21 = 1'h0;
  reg [0:0] v_22 = 1'h0;
  wire [0:0] v_23;
  wire [0:0] v_24;
  function [0:0] mux_24(input [0:0] sel);
    case (sel) 0: mux_24 = 1'h0; 1: mux_24 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_25;
  wire [0:0] v_26;
  wire [0:0] v_27;
  reg [0:0] v_28 = 1'h0;
  reg [0:0] v_29 = 1'h0;
  wire [0:0] v_30;
  wire [0:0] v_31;
  wire [0:0] v_32;
  wire [0:0] v_33;
  wire [0:0] v_34;
  wire [0:0] act_35;
  wire [0:0] v_36;
  wire [0:0] v_37;
  wire [0:0] v_38;
  reg [0:0] v_39 = 1'h0;
  wire [0:0] v_40;
  wire [0:0] v_41;
  wire [0:0] v_42;
  wire [0:0] v_43;
  wire [0:0] v_44;
  wire [0:0] v_45;
  wire [0:0] v_46;
  wire [0:0] v_47;
  wire [0:0] v_48;
  wire [0:0] v_49;
  wire [0:0] v_50;
  reg [31:0] v_51 = 32'h0;
  wire [31:0] v_52;
  wire [8:0] v_53;
  wire [8:0] v_54;
  function [8:0] mux_54(input [0:0] sel);
    case (sel) 0: mux_54 = 9'h0; 1: mux_54 = v_55;
    endcase
  endfunction
  wire [8:0] v_55;
  wire [29:0] v_56;
  wire [31:0] v_57;
  function [31:0] mux_57(input [0:0] sel);
    case (sel) 0: mux_57 = v_58; 1: mux_57 = v_62;
    endcase
  endfunction
  wire [31:0] v_58;
  reg [31:0] v_59 = 32'hfffffffc;
  wire [0:0] v_60;
  wire [0:0] v_61;
  wire [31:0] v_62;
  wire [31:0] v_63;
  wire [31:0] v_64;
  function [31:0] mux_64(input [0:0] sel);
    case (sel) 0: mux_64 = 32'h0; 1: mux_64 = v_2542;
    endcase
  endfunction
  wire [0:0] v_65;
  wire [0:0] v_66;
  wire [0:0] v_67;
  wire [0:0] v_68;
  wire [0:0] v_69;
  reg [0:0] v_70 = 1'h0;
  wire [0:0] v_71;
  wire [0:0] v_72;
  wire [0:0] v_73;
  wire [0:0] v_74;
  wire [0:0] v_75;
  wire [0:0] v_76;
  wire [0:0] v_77;
  wire [0:0] v_78;
  wire [0:0] v_79;
  wire [0:0] v_80;
  wire [0:0] v_81;
  wire [0:0] v_82;
  wire [0:0] v_83;
  wire [0:0] v_84;
  wire [0:0] v_85;
  wire [0:0] v_86;
  wire [0:0] v_87;
  wire [0:0] v_88;
  wire [0:0] v_89;
  wire [0:0] v_90;
  reg [31:0] v_91 = 32'h0;
  wire [0:0] v_92;
  wire [0:0] v_93;
  wire [31:0] v_94;
  function [31:0] mux_94(input [0:0] sel);
    case (sel) 0: mux_94 = v_2437; 1: mux_94 = v_390;
    endcase
  endfunction
  wire [0:0] v_95;
  wire [0:0] act_96;
  wire [0:0] v_97;
  wire [0:0] v_98;
  wire [0:0] v_99;
  wire [0:0] v_100;
  wire [0:0] v_101;
  wire [4:0] v_102;
  wire [0:0] v_103;
  reg [31:0] v_104 = 32'h0;
  wire [3:0] v_105;
  wire [0:0] v_106;
  wire [2:0] v_107;
  wire [0:0] v_108;
  wire [1:0] v_109;
  wire [0:0] v_110;
  wire [0:0] v_111;
  wire [0:0] v_112;
  wire [0:0] v_113;
  wire [11:0] v_114;
  reg [31:0] v_115 = 32'h0;
  wire [31:0] v_116;
  function [31:0] mux_116(input [0:0] sel);
    case (sel) 0: mux_116 = v_257; 1: mux_116 = v_1374;
    endcase
  endfunction
  wire [0:0] v_117;
  wire [0:0] v_118;
  wire [0:0] v_119;
  wire [0:0] v_120;
  wire [0:0] v_121;
  wire [0:0] v_122;
  wire [0:0] v_123;
  wire [0:0] v_124;
  wire [0:0] v_125;
  wire [0:0] v_126;
  wire [0:0] v_127;
  wire [0:0] v_128;
  wire [0:0] v_129;
  wire [0:0] v_130;
  wire [0:0] v_131;
  wire [0:0] v_132;
  wire [0:0] v_133;
  wire [0:0] v_134;
  wire [0:0] v_135;
  wire [0:0] v_136;
  wire [0:0] v_137;
  wire [0:0] v_138;
  wire [0:0] v_139;
  wire [0:0] v_140;
  wire [0:0] v_141;
  wire [0:0] v_142;
  wire [0:0] v_143;
  wire [0:0] v_144;
  wire [0:0] v_145;
  wire [0:0] v_146;
  wire [0:0] v_147;
  wire [0:0] v_148;
  wire [0:0] v_149;
  wire [0:0] v_150;
  wire [0:0] v_151;
  wire [0:0] v_152;
  wire [0:0] v_153;
  wire [0:0] v_154;
  wire [0:0] v_155;
  wire [0:0] v_156;
  wire [0:0] v_157;
  wire [0:0] v_158;
  wire [0:0] v_159;
  wire [0:0] v_160;
  wire [0:0] v_161;
  wire [0:0] v_162;
  wire [0:0] v_163;
  wire [0:0] v_164;
  wire [0:0] v_165;
  wire [0:0] v_166;
  wire [0:0] v_167;
  wire [0:0] v_168;
  wire [0:0] v_169;
  wire [0:0] v_170;
  wire [0:0] v_171;
  wire [0:0] v_172;
  wire [0:0] v_173;
  wire [0:0] v_174;
  wire [0:0] v_175;
  wire [0:0] v_176;
  wire [0:0] v_177;
  wire [0:0] v_178;
  wire [0:0] v_179;
  wire [0:0] v_180;
  wire [0:0] v_181;
  wire [0:0] v_182;
  wire [0:0] v_183;
  wire [0:0] v_184;
  wire [0:0] v_185;
  wire [0:0] v_186;
  wire [0:0] v_187;
  wire [0:0] v_188;
  wire [0:0] v_189;
  wire [0:0] v_190;
  wire [0:0] v_191;
  wire [0:0] v_192;
  wire [0:0] v_193;
  wire [0:0] v_194;
  wire [0:0] v_195;
  wire [0:0] v_196;
  wire [0:0] v_197;
  wire [0:0] v_198;
  wire [0:0] v_199;
  wire [0:0] v_200;
  wire [0:0] v_201;
  wire [0:0] v_202;
  wire [0:0] v_203;
  wire [0:0] v_204;
  wire [0:0] v_205;
  wire [0:0] v_206;
  wire [0:0] v_207;
  wire [0:0] v_208;
  wire [0:0] v_209;
  wire [0:0] v_210;
  wire [0:0] v_211;
  wire [0:0] v_212;
  wire [0:0] v_213;
  wire [0:0] v_214;
  wire [0:0] v_215;
  wire [0:0] v_216;
  wire [0:0] v_217;
  wire [0:0] v_218;
  wire [0:0] v_219;
  wire [0:0] v_220;
  wire [0:0] v_221;
  wire [0:0] v_222;
  wire [0:0] v_223;
  wire [0:0] v_224;
  wire [0:0] v_225;
  wire [0:0] v_226;
  wire [0:0] v_227;
  wire [0:0] v_228;
  wire [0:0] v_229;
  wire [0:0] v_230;
  wire [0:0] v_231;
  wire [0:0] v_232;
  wire [0:0] v_233;
  wire [0:0] v_234;
  wire [0:0] v_235;
  wire [0:0] v_236;
  wire [0:0] v_237;
  wire [0:0] v_238;
  wire [0:0] v_239;
  wire [0:0] v_240;
  wire [0:0] v_241;
  wire [0:0] v_242;
  wire [0:0] v_243;
  wire [0:0] v_244;
  wire [0:0] v_245;
  wire [0:0] v_246;
  wire [0:0] v_247;
  wire [0:0] v_248;
  wire [0:0] v_249;
  wire [0:0] v_250;
  wire [0:0] v_251;
  wire [0:0] v_252;
  wire [0:0] v_253;
  wire [0:0] v_254;
  wire [0:0] v_255;
  wire [0:0] v_256;
  wire [31:0] v_257;
  function [31:0] mux_257(input [0:0] sel);
    case (sel) 0: mux_257 = v_278; 1: mux_257 = v_390;
    endcase
  endfunction
  wire [0:0] v_258;
  wire [0:0] v_259;
  wire [4:0] v_260;
  wire [0:0] v_261;
  wire [3:0] v_262;
  wire [0:0] v_263;
  wire [2:0] v_264;
  wire [0:0] v_265;
  wire [1:0] v_266;
  wire [0:0] v_267;
  wire [0:0] v_268;
  wire [4:0] v_269;
  wire [0:0] v_270;
  wire [3:0] v_271;
  wire [0:0] v_272;
  wire [2:0] v_273;
  wire [0:0] v_274;
  wire [1:0] v_275;
  wire [0:0] v_276;
  wire [0:0] v_277;
  wire [31:0] v_278;
  function [31:0] mux_278(input [0:0] sel);
    case (sel) 0: mux_278 = v_328; 1: mux_278 = v_384;
    endcase
  endfunction
  wire [0:0] v_279;
  wire [0:0] act_280;
  wire [0:0] v_281;
  wire [0:0] v_282;
  wire [0:0] v_283;
  wire [0:0] act_284;
  wire [0:0] v_285;
  wire [4:0] v_286;
  wire [0:0] v_287;
  reg [31:0] v_288 = 32'h0;
  wire [0:0] v_289;
  reg [0:0] v_290 = 1'h0;
  wire [0:0] v_291;
  wire [0:0] v_292;
  wire [0:0] v_293;
  wire [0:0] v_294;
  wire [0:0] v_295;
  wire [0:0] v_296;
  function [0:0] mux_296(input [0:0] sel);
    case (sel) 0: mux_296 = 1'h0; 1: mux_296 = v_297;
    endcase
  endfunction
  wire [0:0] v_297;
  wire [0:0] v_298;
  wire [0:0] v_299;
  function [0:0] mux_299(input [0:0] sel);
    case (sel) 0: mux_299 = 1'h0; 1: mux_299 = 1'h0;
    endcase
  endfunction
  wire [3:0] v_300;
  wire [0:0] v_301;
  wire [2:0] v_302;
  wire [0:0] v_303;
  wire [1:0] v_304;
  wire [0:0] v_305;
  wire [0:0] v_306;
  reg [0:0] v_307 = 1'h0;
  wire [0:0] v_308;
  wire [0:0] v_309;
  wire [4:0] v_310;
  wire [0:0] v_311;
  wire [3:0] v_312;
  wire [0:0] v_313;
  wire [2:0] v_314;
  wire [0:0] v_315;
  wire [1:0] v_316;
  wire [0:0] v_317;
  wire [0:0] v_318;
  wire [4:0] v_319;
  wire [0:0] v_320;
  wire [3:0] v_321;
  wire [0:0] v_322;
  wire [2:0] v_323;
  wire [0:0] v_324;
  wire [1:0] v_325;
  wire [0:0] v_326;
  wire [0:0] v_327;
  wire [31:0] v_328;
  function [31:0] mux_328(input [0:0] sel);
    case (sel) 0: mux_328 = v_373; 1: mux_328 = v_1369;
    endcase
  endfunction
  wire [0:0] v_329;
  wire [0:0] v_330;
  reg [0:0] v_331 = 1'h0;
  reg [0:0] v_332 = 1'h0;
  wire [0:0] act_333;
  wire [0:0] v_334;
  reg [4:0] v_335 = 5'h0;
  wire [4:0] v_336;
  wire [4:0] v_337;
  function [4:0] mux_337(input [0:0] sel);
    case (sel) 0: mux_337 = 5'h0; 1: mux_337 = v_338;
    endcase
  endfunction
  wire [4:0] v_338;
  function [4:0] mux_338(input [0:0] sel);
    case (sel) 0: mux_338 = v_339; 1: mux_338 = v_348;
    endcase
  endfunction
  wire [4:0] v_339;
  wire [0:0] v_340;
  wire [3:0] v_341;
  wire [0:0] v_342;
  wire [2:0] v_343;
  wire [0:0] v_344;
  wire [1:0] v_345;
  wire [0:0] v_346;
  wire [0:0] v_347;
  wire [4:0] v_348;
  wire [0:0] v_349;
  wire [3:0] v_350;
  wire [0:0] v_351;
  wire [2:0] v_352;
  wire [0:0] v_353;
  wire [1:0] v_354;
  wire [0:0] v_355;
  wire [0:0] v_356;
  wire [4:0] v_357;
  function [4:0] mux_357(input [0:0] sel);
    case (sel) 0: mux_357 = 5'h0; 1: mux_357 = 5'bxxxxx;
    endcase
  endfunction
  wire [0:0] v_358;
  reg [4:0] v_359 = 5'h0;
  wire [4:0] v_360;
  wire [4:0] v_361;
  function [4:0] mux_361(input [0:0] sel);
    case (sel) 0: mux_361 = 5'h0; 1: mux_361 = v_362;
    endcase
  endfunction
  wire [4:0] v_362;
  wire [0:0] v_363;
  wire [3:0] v_364;
  wire [0:0] v_365;
  wire [2:0] v_366;
  wire [0:0] v_367;
  wire [1:0] v_368;
  wire [0:0] v_369;
  wire [0:0] v_370;
  wire [4:0] v_371;
  function [4:0] mux_371(input [0:0] sel);
    case (sel) 0: mux_371 = 5'h0; 1: mux_371 = 5'bxxxxx;
    endcase
  endfunction
  wire [0:0] v_372;
  wire [31:0] v_373;
  wire [4:0] v_374;
  wire [4:0] v_375;
  function [4:0] mux_375(input [0:0] sel);
    case (sel) 0: mux_375 = 5'h0; 1: mux_375 = v_338;
    endcase
  endfunction
  wire [4:0] v_376;
  function [4:0] mux_376(input [0:0] sel);
    case (sel) 0: mux_376 = 5'h0; 1: mux_376 = 5'bxxxxx;
    endcase
  endfunction
  wire [0:0] v_377;
  wire [4:0] v_378;
  wire [4:0] v_379;
  function [4:0] mux_379(input [0:0] sel);
    case (sel) 0: mux_379 = 5'h0; 1: mux_379 = v_362;
    endcase
  endfunction
  wire [4:0] v_380;
  function [4:0] mux_380(input [0:0] sel);
    case (sel) 0: mux_380 = 5'h0; 1: mux_380 = 5'bxxxxx;
    endcase
  endfunction
  wire [0:0] v_381;
  wire [31:0] v_382;
  wire [31:0] v_383;
  function [31:0] mux_383(input [0:0] sel);
    case (sel) 0: mux_383 = 32'h0; 1: mux_383 = v_384;
    endcase
  endfunction
  wire [31:0] v_384;
  wire [31:0] v_385;
  function [31:0] mux_385(input [0:0] sel);
    case (sel)
      0: mux_385 = 32'h0;
      1: mux_385 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_386;
  wire [31:0] v_387;
  wire [31:0] v_388;
  function [31:0] mux_388(input [0:0] sel);
    case (sel) 0: mux_388 = 32'h0; 1: mux_388 = v_389;
    endcase
  endfunction
  reg [31:0] v_389 = 32'h0;
  wire [31:0] v_390;
  wire [31:0] v_391;
  wire [31:0] v_392;
  wire [31:0] v_393;
  wire [31:0] v_394;
  function [31:0] mux_394(input [0:0] sel);
    case (sel) 0: mux_394 = 32'h0; 1: mux_394 = v_677;
    endcase
  endfunction
  wire [0:0] v_395;
  wire [0:0] v_396;
  wire [4:0] v_397;
  wire [0:0] v_398;
  wire [3:0] v_399;
  wire [0:0] v_400;
  wire [2:0] v_401;
  wire [0:0] v_402;
  wire [1:0] v_403;
  wire [0:0] v_404;
  wire [0:0] v_405;
  wire [0:0] v_406;
  wire [0:0] v_407;
  wire [0:0] v_408;
  wire [0:0] v_409;
  reg [0:0] v_410 = 1'h0;
  wire [0:0] v_411;
  wire [0:0] v_412;
  reg [0:0] v_413 = 1'h0;
  wire [0:0] v_414;
  wire [0:0] v_415;
  wire [0:0] v_416;
  function [0:0] mux_416(input [0:0] sel);
    case (sel) 0: mux_416 = 1'h0; 1: mux_416 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_417;
  wire [0:0] v_418;
  wire [0:0] v_419;
  reg [0:0] v_420 = 1'h0;
  wire [0:0] v_421;
  wire [0:0] v_422;
  wire [0:0] v_423;
  wire [0:0] v_424;
  wire [0:0] v_425;
  reg [0:0] v_426 = 1'h0;
  wire [0:0] v_427;
  wire [0:0] v_428;
  wire [0:0] v_429;
  wire [0:0] v_430;
  wire [0:0] v_431;
  function [0:0] mux_431(input [0:0] sel);
    case (sel) 0: mux_431 = 1'h0; 1: mux_431 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_432;
  wire [0:0] v_433;
  function [0:0] mux_433(input [0:0] sel);
    case (sel) 0: mux_433 = 1'h0; 1: mux_433 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_434;
  wire [0:0] v_435;
  wire [0:0] act_436;
  wire [0:0] v_437;
  wire [0:0] v_438;
  reg [0:0] v_439 = 1'h0;
  wire [0:0] v_440;
  reg [0:0] v_441 = 1'h0;
  wire [0:0] v_442;
  wire [0:0] v_443;
  wire [0:0] v_444;
  wire [32:0] v_445;
  wire [38:0] v_446;
  wire [77:0] v_447;
  wire [38:0] v_448;
  wire [5:0] v_449;
  wire [38:0] v_450;
  wire [77:0] v_451;
  wire [77:0] v_452;
  wire [38:0] v_453;
  wire [5:0] v_454;
  wire [38:0] v_455;
  wire [77:0] v_456;
  function [77:0] mux_456(input [0:0] sel);
    case (sel) 0: mux_456 = v_457; 1: mux_456 = v_475;
    endcase
  endfunction
  wire [77:0] v_457;
  wire [38:0] v_458;
  wire [5:0] v_459;
  wire [38:0] v_460;
  wire [32:0] v_461;
  wire [0:0] v_462;
  wire [32:0] v_463;
  wire [31:0] v_464;
  wire [38:0] v_465;
  wire [35:0] v_466;
  wire [3:0] v_467;
  wire [35:0] v_468;
  wire [38:0] v_469;
  wire [31:0] v_470;
  wire [2:0] v_471;
  wire [1:0] v_472;
  wire [2:0] v_473;
  wire [0:0] v_474;
  wire [77:0] v_475;
  wire [38:0] v_476;
  wire [5:0] v_477;
  wire [38:0] v_478;
  wire [77:0] v_479;
  wire [38:0] v_480;
  wire [32:0] v_481;
  wire [0:0] v_482;
  wire [31:0] v_483;
  wire [38:0] v_484;
  wire [35:0] v_485;
  wire [3:0] v_486;
  wire [3:0] v_487;
  function [3:0] mux_487(input [0:0] sel);
    case (sel) 0: mux_487 = 4'h0; 1: mux_487 = v_492;
    endcase
  endfunction
  wire [0:0] v_488;
  wire [1:0] v_489;
  reg [0:0] v_490 = 1'h0;
  reg [0:0] v_491 = 1'h0;
  wire [3:0] v_492;
  wire [0:0] v_493;
  wire [1:0] v_494;
  wire [2:0] v_495;
  wire [0:0] v_496;
  wire [1:0] v_497;
  wire [0:0] v_498;
  wire [0:0] v_499;
  wire [3:0] v_500;
  wire [3:0] v_501;
  function [3:0] mux_501(input [0:0] sel);
    case (sel) 0: mux_501 = 4'h0; 1: mux_501 = 4'hf;
    endcase
  endfunction
  wire [0:0] v_502;
  wire [3:0] v_503;
  function [3:0] mux_503(input [0:0] sel);
    case (sel) 0: mux_503 = 4'h0; 1: mux_503 = v_505;
    endcase
  endfunction
  wire [0:0] v_504;
  wire [3:0] v_505;
  wire [0:0] v_506;
  wire [2:0] v_507;
  wire [0:0] v_508;
  wire [1:0] v_509;
  wire [0:0] v_510;
  wire [0:0] v_511;
  wire [31:0] v_512;
  wire [31:0] v_513;
  function [31:0] mux_513(input [0:0] sel);
    case (sel) 0: mux_513 = 32'h0; 1: mux_513 = v_515;
    endcase
  endfunction
  wire [0:0] v_514;
  wire [31:0] v_515;
  wire [7:0] v_516;
  reg [31:0] v_517 = 32'h0;
  wire [23:0] v_518;
  wire [15:0] v_519;
  wire [31:0] v_520;
  wire [31:0] v_521;
  function [31:0] mux_521(input [0:0] sel);
    case (sel) 0: mux_521 = 32'h0; 1: mux_521 = v_523;
    endcase
  endfunction
  wire [0:0] v_522;
  wire [31:0] v_523;
  wire [7:0] v_524;
  wire [23:0] v_525;
  wire [7:0] v_526;
  wire [15:0] v_527;
  wire [7:0] v_528;
  wire [31:0] v_529;
  function [31:0] mux_529(input [0:0] sel);
    case (sel) 0: mux_529 = 32'h0; 1: mux_529 = v_531;
    endcase
  endfunction
  wire [0:0] v_530;
  wire [31:0] v_531;
  wire [23:0] v_532;
  wire [15:0] v_533;
  wire [2:0] v_534;
  reg [0:0] v_535 = 1'h0;
  wire [32:0] v_536;
  wire [0:0] v_537;
  wire [32:0] v_538;
  wire [31:0] v_539;
  wire [38:0] v_540;
  wire [35:0] v_541;
  wire [3:0] v_542;
  wire [35:0] v_543;
  wire [38:0] v_544;
  wire [31:0] v_545;
  wire [2:0] v_546;
  wire [1:0] v_547;
  wire [2:0] v_548;
  wire [0:0] v_549;
  wire [32:0] v_550;
  wire [0:0] v_551;
  wire [32:0] v_552;
  wire [31:0] v_553;
  wire [38:0] v_554;
  wire [35:0] v_555;
  wire [3:0] v_556;
  wire [35:0] v_557;
  wire [38:0] v_558;
  wire [31:0] v_559;
  wire [2:0] v_560;
  wire [1:0] v_561;
  wire [2:0] v_562;
  wire [0:0] v_563;
  wire [77:0] v_564;
  wire [38:0] v_565;
  wire [5:0] v_566;
  wire [38:0] v_567;
  wire [77:0] v_568;
  function [77:0] mux_568(input [0:0] sel);
    case (sel) 0: mux_568 = v_570; 1: mux_568 = v_588;
    endcase
  endfunction
  wire [0:0] v_569;
  wire [77:0] v_570;
  wire [38:0] v_571;
  wire [5:0] v_572;
  wire [38:0] v_573;
  wire [32:0] v_574;
  wire [0:0] v_575;
  wire [32:0] v_576;
  wire [31:0] v_577;
  wire [38:0] v_578;
  wire [35:0] v_579;
  wire [3:0] v_580;
  wire [35:0] v_581;
  wire [38:0] v_582;
  wire [31:0] v_583;
  wire [2:0] v_584;
  wire [1:0] v_585;
  wire [2:0] v_586;
  wire [0:0] v_587;
  wire [77:0] v_588;
  wire [38:0] v_589;
  wire [5:0] v_590;
  wire [38:0] v_591;
  wire [32:0] v_592;
  wire [0:0] v_593;
  wire [32:0] v_594;
  wire [31:0] v_595;
  wire [38:0] v_596;
  wire [35:0] v_597;
  wire [3:0] v_598;
  wire [35:0] v_599;
  wire [38:0] v_600;
  wire [31:0] v_601;
  wire [2:0] v_602;
  wire [1:0] v_603;
  wire [2:0] v_604;
  wire [0:0] v_605;
  wire [32:0] v_606;
  wire [0:0] v_607;
  wire [32:0] v_608;
  wire [31:0] v_609;
  wire [38:0] v_610;
  wire [35:0] v_611;
  wire [3:0] v_612;
  wire [35:0] v_613;
  wire [38:0] v_614;
  wire [31:0] v_615;
  wire [2:0] v_616;
  wire [1:0] v_617;
  wire [2:0] v_618;
  wire [0:0] v_619;
  wire [32:0] v_620;
  wire [0:0] v_621;
  wire [32:0] v_622;
  wire [31:0] v_623;
  wire [38:0] v_624;
  wire [35:0] v_625;
  wire [3:0] v_626;
  wire [35:0] v_627;
  wire [38:0] v_628;
  wire [31:0] v_629;
  wire [2:0] v_630;
  wire [1:0] v_631;
  wire [2:0] v_632;
  wire [0:0] v_633;
  wire [0:0] v_634;
  wire [0:0] v_635;
  wire [0:0] v_636;
  reg [0:0] v_637 = 1'h0;
  wire [0:0] v_638;
  wire [0:0] v_639;
  wire [0:0] v_640;
  wire [0:0] v_641;
  wire [0:0] v_642;
  wire [0:0] v_643;
  wire [0:0] v_644;
  wire [0:0] v_645;
  wire [0:0] v_646;
  wire [0:0] v_647;
  wire [0:0] v_648;
  wire [0:0] v_649;
  wire [0:0] v_650;
  wire [0:0] v_651;
  wire [0:0] v_652;
  wire [0:0] v_653;
  wire [0:0] v_654;
  wire [0:0] v_655;
  wire [0:0] v_656;
  wire [0:0] v_657;
  wire [0:0] v_658;
  wire [0:0] v_659;
  wire [0:0] v_660;
  wire [0:0] v_661;
  wire [0:0] v_662;
  wire [0:0] v_663;
  wire [0:0] v_664;
  function [0:0] mux_664(input [0:0] sel);
    case (sel) 0: mux_664 = 1'h0; 1: mux_664 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_665;
  function [0:0] mux_665(input [0:0] sel);
    case (sel) 0: mux_665 = 1'h0; 1: mux_665 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_666;
  function [0:0] mux_666(input [0:0] sel);
    case (sel) 0: mux_666 = 1'h0; 1: mux_666 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_667;
  wire [0:0] v_668;
  wire [0:0] v_669;
  wire [0:0] v_670;
  function [0:0] mux_670(input [0:0] sel);
    case (sel) 0: mux_670 = 1'h0; 1: mux_670 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_671;
  wire [0:0] v_672;
  wire [0:0] v_673;
  function [0:0] mux_673(input [0:0] sel);
    case (sel) 0: mux_673 = 1'h0; 1: mux_673 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_674;
  wire [0:0] v_675;
  wire [0:0] v_676;
  wire [31:0] v_677;
  wire [0:0] v_678;
  wire [0:0] v_679;
  reg [0:0] v_680 = 1'h0;
  wire [0:0] v_681;
  wire [0:0] v_682;
  wire [0:0] act_683;
  wire [0:0] v_684;
  wire [11:0] v_685;
  wire [0:0] v_686;
  wire [0:0] v_687;
  wire [0:0] v_688;
  wire [0:0] v_689;
  wire [0:0] v_690;
  wire [0:0] v_691;
  function [0:0] mux_691(input [0:0] sel);
    case (sel) 0: mux_691 = 1'h0; 1: mux_691 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_692;
  wire [0:0] v_693;
  wire [0:0] v_694;
  function [0:0] mux_694(input [0:0] sel);
    case (sel) 0: mux_694 = 1'h0; 1: mux_694 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_695;
  wire [0:0] v_696;
  wire [0:0] v_697;
  wire [0:0] v_698;
  function [0:0] mux_698(input [0:0] sel);
    case (sel) 0: mux_698 = 1'h0; 1: mux_698 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_699;
  function [0:0] mux_699(input [0:0] sel);
    case (sel) 0: mux_699 = 1'h0; 1: mux_699 = 1'h0;
    endcase
  endfunction
  wire [31:0] v_700;
  function [31:0] mux_700(input [0:0] sel);
    case (sel) 0: mux_700 = 32'h0; 1: mux_700 = v_714;
    endcase
  endfunction
  wire [0:0] v_701;
  wire [0:0] v_702;
  wire [4:0] v_703;
  wire [0:0] v_704;
  wire [3:0] v_705;
  wire [0:0] v_706;
  wire [2:0] v_707;
  wire [0:0] v_708;
  wire [1:0] v_709;
  wire [0:0] v_710;
  wire [0:0] v_711;
  wire [0:0] v_712;
  wire [0:0] v_713;
  reg [31:0] v_714 = 32'h0;
  wire [0:0] v_715;
  wire [0:0] v_716;
  wire [0:0] v_717;
  reg [0:0] v_718 = 1'h0;
  wire [0:0] v_719;
  wire [0:0] v_720;
  wire [0:0] v_721;
  wire [0:0] v_722;
  wire [0:0] v_723;
  wire [0:0] v_724;
  wire [0:0] v_725;
  wire [0:0] v_726;
  wire [0:0] v_727;
  wire [0:0] v_728;
  wire [0:0] v_729;
  wire [0:0] v_730;
  wire [0:0] v_731;
  wire [0:0] v_732;
  wire [0:0] v_733;
  wire [0:0] v_734;
  wire [0:0] v_735;
  wire [0:0] v_736;
  wire [0:0] v_737;
  wire [0:0] v_738;
  wire [0:0] v_739;
  wire [0:0] v_740;
  wire [0:0] v_741;
  wire [0:0] v_742;
  wire [0:0] v_743;
  wire [0:0] v_744;
  wire [0:0] v_745;
  wire [0:0] v_746;
  wire [0:0] v_747;
  wire [0:0] v_748;
  wire [0:0] v_749;
  wire [0:0] v_750;
  wire [0:0] v_751;
  wire [0:0] v_752;
  wire [0:0] v_753;
  wire [0:0] v_754;
  wire [0:0] v_755;
  wire [0:0] v_756;
  wire [0:0] v_757;
  wire [0:0] v_758;
  wire [0:0] v_759;
  wire [0:0] v_760;
  wire [0:0] v_761;
  wire [0:0] v_762;
  wire [0:0] v_763;
  wire [0:0] v_764;
  wire [0:0] v_765;
  wire [0:0] v_766;
  wire [0:0] v_767;
  reg [0:0] v_768 = 1'h0;
  wire [0:0] v_769;
  wire [31:0] v_770;
  wire [31:0] v_771;
  function [31:0] mux_771(input [0:0] sel);
    case (sel) 0: mux_771 = 32'h0; 1: mux_771 = v_772;
    endcase
  endfunction
  wire [31:0] v_772;
  wire [31:0] v_773;
  wire [31:0] v_774;
  function [31:0] mux_774(input [0:0] sel);
    case (sel) 0: mux_774 = 32'h0; 1: mux_774 = v_91;
    endcase
  endfunction
  wire [31:0] v_775;
  function [31:0] mux_775(input [0:0] sel);
    case (sel) 0: mux_775 = 32'h0; 1: mux_775 = v_776;
    endcase
  endfunction
  wire [31:0] v_776;
  wire [31:0] v_777;
  wire [31:0] v_778;
  function [31:0] mux_778(input [0:0] sel);
    case (sel) 0: mux_778 = 32'h0; 1: mux_778 = v_792;
    endcase
  endfunction
  wire [0:0] v_779;
  wire [0:0] v_780;
  wire [4:0] v_781;
  wire [0:0] v_782;
  wire [3:0] v_783;
  wire [0:0] v_784;
  wire [2:0] v_785;
  wire [0:0] v_786;
  wire [1:0] v_787;
  wire [0:0] v_788;
  wire [0:0] v_789;
  wire [0:0] v_790;
  wire [0:0] v_791;
  reg [31:0] v_792 = 32'h0;
  wire [0:0] v_793;
  wire [0:0] v_794;
  wire [31:0] v_795;
  function [31:0] mux_795(input [0:0] sel);
    case (sel) 0: mux_795 = 32'h0; 1: mux_795 = v_809;
    endcase
  endfunction
  wire [0:0] v_796;
  wire [0:0] v_797;
  wire [4:0] v_798;
  wire [0:0] v_799;
  wire [3:0] v_800;
  wire [0:0] v_801;
  wire [2:0] v_802;
  wire [0:0] v_803;
  wire [1:0] v_804;
  wire [0:0] v_805;
  wire [0:0] v_806;
  wire [0:0] v_807;
  wire [0:0] v_808;
  reg [31:0] v_809 = 32'h0;
  wire [0:0] v_810;
  wire [0:0] v_811;
  wire [31:0] v_812;
  wire [31:0] v_813;
  wire [31:0] v_814;
  function [31:0] mux_814(input [0:0] sel);
    case (sel) 0: mux_814 = 32'h0; 1: mux_814 = v_830;
    endcase
  endfunction
  wire [0:0] v_815;
  wire [0:0] v_816;
  wire [4:0] v_817;
  wire [0:0] v_818;
  wire [3:0] v_819;
  wire [0:0] v_820;
  wire [2:0] v_821;
  wire [0:0] v_822;
  wire [1:0] v_823;
  wire [0:0] v_824;
  wire [0:0] v_825;
  wire [0:0] v_826;
  wire [0:0] v_827;
  reg [0:0] v_828 = 1'h0;
  wire [0:0] v_829;
  wire [31:0] v_830;
  reg [31:0] v_831 = 32'h0;
  reg [31:0] v_832 = 32'h0;
  wire [31:0] v_833;
  function [31:0] mux_833(input [0:0] sel);
    case (sel) 0: mux_833 = 32'h0; 1: mux_833 = v_858;
    endcase
  endfunction
  wire [0:0] v_834;
  wire [0:0] v_835;
  wire [4:0] v_836;
  wire [0:0] v_837;
  wire [3:0] v_838;
  wire [0:0] v_839;
  wire [2:0] v_840;
  wire [0:0] v_841;
  wire [1:0] v_842;
  wire [0:0] v_843;
  wire [0:0] v_844;
  wire [0:0] v_845;
  wire [0:0] v_846;
  reg [0:0] v_847 = 1'h0;
  wire [0:0] v_848;
  wire [0:0] v_849;
  wire [0:0] v_850;
  wire [0:0] v_851;
  wire [0:0] v_852;
  wire [0:0] v_853;
  wire [0:0] v_854;
  reg [0:0] v_855 = 1'h0;
  wire [0:0] v_856;
  wire [0:0] v_857;
  wire [31:0] v_858;
  wire [32:0] v_859;
  wire [32:0] v_860;
  wire [0:0] v_861;
  function [0:0] mux_861(input [0:0] sel);
    case (sel) 0: mux_861 = 1'h0; 1: mux_861 = v_863;
    endcase
  endfunction
  wire [0:0] v_862;
  wire [0:0] v_863;
  wire [4:0] v_864;
  wire [31:0] v_865;
  wire [31:0] v_866;
  function [31:0] mux_866(input [0:0] sel);
    case (sel) 0: mux_866 = 32'h0; 1: mux_866 = v_887;
    endcase
  endfunction
  wire [0:0] v_867;
  wire [0:0] v_868;
  wire [4:0] v_869;
  wire [0:0] v_870;
  wire [3:0] v_871;
  wire [0:0] v_872;
  wire [2:0] v_873;
  wire [0:0] v_874;
  wire [1:0] v_875;
  wire [0:0] v_876;
  wire [0:0] v_877;
  wire [0:0] v_878;
  wire [0:0] v_879;
  reg [0:0] v_880 = 1'h0;
  wire [0:0] v_881;
  wire [0:0] v_882;
  wire [0:0] v_883;
  wire [0:0] v_884;
  wire [0:0] v_885;
  wire [0:0] v_886;
  wire [31:0] v_887;
  wire [4:0] v_888;
  wire [31:0] v_889;
  function [31:0] mux_889(input [0:0] sel);
    case (sel) 0: mux_889 = 32'h0; 1: mux_889 = v_904;
    endcase
  endfunction
  wire [0:0] v_890;
  wire [0:0] v_891;
  wire [4:0] v_892;
  wire [0:0] v_893;
  wire [3:0] v_894;
  wire [0:0] v_895;
  wire [2:0] v_896;
  wire [0:0] v_897;
  wire [1:0] v_898;
  wire [0:0] v_899;
  wire [0:0] v_900;
  wire [0:0] v_901;
  wire [0:0] v_902;
  reg [0:0] v_903 = 1'h0;
  wire [31:0] v_904;
  wire [31:0] v_905;
  wire [31:0] v_906;
  wire [31:0] v_907;
  wire [31:0] v_908;
  function [31:0] mux_908(input [0:0] sel);
    case (sel) 0: mux_908 = 32'h0; 1: mux_908 = v_115;
    endcase
  endfunction
  wire [0:0] v_909;
  wire [0:0] v_910;
  wire [4:0] v_911;
  wire [0:0] v_912;
  wire [3:0] v_913;
  wire [0:0] v_914;
  wire [2:0] v_915;
  wire [0:0] v_916;
  wire [1:0] v_917;
  wire [0:0] v_918;
  wire [0:0] v_919;
  wire [0:0] v_920;
  wire [0:0] v_921;
  reg [0:0] v_922 = 1'h0;
  wire [31:0] v_923;
  function [31:0] mux_923(input [0:0] sel);
    case (sel) 0: mux_923 = 32'h0; 1: mux_923 = v_941;
    endcase
  endfunction
  wire [0:0] v_924;
  wire [0:0] v_925;
  wire [4:0] v_926;
  wire [0:0] v_927;
  wire [3:0] v_928;
  wire [0:0] v_929;
  wire [2:0] v_930;
  wire [0:0] v_931;
  wire [1:0] v_932;
  wire [0:0] v_933;
  wire [0:0] v_934;
  wire [0:0] v_935;
  wire [0:0] v_936;
  reg [0:0] v_937 = 1'h0;
  wire [0:0] v_938;
  wire [0:0] v_939;
  wire [0:0] v_940;
  wire [31:0] v_941;
  wire [31:0] v_942;
  wire [31:0] v_943;
  function [31:0] mux_943(input [0:0] sel);
    case (sel) 0: mux_943 = 32'h0; 1: mux_943 = v_962;
    endcase
  endfunction
  wire [0:0] v_944;
  wire [0:0] v_945;
  wire [4:0] v_946;
  wire [0:0] v_947;
  wire [3:0] v_948;
  wire [0:0] v_949;
  wire [2:0] v_950;
  wire [0:0] v_951;
  wire [1:0] v_952;
  wire [0:0] v_953;
  wire [0:0] v_954;
  wire [0:0] v_955;
  wire [0:0] v_956;
  reg [0:0] v_957 = 1'h0;
  wire [0:0] v_958;
  wire [0:0] v_959;
  wire [0:0] v_960;
  wire [0:0] v_961;
  wire [31:0] v_962;
  wire [31:0] v_963;
  function [31:0] mux_963(input [0:0] sel);
    case (sel) 0: mux_963 = 32'h0; 1: mux_963 = v_980;
    endcase
  endfunction
  wire [0:0] v_964;
  wire [0:0] v_965;
  wire [4:0] v_966;
  wire [0:0] v_967;
  wire [3:0] v_968;
  wire [0:0] v_969;
  wire [2:0] v_970;
  wire [0:0] v_971;
  wire [1:0] v_972;
  wire [0:0] v_973;
  wire [0:0] v_974;
  wire [0:0] v_975;
  wire [0:0] v_976;
  reg [0:0] v_977 = 1'h0;
  wire [0:0] v_978;
  wire [0:0] v_979;
  wire [31:0] v_980;
  wire [31:0] v_981;
  wire [31:0] v_982;
  wire [31:0] v_983;
  function [31:0] mux_983(input [0:0] sel);
    case (sel) 0: mux_983 = 32'h0; 1: mux_983 = v_1006;
    endcase
  endfunction
  wire [0:0] v_984;
  wire [0:0] v_985;
  wire [4:0] v_986;
  wire [0:0] v_987;
  wire [3:0] v_988;
  wire [0:0] v_989;
  wire [2:0] v_990;
  wire [0:0] v_991;
  wire [1:0] v_992;
  wire [0:0] v_993;
  wire [0:0] v_994;
  wire [0:0] v_995;
  wire [0:0] v_996;
  reg [0:0] v_997 = 1'h0;
  wire [0:0] v_998;
  wire [0:0] v_999;
  wire [0:0] v_1000;
  wire [0:0] v_1001;
  wire [0:0] v_1002;
  reg [0:0] v_1003 = 1'h0;
  wire [0:0] v_1004;
  wire [0:0] v_1005;
  wire [31:0] v_1006;
  wire [0:0] v_1007;
  wire [32:0] v_1008;
  wire [32:0] v_1009;
  wire [32:0] v_1010;
  wire [0:0] v_1011;
  function [0:0] mux_1011(input [0:0] sel);
    case (sel) 0: mux_1011 = v_1025; 1: mux_1011 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1012;
  wire [0:0] v_1013;
  reg [0:0] v_1014 = 1'h0;
  wire [0:0] v_1015;
  wire [0:0] v_1016;
  wire [0:0] v_1017;
  wire [0:0] v_1018;
  wire [0:0] v_1019;
  reg [0:0] v_1020 = 1'h0;
  wire [0:0] v_1021;
  wire [0:0] v_1022;
  wire [0:0] v_1023;
  wire [0:0] v_1024;
  wire [0:0] v_1025;
  wire [32:0] v_1026;
  function [32:0] mux_1026(input [0:0] sel);
    case (sel) 0: mux_1026 = v_1032; 1: mux_1026 = v_1033;
    endcase
  endfunction
  wire [0:0] v_1027;
  reg [0:0] v_1028 = 1'h0;
  wire [0:0] v_1029;
  wire [0:0] v_1030;
  wire [0:0] v_1031;
  wire [32:0] v_1032;
  wire [32:0] v_1033;
  wire [0:0] v_1034;
  function [0:0] mux_1034(input [0:0] sel);
    case (sel) 0: mux_1034 = v_1035; 1: mux_1034 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1035;
  wire [32:0] v_1036;
  function [32:0] mux_1036(input [0:0] sel);
    case (sel) 0: mux_1036 = 33'h1; 1: mux_1036 = 33'h0;
    endcase
  endfunction
  wire [31:0] v_1037;
  function [31:0] mux_1037(input [0:0] sel);
    case (sel) 0: mux_1037 = 32'h0; 1: mux_1037 = v_1058;
    endcase
  endfunction
  wire [0:0] v_1038;
  wire [0:0] v_1039;
  wire [4:0] v_1040;
  wire [0:0] v_1041;
  wire [3:0] v_1042;
  wire [0:0] v_1043;
  wire [2:0] v_1044;
  wire [0:0] v_1045;
  wire [1:0] v_1046;
  wire [0:0] v_1047;
  wire [0:0] v_1048;
  wire [0:0] v_1049;
  wire [0:0] v_1050;
  wire [0:0] v_1051;
  reg [0:0] v_1052 = 1'h0;
  wire [0:0] v_1053;
  wire [0:0] v_1054;
  wire [0:0] v_1055;
  wire [0:0] v_1056;
  wire [0:0] v_1057;
  wire [31:0] v_1058;
  wire [31:0] v_1059;
  wire [31:0] v_1060;
  function [31:0] mux_1060(input [0:0] sel);
    case (sel)
      0: mux_1060 = 32'h0;
      1: mux_1060 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_1061;
  wire [31:0] v_1062;
  wire [31:0] v_1063;
  function [31:0] mux_1063(input [0:0] sel);
    case (sel) 0: mux_1063 = 32'h0; 1: mux_1063 = v_1064;
    endcase
  endfunction
  wire [31:0] v_1064;
  wire [7:0] v_1065;
  wire [31:0] v_1066;
  function [31:0] mux_1066(input [0:0] sel);
    case (sel) 0: mux_1066 = 32'h0; 1: mux_1066 = v_1080;
    endcase
  endfunction
  wire [0:0] v_1067;
  wire [0:0] v_1068;
  wire [4:0] v_1069;
  wire [0:0] v_1070;
  wire [3:0] v_1071;
  wire [0:0] v_1072;
  wire [2:0] v_1073;
  wire [0:0] v_1074;
  wire [1:0] v_1075;
  wire [0:0] v_1076;
  wire [0:0] v_1077;
  wire [0:0] v_1078;
  wire [0:0] v_1079;
  wire [31:0] v_1080;
  wire [0:0] v_1081;
  wire [31:0] v_1082;
  function [31:0] mux_1082(input [0:0] sel);
    case (sel) 0: mux_1082 = 32'h0; 1: mux_1082 = v_1083;
    endcase
  endfunction
  wire [31:0] v_1083;
  wire [31:0] v_1084;
  function [31:0] mux_1084(input [0:0] sel);
    case (sel) 0: mux_1084 = 32'h0; 1: mux_1084 = v_1085;
    endcase
  endfunction
  wire [31:0] v_1085;
  wire [37:0] v_1086;
  function [37:0] mux_1086(input [0:0] sel);
    case (sel) 0: mux_1086 = v_1087; 1: mux_1086 = v_1282;
    endcase
  endfunction
  wire [37:0] v_1087;
  wire [5:0] v_1088;
  wire [37:0] v_1089;
  function [37:0] mux_1089(input [0:0] sel);
    case (sel) 0: mux_1089 = v_1090; 1: mux_1089 = v_1149;
    endcase
  endfunction
  wire [37:0] v_1090;
  wire [5:0] v_1091;
  wire [69:0] v_1092;
  wire [72:0] v_1093;
  wire [69:0] v_1094;
  wire [5:0] v_1095;
  wire [69:0] v_1096;
  reg [72:0] v_1097 = 73'h0;
  wire [72:0] v_1098;
  wire [69:0] v_1099;
  wire [5:0] v_1100;
  wire [69:0] v_1101;
  wire [72:0] v_1102;
  wire [69:0] v_1103;
  wire [63:0] v_1104;
  wire [2:0] v_1105;
  wire [0:0] v_1106;
  wire [1:0] v_1107;
  reg [0:0] v_1108 = 1'h0;
  reg [0:0] v_1109 = 1'h0;
  wire [1:0] v_1110;
  wire [0:0] v_1111;
  wire [0:0] v_1112;
  wire [63:0] v_1113;
  wire [31:0] v_1114;
  wire [63:0] v_1115;
  wire [31:0] v_1116;
  wire [2:0] v_1117;
  wire [0:0] v_1118;
  wire [2:0] v_1119;
  wire [1:0] v_1120;
  wire [0:0] v_1121;
  wire [1:0] v_1122;
  wire [0:0] v_1123;
  wire [63:0] v_1124;
  wire [31:0] v_1125;
  wire [63:0] v_1126;
  wire [31:0] v_1127;
  wire [2:0] v_1128;
  wire [0:0] v_1129;
  wire [2:0] v_1130;
  wire [1:0] v_1131;
  wire [0:0] v_1132;
  wire [1:0] v_1133;
  wire [0:0] v_1134;
  wire [31:0] v_1135;
  function [31:0] mux_1135(input [0:0] sel);
    case (sel) 0: mux_1135 = v_1138; 1: mux_1135 = v_1148;
    endcase
  endfunction
  wire [0:0] v_1136;
  wire [2:0] v_1137;
  wire [31:0] v_1138;
  reg [63:0] v_1139 = 64'h0;
  wire [63:0] v_1140;
  wire [65:0] v_1141;
  wire [32:0] v_1142;
  wire [0:0] v_1143;
  function [0:0] mux_1143(input [0:0] sel);
    case (sel) 0: mux_1143 = v_1144; 1: mux_1143 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1144;
  wire [32:0] v_1145;
  wire [0:0] v_1146;
  function [0:0] mux_1146(input [0:0] sel);
    case (sel) 0: mux_1146 = v_1147; 1: mux_1146 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1147;
  wire [31:0] v_1148;
  wire [37:0] v_1149;
  wire [5:0] v_1150;
  wire [38:0] v_1151;
  wire [77:0] v_1152;
  wire [38:0] v_1153;
  wire [5:0] v_1154;
  wire [38:0] v_1155;
  reg [77:0] v_1156 = 78'h0;
  wire [0:0] v_1157;
  wire [77:0] v_1158;
  wire [38:0] v_1159;
  wire [5:0] v_1160;
  wire [38:0] v_1161;
  wire [77:0] v_1162;
  wire [38:0] v_1163;
  wire [5:0] v_1164;
  wire [32:0] v_1165;
  wire [31:0] v_1166;
  wire [38:0] v_1167;
  wire [35:0] v_1168;
  wire [3:0] v_1169;
  wire [35:0] v_1170;
  wire [38:0] v_1171;
  wire [31:0] v_1172;
  wire [2:0] v_1173;
  wire [1:0] v_1174;
  wire [2:0] v_1175;
  wire [0:0] v_1176;
  wire [32:0] v_1177;
  wire [0:0] v_1178;
  wire [32:0] v_1179;
  wire [31:0] v_1180;
  wire [38:0] v_1181;
  wire [35:0] v_1182;
  wire [3:0] v_1183;
  wire [35:0] v_1184;
  wire [38:0] v_1185;
  wire [31:0] v_1186;
  wire [2:0] v_1187;
  wire [1:0] v_1188;
  wire [2:0] v_1189;
  wire [0:0] v_1190;
  wire [32:0] v_1191;
  wire [0:0] v_1192;
  wire [32:0] v_1193;
  wire [31:0] v_1194;
  wire [38:0] v_1195;
  wire [35:0] v_1196;
  wire [3:0] v_1197;
  wire [35:0] v_1198;
  wire [38:0] v_1199;
  wire [31:0] v_1200;
  wire [2:0] v_1201;
  wire [1:0] v_1202;
  wire [2:0] v_1203;
  wire [0:0] v_1204;
  wire [31:0] v_1205;
  wire [31:0] v_1206;
  function [31:0] mux_1206(input [0:0] sel);
    case (sel) 0: mux_1206 = 32'h0; 1: mux_1206 = v_1211;
    endcase
  endfunction
  wire [0:0] v_1207;
  wire [1:0] v_1208;
  wire [2:0] v_1209;
  wire [38:0] v_1210;
  wire [31:0] v_1211;
  wire [23:0] v_1212;
  function [23:0] mux_1212(input [0:0] sel);
    case (sel) 0: mux_1212 = v_1214; 1: mux_1212 = 24'h0;
    endcase
  endfunction
  wire [0:0] v_1213;
  wire [23:0] v_1214;
  wire [0:0] v_1215;
  wire [7:0] v_1216;
  wire [7:0] v_1217;
  wire [7:0] v_1218;
  function [7:0] mux_1218(input [0:0] sel);
    case (sel) 0: mux_1218 = 8'h0; 1: mux_1218 = v_1223;
    endcase
  endfunction
  wire [0:0] v_1219;
  wire [1:0] v_1220;
  wire [31:0] v_1221;
  wire [32:0] v_1222;
  wire [7:0] v_1223;
  wire [31:0] v_1224;
  wire [8:0] v_1225;
  wire [8:0] v_1226;
  function [8:0] mux_1226(input [0:0] sel);
    case (sel) 0: mux_1226 = 9'h0; 1: mux_1226 = 9'bxxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_1227;
  wire [0:0] v_1228;
  wire [0:0] v_1229;
  wire [0:0] v_1230;
  wire [0:0] v_1231;
  wire [8:0] v_1232;
  wire [8:0] v_1233;
  function [8:0] mux_1233(input [0:0] sel);
    case (sel) 0: mux_1233 = 9'h0; 1: mux_1233 = v_1234;
    endcase
  endfunction
  wire [8:0] v_1234;
  wire [29:0] v_1235;
  wire [8:0] v_1236;
  function [8:0] mux_1236(input [0:0] sel);
    case (sel) 0: mux_1236 = 9'h0; 1: mux_1236 = v_1234;
    endcase
  endfunction
  wire [31:0] v_1237;
  wire [31:0] v_1238;
  function [31:0] mux_1238(input [0:0] sel);
    case (sel) 0: mux_1238 = 32'h0; 1: mux_1238 = v_1172;
    endcase
  endfunction
  wire [31:0] v_1239;
  function [31:0] mux_1239(input [0:0] sel);
    case (sel)
      0: mux_1239 = 32'h0;
      1: mux_1239 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_1240;
  wire [0:0] v_1241;
  wire [0:0] v_1242;
  function [0:0] mux_1242(input [0:0] sel);
    case (sel) 0: mux_1242 = 1'h0; 1: mux_1242 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1243;
  function [0:0] mux_1243(input [0:0] sel);
    case (sel) 0: mux_1243 = 1'h0; 1: mux_1243 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1244;
  wire [0:0] v_1245;
  wire [0:0] v_1246;
  function [0:0] mux_1246(input [0:0] sel);
    case (sel) 0: mux_1246 = 1'h0; 1: mux_1246 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1247;
  wire [0:0] v_1248;
  function [0:0] mux_1248(input [0:0] sel);
    case (sel) 0: mux_1248 = 1'h0; 1: mux_1248 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1249;
  wire [3:0] v_1250;
  wire [3:0] v_1251;
  function [3:0] mux_1251(input [0:0] sel);
    case (sel) 0: mux_1251 = 4'h0; 1: mux_1251 = v_1169;
    endcase
  endfunction
  wire [3:0] v_1252;
  function [3:0] mux_1252(input [0:0] sel);
    case (sel) 0: mux_1252 = 4'h0; 1: mux_1252 = 4'h0;
    endcase
  endfunction
  wire [0:0] v_1253;
  wire [7:0] v_1254;
  function [7:0] mux_1254(input [0:0] sel);
    case (sel) 0: mux_1254 = 8'h0; 1: mux_1254 = v_1256;
    endcase
  endfunction
  wire [0:0] v_1255;
  wire [7:0] v_1256;
  wire [7:0] v_1257;
  wire [7:0] v_1258;
  function [7:0] mux_1258(input [0:0] sel);
    case (sel) 0: mux_1258 = 8'h0; 1: mux_1258 = v_1260;
    endcase
  endfunction
  wire [0:0] v_1259;
  wire [7:0] v_1260;
  wire [7:0] v_1261;
  function [7:0] mux_1261(input [0:0] sel);
    case (sel) 0: mux_1261 = 8'h0; 1: mux_1261 = v_1263;
    endcase
  endfunction
  wire [0:0] v_1262;
  wire [7:0] v_1263;
  wire [31:0] v_1264;
  wire [31:0] v_1265;
  function [31:0] mux_1265(input [0:0] sel);
    case (sel) 0: mux_1265 = 32'h0; 1: mux_1265 = v_1267;
    endcase
  endfunction
  wire [0:0] v_1266;
  wire [31:0] v_1267;
  wire [23:0] v_1268;
  wire [15:0] v_1269;
  wire [31:0] v_1270;
  function [31:0] mux_1270(input [0:0] sel);
    case (sel) 0: mux_1270 = 32'h0; 1: mux_1270 = v_1272;
    endcase
  endfunction
  wire [0:0] v_1271;
  wire [31:0] v_1272;
  wire [15:0] v_1273;
  function [15:0] mux_1273(input [0:0] sel);
    case (sel) 0: mux_1273 = v_1274; 1: mux_1273 = 16'h0;
    endcase
  endfunction
  wire [15:0] v_1274;
  wire [0:0] v_1275;
  wire [15:0] v_1276;
  function [15:0] mux_1276(input [0:0] sel);
    case (sel) 0: mux_1276 = v_1279; 1: mux_1276 = v_1280;
    endcase
  endfunction
  wire [0:0] v_1277;
  wire [0:0] v_1278;
  wire [15:0] v_1279;
  wire [15:0] v_1280;
  wire [31:0] v_1281;
  wire [37:0] v_1282;
  reg [5:0] v_1283 = 6'h0;
  reg [31:0] v_1284 = 32'h0;
  wire [31:0] v_1285;
  function [31:0] mux_1285(input [0:0] sel);
    case (sel) 0: mux_1285 = v_1336; 1: mux_1285 = v_1357;
    endcase
  endfunction
  reg [0:0] v_1286 = 1'h0;
  wire [0:0] v_1287;
  wire [0:0] v_1288;
  wire [0:0] v_1289;
  reg [0:0] v_1290 = 1'h0;
  wire [0:0] v_1291;
  wire [1:0] v_1292;
  wire [1:0] v_1293;
  reg [0:0] v_1294 = 1'h0;
  reg [0:0] v_1295 = 1'h0;
  wire [0:0] v_1296;
  wire [0:0] v_1297;
  reg [31:0] v_1298 = 32'h0;
  wire [0:0] v_1299;
  wire [0:0] v_1300;
  wire [0:0] v_1301;
  wire [0:0] v_1302;
  wire [0:0] v_1303;
  wire [0:0] v_1304;
  wire [31:0] v_1305;
  wire [31:0] v_1306;
  function [31:0] mux_1306(input [0:0] sel);
    case (sel) 0: mux_1306 = 32'h0; 1: mux_1306 = v_517;
    endcase
  endfunction
  wire [31:0] v_1307;
  function [31:0] mux_1307(input [0:0] sel);
    case (sel) 0: mux_1307 = 32'h0; 1: mux_1307 = v_1308;
    endcase
  endfunction
  wire [31:0] v_1308;
  wire [31:0] v_1309;
  wire [0:0] v_1310;
  function [0:0] mux_1310(input [0:0] sel);
    case (sel) 0: mux_1310 = v_1313; 1: mux_1310 = v_1314;
    endcase
  endfunction
  reg [0:0] v_1311 = 1'h0;
  wire [0:0] v_1312;
  wire [0:0] v_1313;
  wire [0:0] v_1314;
  reg [31:0] v_1315 = 32'h0;
  wire [0:0] v_1316;
  wire [0:0] v_1317;
  wire [0:0] v_1318;
  wire [0:0] v_1319;
  wire [0:0] v_1320;
  wire [0:0] v_1321;
  reg [5:0] v_1322 = 6'h0;
  wire [0:0] v_1323;
  wire [5:0] v_1324;
  wire [5:0] v_1325;
  function [5:0] mux_1325(input [0:0] sel);
    case (sel) 0: mux_1325 = 6'h0; 1: mux_1325 = v_1326;
    endcase
  endfunction
  wire [5:0] v_1326;
  wire [5:0] v_1327;
  function [5:0] mux_1327(input [0:0] sel);
    case (sel) 0: mux_1327 = 6'h0; 1: mux_1327 = 6'h20;
    endcase
  endfunction
  wire [31:0] v_1328;
  wire [31:0] v_1329;
  function [31:0] mux_1329(input [0:0] sel);
    case (sel) 0: mux_1329 = 32'h0; 1: mux_1329 = v_1330;
    endcase
  endfunction
  wire [31:0] v_1330;
  wire [31:0] v_1331;
  wire [31:0] v_1332;
  wire [31:0] v_1333;
  function [31:0] mux_1333(input [0:0] sel);
    case (sel) 0: mux_1333 = 32'h0; 1: mux_1333 = v_91;
    endcase
  endfunction
  wire [31:0] v_1334;
  function [31:0] mux_1334(input [0:0] sel);
    case (sel) 0: mux_1334 = 32'h0; 1: mux_1334 = v_1335;
    endcase
  endfunction
  wire [31:0] v_1335;
  wire [31:0] v_1336;
  function [31:0] mux_1336(input [0:0] sel);
    case (sel) 0: mux_1336 = v_1337; 1: mux_1336 = v_1347;
    endcase
  endfunction
  reg [31:0] v_1337 = 32'h0;
  wire [0:0] v_1338;
  wire [31:0] v_1339;
  wire [31:0] v_1340;
  function [31:0] mux_1340(input [0:0] sel);
    case (sel) 0: mux_1340 = 32'h0; 1: mux_1340 = v_1341;
    endcase
  endfunction
  wire [31:0] v_1341;
  wire [31:0] v_1342;
  wire [31:0] v_1343;
  function [31:0] mux_1343(input [0:0] sel);
    case (sel) 0: mux_1343 = 32'h0; 1: mux_1343 = 32'h1;
    endcase
  endfunction
  wire [0:0] v_1344;
  wire [31:0] v_1345;
  wire [31:0] v_1346;
  reg [31:0] v_1347 = 32'h0;
  wire [0:0] v_1348;
  wire [31:0] v_1349;
  wire [31:0] v_1350;
  function [31:0] mux_1350(input [0:0] sel);
    case (sel) 0: mux_1350 = 32'h0; 1: mux_1350 = v_1351;
    endcase
  endfunction
  wire [31:0] v_1351;
  wire [31:0] v_1352;
  function [31:0] mux_1352(input [0:0] sel);
    case (sel) 0: mux_1352 = 32'h0; 1: mux_1352 = v_1298;
    endcase
  endfunction
  wire [31:0] v_1353;
  function [31:0] mux_1353(input [0:0] sel);
    case (sel) 0: mux_1353 = 32'h0; 1: mux_1353 = 32'h0;
    endcase
  endfunction
  wire [31:0] v_1354;
  wire [0:0] v_1355;
  wire [31:0] v_1356;
  function [31:0] mux_1356(input [0:0] sel);
    case (sel) 0: mux_1356 = 32'h0; 1: mux_1356 = 32'h0;
    endcase
  endfunction
  wire [31:0] v_1357;
  wire [31:0] v_1358;
  wire [31:0] v_1359;
  function [31:0] mux_1359(input [0:0] sel);
    case (sel)
      0: mux_1359 = 32'h0;
      1: mux_1359 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_1360;
  wire [31:0] v_1361;
  function [31:0] mux_1361(input [0:0] sel);
    case (sel)
      0: mux_1361 = 32'h0;
      1: mux_1361 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_1362;
  wire [0:0] v_1363;
  wire [0:0] v_1364;
  function [0:0] mux_1364(input [0:0] sel);
    case (sel) 0: mux_1364 = 1'h0; 1: mux_1364 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1365;
  function [0:0] mux_1365(input [0:0] sel);
    case (sel) 0: mux_1365 = 1'h0; 1: mux_1365 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1366;
  wire [0:0] v_1367;
  function [0:0] mux_1367(input [0:0] sel);
    case (sel) 0: mux_1367 = 1'h0; 1: mux_1367 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1368;
  reg [31:0] v_1369 = 32'h0;
  wire [31:0] v_1370;
  wire [31:0] v_1371;
  function [31:0] mux_1371(input [0:0] sel);
    case (sel) 0: mux_1371 = 32'h0; 1: mux_1371 = v_384;
    endcase
  endfunction
  wire [31:0] v_1372;
  function [31:0] mux_1372(input [0:0] sel);
    case (sel)
      0: mux_1372 = 32'h0;
      1: mux_1372 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_1373;
  wire [31:0] v_1374;
  wire [0:0] v_1375;
  wire [0:0] v_1376;
  wire [0:0] v_1377;
  wire [0:0] v_1378;
  wire [0:0] v_1379;
  wire [0:0] v_1380;
  wire [0:0] v_1381;
  wire [0:0] v_1382;
  wire [0:0] v_1383;
  wire [0:0] v_1384;
  wire [0:0] v_1385;
  wire [0:0] v_1386;
  wire [0:0] v_1387;
  wire [0:0] v_1388;
  wire [0:0] v_1389;
  wire [0:0] v_1390;
  wire [0:0] v_1391;
  wire [0:0] v_1392;
  wire [0:0] v_1393;
  wire [0:0] v_1394;
  wire [0:0] v_1395;
  wire [0:0] v_1396;
  wire [0:0] v_1397;
  wire [0:0] v_1398;
  wire [0:0] v_1399;
  wire [0:0] v_1400;
  wire [0:0] v_1401;
  wire [0:0] v_1402;
  wire [0:0] v_1403;
  wire [0:0] v_1404;
  wire [0:0] v_1405;
  wire [30:0] v_1406;
  wire [0:0] v_1407;
  wire [0:0] v_1408;
  wire [0:0] v_1409;
  wire [0:0] v_1410;
  wire [0:0] v_1411;
  wire [0:0] v_1412;
  wire [0:0] v_1413;
  wire [0:0] v_1414;
  wire [0:0] v_1415;
  wire [0:0] v_1416;
  wire [0:0] v_1417;
  wire [0:0] v_1418;
  wire [0:0] v_1419;
  wire [0:0] v_1420;
  wire [0:0] v_1421;
  wire [0:0] v_1422;
  wire [0:0] v_1423;
  wire [0:0] v_1424;
  wire [0:0] v_1425;
  wire [0:0] v_1426;
  wire [0:0] v_1427;
  wire [0:0] v_1428;
  wire [0:0] v_1429;
  wire [0:0] v_1430;
  wire [0:0] v_1431;
  wire [0:0] v_1432;
  wire [0:0] v_1433;
  wire [0:0] v_1434;
  wire [0:0] v_1435;
  wire [0:0] v_1436;
  wire [0:0] v_1437;
  wire [29:0] v_1438;
  wire [0:0] v_1439;
  wire [0:0] v_1440;
  wire [0:0] v_1441;
  wire [0:0] v_1442;
  wire [0:0] v_1443;
  wire [0:0] v_1444;
  wire [0:0] v_1445;
  wire [0:0] v_1446;
  wire [0:0] v_1447;
  wire [0:0] v_1448;
  wire [0:0] v_1449;
  wire [0:0] v_1450;
  wire [0:0] v_1451;
  wire [0:0] v_1452;
  wire [0:0] v_1453;
  wire [0:0] v_1454;
  wire [0:0] v_1455;
  wire [0:0] v_1456;
  wire [0:0] v_1457;
  wire [0:0] v_1458;
  wire [0:0] v_1459;
  wire [0:0] v_1460;
  wire [0:0] v_1461;
  wire [0:0] v_1462;
  wire [0:0] v_1463;
  wire [0:0] v_1464;
  wire [0:0] v_1465;
  wire [0:0] v_1466;
  wire [0:0] v_1467;
  wire [0:0] v_1468;
  wire [0:0] v_1469;
  wire [28:0] v_1470;
  wire [0:0] v_1471;
  wire [0:0] v_1472;
  wire [0:0] v_1473;
  wire [0:0] v_1474;
  wire [0:0] v_1475;
  wire [0:0] v_1476;
  wire [0:0] v_1477;
  wire [0:0] v_1478;
  wire [0:0] v_1479;
  wire [0:0] v_1480;
  wire [0:0] v_1481;
  wire [0:0] v_1482;
  wire [0:0] v_1483;
  wire [0:0] v_1484;
  wire [0:0] v_1485;
  wire [0:0] v_1486;
  wire [0:0] v_1487;
  wire [0:0] v_1488;
  wire [0:0] v_1489;
  wire [0:0] v_1490;
  wire [0:0] v_1491;
  wire [0:0] v_1492;
  wire [0:0] v_1493;
  wire [0:0] v_1494;
  wire [0:0] v_1495;
  wire [0:0] v_1496;
  wire [0:0] v_1497;
  wire [0:0] v_1498;
  wire [0:0] v_1499;
  wire [0:0] v_1500;
  wire [0:0] v_1501;
  wire [27:0] v_1502;
  wire [0:0] v_1503;
  wire [0:0] v_1504;
  wire [0:0] v_1505;
  wire [0:0] v_1506;
  wire [0:0] v_1507;
  wire [0:0] v_1508;
  wire [0:0] v_1509;
  wire [0:0] v_1510;
  wire [0:0] v_1511;
  wire [0:0] v_1512;
  wire [0:0] v_1513;
  wire [0:0] v_1514;
  wire [0:0] v_1515;
  wire [0:0] v_1516;
  wire [0:0] v_1517;
  wire [0:0] v_1518;
  wire [0:0] v_1519;
  wire [0:0] v_1520;
  wire [0:0] v_1521;
  wire [0:0] v_1522;
  wire [0:0] v_1523;
  wire [0:0] v_1524;
  wire [0:0] v_1525;
  wire [0:0] v_1526;
  wire [0:0] v_1527;
  wire [0:0] v_1528;
  wire [0:0] v_1529;
  wire [0:0] v_1530;
  wire [0:0] v_1531;
  wire [0:0] v_1532;
  wire [0:0] v_1533;
  wire [26:0] v_1534;
  wire [0:0] v_1535;
  wire [0:0] v_1536;
  wire [0:0] v_1537;
  wire [0:0] v_1538;
  wire [0:0] v_1539;
  wire [0:0] v_1540;
  wire [0:0] v_1541;
  wire [0:0] v_1542;
  wire [0:0] v_1543;
  wire [0:0] v_1544;
  wire [0:0] v_1545;
  wire [0:0] v_1546;
  wire [0:0] v_1547;
  wire [0:0] v_1548;
  wire [0:0] v_1549;
  wire [0:0] v_1550;
  wire [0:0] v_1551;
  wire [0:0] v_1552;
  wire [0:0] v_1553;
  wire [0:0] v_1554;
  wire [0:0] v_1555;
  wire [0:0] v_1556;
  wire [0:0] v_1557;
  wire [0:0] v_1558;
  wire [0:0] v_1559;
  wire [0:0] v_1560;
  wire [0:0] v_1561;
  wire [0:0] v_1562;
  wire [0:0] v_1563;
  wire [0:0] v_1564;
  wire [0:0] v_1565;
  wire [25:0] v_1566;
  wire [0:0] v_1567;
  wire [0:0] v_1568;
  wire [0:0] v_1569;
  wire [0:0] v_1570;
  wire [0:0] v_1571;
  wire [0:0] v_1572;
  wire [0:0] v_1573;
  wire [0:0] v_1574;
  wire [0:0] v_1575;
  wire [0:0] v_1576;
  wire [0:0] v_1577;
  wire [0:0] v_1578;
  wire [0:0] v_1579;
  wire [0:0] v_1580;
  wire [0:0] v_1581;
  wire [0:0] v_1582;
  wire [0:0] v_1583;
  wire [0:0] v_1584;
  wire [0:0] v_1585;
  wire [0:0] v_1586;
  wire [0:0] v_1587;
  wire [0:0] v_1588;
  wire [0:0] v_1589;
  wire [0:0] v_1590;
  wire [0:0] v_1591;
  wire [0:0] v_1592;
  wire [0:0] v_1593;
  wire [0:0] v_1594;
  wire [0:0] v_1595;
  wire [0:0] v_1596;
  wire [0:0] v_1597;
  wire [24:0] v_1598;
  wire [0:0] v_1599;
  wire [0:0] v_1600;
  wire [0:0] v_1601;
  wire [0:0] v_1602;
  wire [0:0] v_1603;
  wire [0:0] v_1604;
  wire [0:0] v_1605;
  wire [0:0] v_1606;
  wire [0:0] v_1607;
  wire [0:0] v_1608;
  wire [0:0] v_1609;
  wire [0:0] v_1610;
  wire [0:0] v_1611;
  wire [0:0] v_1612;
  wire [0:0] v_1613;
  wire [0:0] v_1614;
  wire [0:0] v_1615;
  wire [0:0] v_1616;
  wire [0:0] v_1617;
  wire [0:0] v_1618;
  wire [0:0] v_1619;
  wire [0:0] v_1620;
  wire [0:0] v_1621;
  wire [0:0] v_1622;
  wire [0:0] v_1623;
  wire [0:0] v_1624;
  wire [0:0] v_1625;
  wire [0:0] v_1626;
  wire [0:0] v_1627;
  wire [0:0] v_1628;
  wire [0:0] v_1629;
  wire [23:0] v_1630;
  wire [0:0] v_1631;
  wire [0:0] v_1632;
  wire [0:0] v_1633;
  wire [0:0] v_1634;
  wire [0:0] v_1635;
  wire [0:0] v_1636;
  wire [0:0] v_1637;
  wire [0:0] v_1638;
  wire [0:0] v_1639;
  wire [0:0] v_1640;
  wire [0:0] v_1641;
  wire [0:0] v_1642;
  wire [0:0] v_1643;
  wire [0:0] v_1644;
  wire [0:0] v_1645;
  wire [0:0] v_1646;
  wire [0:0] v_1647;
  wire [0:0] v_1648;
  wire [0:0] v_1649;
  wire [0:0] v_1650;
  wire [0:0] v_1651;
  wire [0:0] v_1652;
  wire [0:0] v_1653;
  wire [0:0] v_1654;
  wire [0:0] v_1655;
  wire [0:0] v_1656;
  wire [0:0] v_1657;
  wire [0:0] v_1658;
  wire [0:0] v_1659;
  wire [0:0] v_1660;
  wire [0:0] v_1661;
  wire [22:0] v_1662;
  wire [0:0] v_1663;
  wire [0:0] v_1664;
  wire [0:0] v_1665;
  wire [0:0] v_1666;
  wire [0:0] v_1667;
  wire [0:0] v_1668;
  wire [0:0] v_1669;
  wire [0:0] v_1670;
  wire [0:0] v_1671;
  wire [0:0] v_1672;
  wire [0:0] v_1673;
  wire [0:0] v_1674;
  wire [0:0] v_1675;
  wire [0:0] v_1676;
  wire [0:0] v_1677;
  wire [0:0] v_1678;
  wire [0:0] v_1679;
  wire [0:0] v_1680;
  wire [0:0] v_1681;
  wire [0:0] v_1682;
  wire [0:0] v_1683;
  wire [0:0] v_1684;
  wire [0:0] v_1685;
  wire [0:0] v_1686;
  wire [0:0] v_1687;
  wire [0:0] v_1688;
  wire [0:0] v_1689;
  wire [0:0] v_1690;
  wire [0:0] v_1691;
  wire [0:0] v_1692;
  wire [0:0] v_1693;
  wire [21:0] v_1694;
  wire [0:0] v_1695;
  wire [0:0] v_1696;
  wire [0:0] v_1697;
  wire [0:0] v_1698;
  wire [0:0] v_1699;
  wire [0:0] v_1700;
  wire [0:0] v_1701;
  wire [0:0] v_1702;
  wire [0:0] v_1703;
  wire [0:0] v_1704;
  wire [0:0] v_1705;
  wire [0:0] v_1706;
  wire [0:0] v_1707;
  wire [0:0] v_1708;
  wire [0:0] v_1709;
  wire [0:0] v_1710;
  wire [0:0] v_1711;
  wire [0:0] v_1712;
  wire [0:0] v_1713;
  wire [0:0] v_1714;
  wire [0:0] v_1715;
  wire [0:0] v_1716;
  wire [0:0] v_1717;
  wire [0:0] v_1718;
  wire [0:0] v_1719;
  wire [0:0] v_1720;
  wire [0:0] v_1721;
  wire [0:0] v_1722;
  wire [0:0] v_1723;
  wire [0:0] v_1724;
  wire [0:0] v_1725;
  wire [20:0] v_1726;
  wire [0:0] v_1727;
  wire [0:0] v_1728;
  wire [0:0] v_1729;
  wire [0:0] v_1730;
  wire [0:0] v_1731;
  wire [0:0] v_1732;
  wire [0:0] v_1733;
  wire [0:0] v_1734;
  wire [0:0] v_1735;
  wire [0:0] v_1736;
  wire [0:0] v_1737;
  wire [0:0] v_1738;
  wire [0:0] v_1739;
  wire [0:0] v_1740;
  wire [0:0] v_1741;
  wire [0:0] v_1742;
  wire [0:0] v_1743;
  wire [0:0] v_1744;
  wire [0:0] v_1745;
  wire [0:0] v_1746;
  wire [0:0] v_1747;
  wire [0:0] v_1748;
  wire [0:0] v_1749;
  wire [0:0] v_1750;
  wire [0:0] v_1751;
  wire [0:0] v_1752;
  wire [0:0] v_1753;
  wire [0:0] v_1754;
  wire [0:0] v_1755;
  wire [0:0] v_1756;
  wire [0:0] v_1757;
  wire [19:0] v_1758;
  wire [0:0] v_1759;
  wire [0:0] v_1760;
  wire [0:0] v_1761;
  wire [0:0] v_1762;
  wire [0:0] v_1763;
  wire [0:0] v_1764;
  wire [0:0] v_1765;
  wire [0:0] v_1766;
  wire [0:0] v_1767;
  wire [0:0] v_1768;
  wire [0:0] v_1769;
  wire [0:0] v_1770;
  wire [0:0] v_1771;
  wire [0:0] v_1772;
  wire [0:0] v_1773;
  wire [0:0] v_1774;
  wire [0:0] v_1775;
  wire [0:0] v_1776;
  wire [0:0] v_1777;
  wire [0:0] v_1778;
  wire [0:0] v_1779;
  wire [0:0] v_1780;
  wire [0:0] v_1781;
  wire [0:0] v_1782;
  wire [0:0] v_1783;
  wire [0:0] v_1784;
  wire [0:0] v_1785;
  wire [0:0] v_1786;
  wire [0:0] v_1787;
  wire [0:0] v_1788;
  wire [0:0] v_1789;
  wire [0:0] v_1790;
  wire [18:0] v_1791;
  wire [0:0] v_1792;
  wire [0:0] v_1793;
  wire [0:0] v_1794;
  wire [0:0] v_1795;
  wire [0:0] v_1796;
  wire [0:0] v_1797;
  wire [0:0] v_1798;
  wire [0:0] v_1799;
  wire [0:0] v_1800;
  wire [0:0] v_1801;
  wire [0:0] v_1802;
  wire [0:0] v_1803;
  wire [0:0] v_1804;
  wire [0:0] v_1805;
  wire [0:0] v_1806;
  wire [0:0] v_1807;
  wire [0:0] v_1808;
  wire [0:0] v_1809;
  wire [0:0] v_1810;
  wire [0:0] v_1811;
  wire [0:0] v_1812;
  wire [0:0] v_1813;
  wire [0:0] v_1814;
  wire [0:0] v_1815;
  wire [0:0] v_1816;
  wire [0:0] v_1817;
  wire [0:0] v_1818;
  wire [0:0] v_1819;
  wire [0:0] v_1820;
  wire [0:0] v_1821;
  wire [0:0] v_1822;
  wire [0:0] v_1823;
  wire [17:0] v_1824;
  wire [0:0] v_1825;
  wire [0:0] v_1826;
  wire [0:0] v_1827;
  wire [0:0] v_1828;
  wire [0:0] v_1829;
  wire [0:0] v_1830;
  wire [0:0] v_1831;
  wire [0:0] v_1832;
  wire [0:0] v_1833;
  wire [0:0] v_1834;
  wire [0:0] v_1835;
  wire [0:0] v_1836;
  wire [0:0] v_1837;
  wire [0:0] v_1838;
  wire [0:0] v_1839;
  wire [0:0] v_1840;
  wire [0:0] v_1841;
  wire [0:0] v_1842;
  wire [0:0] v_1843;
  wire [0:0] v_1844;
  wire [0:0] v_1845;
  wire [0:0] v_1846;
  wire [0:0] v_1847;
  wire [0:0] v_1848;
  wire [0:0] v_1849;
  wire [0:0] v_1850;
  wire [0:0] v_1851;
  wire [0:0] v_1852;
  wire [0:0] v_1853;
  wire [0:0] v_1854;
  wire [0:0] v_1855;
  wire [0:0] v_1856;
  wire [16:0] v_1857;
  wire [0:0] v_1858;
  wire [0:0] v_1859;
  wire [0:0] v_1860;
  wire [0:0] v_1861;
  wire [0:0] v_1862;
  wire [0:0] v_1863;
  wire [0:0] v_1864;
  wire [0:0] v_1865;
  wire [0:0] v_1866;
  wire [0:0] v_1867;
  wire [0:0] v_1868;
  wire [0:0] v_1869;
  wire [0:0] v_1870;
  wire [0:0] v_1871;
  wire [0:0] v_1872;
  wire [0:0] v_1873;
  wire [0:0] v_1874;
  wire [0:0] v_1875;
  wire [0:0] v_1876;
  wire [0:0] v_1877;
  wire [0:0] v_1878;
  wire [0:0] v_1879;
  wire [0:0] v_1880;
  wire [0:0] v_1881;
  wire [0:0] v_1882;
  wire [0:0] v_1883;
  wire [0:0] v_1884;
  wire [0:0] v_1885;
  wire [0:0] v_1886;
  wire [0:0] v_1887;
  wire [0:0] v_1888;
  wire [0:0] v_1889;
  wire [15:0] v_1890;
  wire [0:0] v_1891;
  wire [0:0] v_1892;
  wire [0:0] v_1893;
  wire [0:0] v_1894;
  wire [0:0] v_1895;
  wire [0:0] v_1896;
  wire [0:0] v_1897;
  wire [0:0] v_1898;
  wire [0:0] v_1899;
  wire [0:0] v_1900;
  wire [0:0] v_1901;
  wire [0:0] v_1902;
  wire [0:0] v_1903;
  wire [0:0] v_1904;
  wire [0:0] v_1905;
  wire [0:0] v_1906;
  wire [0:0] v_1907;
  wire [0:0] v_1908;
  wire [0:0] v_1909;
  wire [0:0] v_1910;
  wire [0:0] v_1911;
  wire [0:0] v_1912;
  wire [0:0] v_1913;
  wire [0:0] v_1914;
  wire [0:0] v_1915;
  wire [0:0] v_1916;
  wire [0:0] v_1917;
  wire [0:0] v_1918;
  wire [0:0] v_1919;
  wire [0:0] v_1920;
  wire [0:0] v_1921;
  wire [0:0] v_1922;
  wire [14:0] v_1923;
  wire [0:0] v_1924;
  wire [0:0] v_1925;
  wire [0:0] v_1926;
  wire [0:0] v_1927;
  wire [0:0] v_1928;
  wire [0:0] v_1929;
  wire [0:0] v_1930;
  wire [0:0] v_1931;
  wire [0:0] v_1932;
  wire [0:0] v_1933;
  wire [0:0] v_1934;
  wire [0:0] v_1935;
  wire [0:0] v_1936;
  wire [0:0] v_1937;
  wire [0:0] v_1938;
  wire [0:0] v_1939;
  wire [0:0] v_1940;
  wire [0:0] v_1941;
  wire [0:0] v_1942;
  wire [0:0] v_1943;
  wire [0:0] v_1944;
  wire [0:0] v_1945;
  wire [0:0] v_1946;
  wire [0:0] v_1947;
  wire [0:0] v_1948;
  wire [0:0] v_1949;
  wire [0:0] v_1950;
  wire [0:0] v_1951;
  wire [0:0] v_1952;
  wire [0:0] v_1953;
  wire [0:0] v_1954;
  wire [13:0] v_1955;
  wire [0:0] v_1956;
  wire [0:0] v_1957;
  wire [0:0] v_1958;
  wire [0:0] v_1959;
  wire [0:0] v_1960;
  wire [0:0] v_1961;
  wire [0:0] v_1962;
  wire [0:0] v_1963;
  wire [0:0] v_1964;
  wire [0:0] v_1965;
  wire [0:0] v_1966;
  wire [0:0] v_1967;
  wire [0:0] v_1968;
  wire [0:0] v_1969;
  wire [0:0] v_1970;
  wire [0:0] v_1971;
  wire [0:0] v_1972;
  wire [0:0] v_1973;
  wire [0:0] v_1974;
  wire [0:0] v_1975;
  wire [0:0] v_1976;
  wire [0:0] v_1977;
  wire [0:0] v_1978;
  wire [0:0] v_1979;
  wire [0:0] v_1980;
  wire [0:0] v_1981;
  wire [0:0] v_1982;
  wire [0:0] v_1983;
  wire [0:0] v_1984;
  wire [0:0] v_1985;
  wire [0:0] v_1986;
  wire [12:0] v_1987;
  wire [0:0] v_1988;
  wire [0:0] v_1989;
  wire [0:0] v_1990;
  wire [0:0] v_1991;
  wire [0:0] v_1992;
  wire [0:0] v_1993;
  wire [0:0] v_1994;
  wire [0:0] v_1995;
  wire [0:0] v_1996;
  wire [0:0] v_1997;
  wire [0:0] v_1998;
  wire [0:0] v_1999;
  wire [0:0] v_2000;
  wire [0:0] v_2001;
  wire [0:0] v_2002;
  wire [0:0] v_2003;
  wire [0:0] v_2004;
  wire [0:0] v_2005;
  wire [0:0] v_2006;
  wire [0:0] v_2007;
  wire [0:0] v_2008;
  wire [0:0] v_2009;
  wire [0:0] v_2010;
  wire [0:0] v_2011;
  wire [0:0] v_2012;
  wire [0:0] v_2013;
  wire [0:0] v_2014;
  wire [0:0] v_2015;
  wire [0:0] v_2016;
  wire [0:0] v_2017;
  wire [0:0] v_2018;
  wire [11:0] v_2019;
  wire [0:0] v_2020;
  wire [0:0] v_2021;
  wire [0:0] v_2022;
  wire [0:0] v_2023;
  wire [0:0] v_2024;
  wire [0:0] v_2025;
  wire [0:0] v_2026;
  wire [0:0] v_2027;
  wire [0:0] v_2028;
  wire [0:0] v_2029;
  wire [0:0] v_2030;
  wire [0:0] v_2031;
  wire [0:0] v_2032;
  wire [0:0] v_2033;
  wire [0:0] v_2034;
  wire [0:0] v_2035;
  wire [0:0] v_2036;
  wire [0:0] v_2037;
  wire [0:0] v_2038;
  wire [0:0] v_2039;
  wire [0:0] v_2040;
  wire [0:0] v_2041;
  wire [0:0] v_2042;
  wire [0:0] v_2043;
  wire [0:0] v_2044;
  wire [0:0] v_2045;
  wire [0:0] v_2046;
  wire [0:0] v_2047;
  wire [0:0] v_2048;
  wire [0:0] v_2049;
  wire [0:0] v_2050;
  wire [10:0] v_2051;
  wire [0:0] v_2052;
  wire [0:0] v_2053;
  wire [0:0] v_2054;
  wire [0:0] v_2055;
  wire [0:0] v_2056;
  wire [0:0] v_2057;
  wire [0:0] v_2058;
  wire [0:0] v_2059;
  wire [0:0] v_2060;
  wire [0:0] v_2061;
  wire [0:0] v_2062;
  wire [0:0] v_2063;
  wire [0:0] v_2064;
  wire [0:0] v_2065;
  wire [0:0] v_2066;
  wire [0:0] v_2067;
  wire [0:0] v_2068;
  wire [0:0] v_2069;
  wire [0:0] v_2070;
  wire [0:0] v_2071;
  wire [0:0] v_2072;
  wire [0:0] v_2073;
  wire [0:0] v_2074;
  wire [0:0] v_2075;
  wire [0:0] v_2076;
  wire [0:0] v_2077;
  wire [0:0] v_2078;
  wire [0:0] v_2079;
  wire [0:0] v_2080;
  wire [0:0] v_2081;
  wire [0:0] v_2082;
  wire [9:0] v_2083;
  wire [0:0] v_2084;
  wire [0:0] v_2085;
  wire [0:0] v_2086;
  wire [0:0] v_2087;
  wire [0:0] v_2088;
  wire [0:0] v_2089;
  wire [0:0] v_2090;
  wire [0:0] v_2091;
  wire [0:0] v_2092;
  wire [0:0] v_2093;
  wire [0:0] v_2094;
  wire [0:0] v_2095;
  wire [0:0] v_2096;
  wire [0:0] v_2097;
  wire [0:0] v_2098;
  wire [0:0] v_2099;
  wire [0:0] v_2100;
  wire [0:0] v_2101;
  wire [0:0] v_2102;
  wire [0:0] v_2103;
  wire [0:0] v_2104;
  wire [0:0] v_2105;
  wire [0:0] v_2106;
  wire [0:0] v_2107;
  wire [0:0] v_2108;
  wire [0:0] v_2109;
  wire [0:0] v_2110;
  wire [0:0] v_2111;
  wire [0:0] v_2112;
  wire [0:0] v_2113;
  wire [0:0] v_2114;
  wire [8:0] v_2115;
  wire [0:0] v_2116;
  wire [0:0] v_2117;
  wire [0:0] v_2118;
  wire [0:0] v_2119;
  wire [0:0] v_2120;
  wire [0:0] v_2121;
  wire [0:0] v_2122;
  wire [0:0] v_2123;
  wire [0:0] v_2124;
  wire [0:0] v_2125;
  wire [0:0] v_2126;
  wire [0:0] v_2127;
  wire [0:0] v_2128;
  wire [0:0] v_2129;
  wire [0:0] v_2130;
  wire [0:0] v_2131;
  wire [0:0] v_2132;
  wire [0:0] v_2133;
  wire [0:0] v_2134;
  wire [0:0] v_2135;
  wire [0:0] v_2136;
  wire [0:0] v_2137;
  wire [0:0] v_2138;
  wire [0:0] v_2139;
  wire [0:0] v_2140;
  wire [0:0] v_2141;
  wire [0:0] v_2142;
  wire [0:0] v_2143;
  wire [0:0] v_2144;
  wire [0:0] v_2145;
  wire [0:0] v_2146;
  wire [7:0] v_2147;
  wire [0:0] v_2148;
  wire [0:0] v_2149;
  wire [0:0] v_2150;
  wire [0:0] v_2151;
  wire [0:0] v_2152;
  wire [0:0] v_2153;
  wire [0:0] v_2154;
  wire [0:0] v_2155;
  wire [0:0] v_2156;
  wire [0:0] v_2157;
  wire [0:0] v_2158;
  wire [0:0] v_2159;
  wire [0:0] v_2160;
  wire [0:0] v_2161;
  wire [0:0] v_2162;
  wire [0:0] v_2163;
  wire [0:0] v_2164;
  wire [0:0] v_2165;
  wire [0:0] v_2166;
  wire [0:0] v_2167;
  wire [0:0] v_2168;
  wire [0:0] v_2169;
  wire [0:0] v_2170;
  wire [0:0] v_2171;
  wire [0:0] v_2172;
  wire [0:0] v_2173;
  wire [0:0] v_2174;
  wire [0:0] v_2175;
  wire [0:0] v_2176;
  wire [0:0] v_2177;
  wire [0:0] v_2178;
  wire [6:0] v_2179;
  wire [0:0] v_2180;
  wire [0:0] v_2181;
  wire [0:0] v_2182;
  wire [0:0] v_2183;
  wire [0:0] v_2184;
  wire [0:0] v_2185;
  wire [0:0] v_2186;
  wire [0:0] v_2187;
  wire [0:0] v_2188;
  wire [0:0] v_2189;
  wire [0:0] v_2190;
  wire [0:0] v_2191;
  wire [0:0] v_2192;
  wire [0:0] v_2193;
  wire [0:0] v_2194;
  wire [0:0] v_2195;
  wire [0:0] v_2196;
  wire [0:0] v_2197;
  wire [0:0] v_2198;
  wire [0:0] v_2199;
  wire [0:0] v_2200;
  wire [0:0] v_2201;
  wire [0:0] v_2202;
  wire [0:0] v_2203;
  wire [0:0] v_2204;
  wire [0:0] v_2205;
  wire [0:0] v_2206;
  wire [0:0] v_2207;
  wire [0:0] v_2208;
  wire [0:0] v_2209;
  wire [0:0] v_2210;
  wire [5:0] v_2211;
  wire [0:0] v_2212;
  wire [0:0] v_2213;
  wire [0:0] v_2214;
  wire [0:0] v_2215;
  wire [0:0] v_2216;
  wire [0:0] v_2217;
  wire [0:0] v_2218;
  wire [0:0] v_2219;
  wire [0:0] v_2220;
  wire [0:0] v_2221;
  wire [0:0] v_2222;
  wire [0:0] v_2223;
  wire [0:0] v_2224;
  wire [0:0] v_2225;
  wire [0:0] v_2226;
  wire [0:0] v_2227;
  wire [0:0] v_2228;
  wire [0:0] v_2229;
  wire [0:0] v_2230;
  wire [0:0] v_2231;
  wire [0:0] v_2232;
  wire [0:0] v_2233;
  wire [0:0] v_2234;
  wire [0:0] v_2235;
  wire [0:0] v_2236;
  wire [0:0] v_2237;
  wire [0:0] v_2238;
  wire [0:0] v_2239;
  wire [0:0] v_2240;
  wire [0:0] v_2241;
  wire [0:0] v_2242;
  wire [4:0] v_2243;
  wire [0:0] v_2244;
  wire [0:0] v_2245;
  wire [0:0] v_2246;
  wire [0:0] v_2247;
  wire [0:0] v_2248;
  wire [0:0] v_2249;
  wire [0:0] v_2250;
  wire [0:0] v_2251;
  wire [0:0] v_2252;
  wire [0:0] v_2253;
  wire [0:0] v_2254;
  wire [0:0] v_2255;
  wire [0:0] v_2256;
  wire [0:0] v_2257;
  wire [0:0] v_2258;
  wire [0:0] v_2259;
  wire [0:0] v_2260;
  wire [0:0] v_2261;
  wire [0:0] v_2262;
  wire [0:0] v_2263;
  wire [0:0] v_2264;
  wire [0:0] v_2265;
  wire [0:0] v_2266;
  wire [0:0] v_2267;
  wire [0:0] v_2268;
  wire [0:0] v_2269;
  wire [0:0] v_2270;
  wire [0:0] v_2271;
  wire [0:0] v_2272;
  wire [0:0] v_2273;
  wire [0:0] v_2274;
  wire [0:0] v_2275;
  wire [3:0] v_2276;
  wire [0:0] v_2277;
  wire [0:0] v_2278;
  wire [0:0] v_2279;
  wire [0:0] v_2280;
  wire [0:0] v_2281;
  wire [0:0] v_2282;
  wire [0:0] v_2283;
  wire [0:0] v_2284;
  wire [0:0] v_2285;
  wire [0:0] v_2286;
  wire [0:0] v_2287;
  wire [0:0] v_2288;
  wire [0:0] v_2289;
  wire [0:0] v_2290;
  wire [0:0] v_2291;
  wire [0:0] v_2292;
  wire [0:0] v_2293;
  wire [0:0] v_2294;
  wire [0:0] v_2295;
  wire [0:0] v_2296;
  wire [0:0] v_2297;
  wire [0:0] v_2298;
  wire [0:0] v_2299;
  wire [0:0] v_2300;
  wire [0:0] v_2301;
  wire [0:0] v_2302;
  wire [0:0] v_2303;
  wire [0:0] v_2304;
  wire [0:0] v_2305;
  wire [0:0] v_2306;
  wire [0:0] v_2307;
  wire [0:0] v_2308;
  wire [2:0] v_2309;
  wire [0:0] v_2310;
  wire [0:0] v_2311;
  wire [0:0] v_2312;
  wire [0:0] v_2313;
  wire [0:0] v_2314;
  wire [0:0] v_2315;
  wire [0:0] v_2316;
  wire [0:0] v_2317;
  wire [0:0] v_2318;
  wire [0:0] v_2319;
  wire [0:0] v_2320;
  wire [0:0] v_2321;
  wire [0:0] v_2322;
  wire [0:0] v_2323;
  wire [0:0] v_2324;
  wire [0:0] v_2325;
  wire [0:0] v_2326;
  wire [0:0] v_2327;
  wire [0:0] v_2328;
  wire [0:0] v_2329;
  wire [0:0] v_2330;
  wire [0:0] v_2331;
  wire [0:0] v_2332;
  wire [0:0] v_2333;
  wire [0:0] v_2334;
  wire [0:0] v_2335;
  wire [0:0] v_2336;
  wire [0:0] v_2337;
  wire [0:0] v_2338;
  wire [0:0] v_2339;
  wire [0:0] v_2340;
  wire [0:0] v_2341;
  wire [1:0] v_2342;
  wire [0:0] v_2343;
  wire [0:0] v_2344;
  wire [0:0] v_2345;
  wire [0:0] v_2346;
  wire [0:0] v_2347;
  wire [0:0] v_2348;
  wire [0:0] v_2349;
  wire [0:0] v_2350;
  wire [0:0] v_2351;
  wire [0:0] v_2352;
  wire [0:0] v_2353;
  wire [0:0] v_2354;
  wire [0:0] v_2355;
  wire [0:0] v_2356;
  wire [0:0] v_2357;
  wire [0:0] v_2358;
  wire [0:0] v_2359;
  wire [0:0] v_2360;
  wire [0:0] v_2361;
  wire [0:0] v_2362;
  wire [0:0] v_2363;
  wire [0:0] v_2364;
  wire [0:0] v_2365;
  wire [0:0] v_2366;
  wire [0:0] v_2367;
  wire [0:0] v_2368;
  wire [0:0] v_2369;
  wire [0:0] v_2370;
  wire [0:0] v_2371;
  wire [0:0] v_2372;
  wire [0:0] v_2373;
  wire [0:0] v_2374;
  wire [0:0] v_2375;
  wire [0:0] v_2376;
  wire [0:0] v_2377;
  wire [0:0] v_2378;
  wire [0:0] v_2379;
  wire [0:0] v_2380;
  wire [0:0] v_2381;
  wire [0:0] v_2382;
  wire [0:0] v_2383;
  wire [0:0] v_2384;
  wire [0:0] v_2385;
  wire [0:0] v_2386;
  wire [0:0] v_2387;
  wire [0:0] v_2388;
  wire [0:0] v_2389;
  wire [0:0] v_2390;
  wire [0:0] v_2391;
  wire [0:0] v_2392;
  wire [0:0] v_2393;
  wire [0:0] v_2394;
  wire [0:0] v_2395;
  wire [0:0] v_2396;
  wire [0:0] v_2397;
  wire [0:0] v_2398;
  wire [0:0] v_2399;
  wire [0:0] v_2400;
  wire [0:0] v_2401;
  wire [0:0] v_2402;
  wire [0:0] v_2403;
  wire [0:0] v_2404;
  wire [0:0] v_2405;
  wire [0:0] v_2406;
  wire [0:0] v_2407;
  wire [0:0] v_2408;
  wire [0:0] v_2409;
  wire [0:0] v_2410;
  wire [0:0] v_2411;
  wire [0:0] v_2412;
  wire [0:0] v_2413;
  wire [0:0] v_2414;
  wire [0:0] v_2415;
  wire [0:0] v_2416;
  wire [0:0] v_2417;
  wire [0:0] v_2418;
  wire [4:0] v_2419;
  wire [0:0] v_2420;
  wire [3:0] v_2421;
  wire [0:0] v_2422;
  wire [2:0] v_2423;
  wire [0:0] v_2424;
  wire [1:0] v_2425;
  wire [0:0] v_2426;
  wire [0:0] v_2427;
  wire [4:0] v_2428;
  wire [0:0] v_2429;
  wire [3:0] v_2430;
  wire [0:0] v_2431;
  wire [2:0] v_2432;
  wire [0:0] v_2433;
  wire [1:0] v_2434;
  wire [0:0] v_2435;
  wire [0:0] v_2436;
  wire [31:0] v_2437;
  function [31:0] mux_2437(input [0:0] sel);
    case (sel) 0: mux_2437 = v_2458; 1: mux_2437 = v_384;
    endcase
  endfunction
  wire [0:0] v_2438;
  wire [0:0] v_2439;
  wire [4:0] v_2440;
  wire [0:0] v_2441;
  wire [3:0] v_2442;
  wire [0:0] v_2443;
  wire [2:0] v_2444;
  wire [0:0] v_2445;
  wire [1:0] v_2446;
  wire [0:0] v_2447;
  wire [0:0] v_2448;
  wire [4:0] v_2449;
  wire [0:0] v_2450;
  wire [3:0] v_2451;
  wire [0:0] v_2452;
  wire [2:0] v_2453;
  wire [0:0] v_2454;
  wire [1:0] v_2455;
  wire [0:0] v_2456;
  wire [0:0] v_2457;
  wire [31:0] v_2458;
  function [31:0] mux_2458(input [0:0] sel);
    case (sel) 0: mux_2458 = v_2493; 1: mux_2458 = v_2512;
    endcase
  endfunction
  wire [0:0] v_2459;
  wire [0:0] v_2460;
  reg [0:0] v_2461 = 1'h0;
  reg [0:0] v_2462 = 1'h0;
  wire [0:0] v_2463;
  reg [4:0] v_2464 = 5'h0;
  wire [4:0] v_2465;
  wire [4:0] v_2466;
  function [4:0] mux_2466(input [0:0] sel);
    case (sel) 0: mux_2466 = 5'h0; 1: mux_2466 = v_2467;
    endcase
  endfunction
  wire [4:0] v_2467;
  function [4:0] mux_2467(input [0:0] sel);
    case (sel) 0: mux_2467 = v_2468; 1: mux_2467 = v_2477;
    endcase
  endfunction
  wire [4:0] v_2468;
  wire [0:0] v_2469;
  wire [3:0] v_2470;
  wire [0:0] v_2471;
  wire [2:0] v_2472;
  wire [0:0] v_2473;
  wire [1:0] v_2474;
  wire [0:0] v_2475;
  wire [0:0] v_2476;
  wire [4:0] v_2477;
  wire [0:0] v_2478;
  wire [3:0] v_2479;
  wire [0:0] v_2480;
  wire [2:0] v_2481;
  wire [0:0] v_2482;
  wire [1:0] v_2483;
  wire [0:0] v_2484;
  wire [0:0] v_2485;
  wire [4:0] v_2486;
  function [4:0] mux_2486(input [0:0] sel);
    case (sel) 0: mux_2486 = 5'h0; 1: mux_2486 = 5'bxxxxx;
    endcase
  endfunction
  wire [0:0] v_2487;
  reg [4:0] v_2488 = 5'h0;
  wire [4:0] v_2489;
  wire [4:0] v_2490;
  function [4:0] mux_2490(input [0:0] sel);
    case (sel) 0: mux_2490 = 5'h0; 1: mux_2490 = v_362;
    endcase
  endfunction
  wire [4:0] v_2491;
  function [4:0] mux_2491(input [0:0] sel);
    case (sel) 0: mux_2491 = 5'h0; 1: mux_2491 = 5'bxxxxx;
    endcase
  endfunction
  wire [0:0] v_2492;
  wire [31:0] v_2493;
  wire [4:0] v_2494;
  wire [4:0] v_2495;
  function [4:0] mux_2495(input [0:0] sel);
    case (sel) 0: mux_2495 = 5'h0; 1: mux_2495 = v_2467;
    endcase
  endfunction
  wire [4:0] v_2496;
  function [4:0] mux_2496(input [0:0] sel);
    case (sel) 0: mux_2496 = 5'h0; 1: mux_2496 = 5'bxxxxx;
    endcase
  endfunction
  wire [0:0] v_2497;
  wire [4:0] v_2498;
  wire [4:0] v_2499;
  function [4:0] mux_2499(input [0:0] sel);
    case (sel) 0: mux_2499 = 5'h0; 1: mux_2499 = v_362;
    endcase
  endfunction
  wire [4:0] v_2500;
  function [4:0] mux_2500(input [0:0] sel);
    case (sel) 0: mux_2500 = 5'h0; 1: mux_2500 = 5'bxxxxx;
    endcase
  endfunction
  wire [0:0] v_2501;
  wire [31:0] v_2502;
  wire [31:0] v_2503;
  function [31:0] mux_2503(input [0:0] sel);
    case (sel) 0: mux_2503 = 32'h0; 1: mux_2503 = v_384;
    endcase
  endfunction
  wire [31:0] v_2504;
  function [31:0] mux_2504(input [0:0] sel);
    case (sel)
      0: mux_2504 = 32'h0;
      1: mux_2504 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_2505;
  wire [0:0] v_2506;
  wire [0:0] v_2507;
  function [0:0] mux_2507(input [0:0] sel);
    case (sel) 0: mux_2507 = 1'h0; 1: mux_2507 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2508;
  function [0:0] mux_2508(input [0:0] sel);
    case (sel) 0: mux_2508 = 1'h0; 1: mux_2508 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2509;
  wire [0:0] v_2510;
  function [0:0] mux_2510(input [0:0] sel);
    case (sel) 0: mux_2510 = 1'h0; 1: mux_2510 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2511;
  reg [31:0] v_2512 = 32'h0;
  wire [31:0] v_2513;
  wire [31:0] v_2514;
  function [31:0] mux_2514(input [0:0] sel);
    case (sel) 0: mux_2514 = 32'h0; 1: mux_2514 = v_384;
    endcase
  endfunction
  wire [31:0] v_2515;
  function [31:0] mux_2515(input [0:0] sel);
    case (sel)
      0: mux_2515 = 32'h0;
      1: mux_2515 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_2516;
  wire [0:0] v_2517;
  wire [0:0] v_2518;
  reg [0:0] v_2519 = 1'h0;
  wire [0:0] v_2520;
  wire [0:0] v_2521;
  wire [0:0] v_2522;
  wire [0:0] v_2523;
  wire [0:0] v_2524;
  wire [0:0] v_2525;
  reg [0:0] v_2526 = 1'h0;
  wire [0:0] v_2527;
  wire [0:0] v_2528;
  wire [0:0] v_2529;
  wire [0:0] v_2530;
  wire [0:0] v_2531;
  wire [0:0] v_2532;
  wire [0:0] v_2533;
  reg [0:0] v_2534 = 1'h0;
  wire [0:0] v_2535;
  wire [0:0] v_2536;
  wire [0:0] v_2537;
  wire [0:0] v_2538;
  wire [0:0] v_2539;
  wire [0:0] v_2540;
  wire [0:0] v_2541;
  wire [31:0] v_2542;
  wire [31:0] v_2543;
  reg [0:0] v_2544 = 1'h0;
  wire [30:0] v_2545;
  wire [29:0] v_2546;
  wire [28:0] v_2547;
  wire [27:0] v_2548;
  wire [26:0] v_2549;
  wire [25:0] v_2550;
  wire [24:0] v_2551;
  wire [23:0] v_2552;
  wire [22:0] v_2553;
  wire [21:0] v_2554;
  wire [20:0] v_2555;
  wire [19:0] v_2556;
  wire [18:0] v_2557;
  wire [17:0] v_2558;
  wire [16:0] v_2559;
  wire [15:0] v_2560;
  wire [14:0] v_2561;
  wire [13:0] v_2562;
  wire [12:0] v_2563;
  wire [11:0] v_2564;
  reg [0:0] v_2565 = 1'h0;
  wire [10:0] v_2566;
  reg [0:0] v_2567 = 1'h0;
  wire [9:0] v_2568;
  reg [0:0] v_2569 = 1'h0;
  wire [8:0] v_2570;
  reg [0:0] v_2571 = 1'h0;
  wire [7:0] v_2572;
  reg [0:0] v_2573 = 1'h0;
  wire [6:0] v_2574;
  reg [0:0] v_2575 = 1'h0;
  wire [5:0] v_2576;
  reg [0:0] v_2577 = 1'h0;
  wire [4:0] v_2578;
  reg [0:0] v_2579 = 1'h0;
  wire [3:0] v_2580;
  reg [0:0] v_2581 = 1'h0;
  wire [2:0] v_2582;
  reg [0:0] v_2583 = 1'h0;
  wire [1:0] v_2584;
  reg [0:0] v_2585 = 1'h0;
  reg [0:0] v_2586 = 1'h0;
  wire [31:0] v_2587;
  function [31:0] mux_2587(input [0:0] sel);
    case (sel)
      0: mux_2587 = 32'h0;
      1: mux_2587 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_2588;
  wire [31:0] v_2589;
  wire [31:0] v_2590;
  wire [31:0] v_2591;
  function [31:0] mux_2591(input [0:0] sel);
    case (sel) 0: mux_2591 = 32'h0; 1: mux_2591 = v_792;
    endcase
  endfunction
  wire [31:0] v_2592;
  function [31:0] mux_2592(input [0:0] sel);
    case (sel) 0: mux_2592 = 32'h0; 1: mux_2592 = v_792;
    endcase
  endfunction
  wire [31:0] v_2593;
  wire [31:0] v_2594;
  function [31:0] mux_2594(input [0:0] sel);
    case (sel) 0: mux_2594 = 32'h0; 1: mux_2594 = v_2595;
    endcase
  endfunction
  wire [31:0] v_2595;
  wire [30:0] v_2596;
  wire [31:0] v_2597;
  wire [31:0] v_2598;
  function [31:0] mux_2598(input [0:0] sel);
    case (sel) 0: mux_2598 = 32'h0; 1: mux_2598 = v_2601;
    endcase
  endfunction
  wire [0:0] v_2599;
  wire [0:0] v_2600;
  wire [31:0] v_2601;
  wire [8:0] v_2602;
  function [8:0] mux_2602(input [0:0] sel);
    case (sel) 0: mux_2602 = 9'h0; 1: mux_2602 = 9'bxxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_2603;
  wire [31:0] v_2604;
  function [31:0] mux_2604(input [0:0] sel);
    case (sel)
      0: mux_2604 = 32'h0;
      1: mux_2604 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_2605;
  wire [0:0] v_2606;
  function [0:0] mux_2606(input [0:0] sel);
    case (sel) 0: mux_2606 = 1'h0; 1: mux_2606 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2607;
  wire [0:0] v_2608;
  wire [0:0] v_2609;
  function [0:0] mux_2609(input [0:0] sel);
    case (sel) 0: mux_2609 = 1'h0; 1: mux_2609 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2610;
  wire [0:0] v_2611;
  function [0:0] mux_2611(input [0:0] sel);
    case (sel) 0: mux_2611 = 1'h0; 1: mux_2611 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2612;
  wire [0:0] v_2613;
  wire [0:0] v_2614;
  wire [0:0] v_2615;
  wire [0:0] v_2616;
  wire [0:0] v_2617;
  wire [0:0] v_2618;
  wire [0:0] v_2619;
  wire [0:0] v_2620;
  wire [0:0] v_2621;
  wire [0:0] v_2622;
  function [0:0] mux_2622(input [0:0] sel);
    case (sel) 0: mux_2622 = 1'h0; 1: mux_2622 = v_2623;
    endcase
  endfunction
  reg [0:0] v_2623 = 1'h0;
  wire [0:0] v_2624;
  function [0:0] mux_2624(input [0:0] sel);
    case (sel) 0: mux_2624 = 1'h0; 1: mux_2624 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2625;
  wire [0:0] v_2626;
  function [0:0] mux_2626(input [0:0] sel);
    case (sel) 0: mux_2626 = 1'h0; 1: mux_2626 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2627;
  reg [0:0] v_2628 = 1'h0;
  wire [0:0] v_2629;
  function [0:0] mux_2629(input [0:0] sel);
    case (sel) 0: mux_2629 = 1'h0; 1: mux_2629 = 1'bx;
    endcase
  endfunction
  wire [0:0] v_2630;
  wire [0:0] v_2631;
  wire [0:0] v_2632;
  wire [0:0] v_2633;
  function [0:0] mux_2633(input [0:0] sel);
    case (sel) 0: mux_2633 = 1'h0; 1: mux_2633 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2634;
  function [0:0] mux_2634(input [0:0] sel);
    case (sel) 0: mux_2634 = 1'h0; 1: mux_2634 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2635;
  wire [0:0] v_2636;
  wire [0:0] v_2637;
  wire [0:0] v_2638;
  wire [0:0] v_2639;
  wire [0:0] v_2640;
  wire [0:0] v_2641;
  function [0:0] mux_2641(input [0:0] sel);
    case (sel) 0: mux_2641 = 1'h0; 1: mux_2641 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2642;
  function [0:0] mux_2642(input [0:0] sel);
    case (sel) 0: mux_2642 = 1'h0; 1: mux_2642 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2643;
  wire [0:0] v_2644;
  function [0:0] mux_2644(input [0:0] sel);
    case (sel) 0: mux_2644 = 1'h0; 1: mux_2644 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2645;
  function [0:0] mux_2645(input [0:0] sel);
    case (sel) 0: mux_2645 = 1'h0; 1: mux_2645 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2646;
  wire [0:0] v_2647;
  wire [0:0] v_2648;
  function [0:0] mux_2648(input [0:0] sel);
    case (sel) 0: mux_2648 = 1'h0; 1: mux_2648 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2649;
  wire [0:0] v_2650;
  function [0:0] mux_2650(input [0:0] sel);
    case (sel) 0: mux_2650 = 1'h0; 1: mux_2650 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2651;
  function [0:0] mux_2651(input [0:0] sel);
    case (sel) 0: mux_2651 = 1'h0; 1: mux_2651 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2652;
  wire [0:0] v_2653;
  wire [0:0] v_2654;
  function [0:0] mux_2654(input [0:0] sel);
    case (sel) 0: mux_2654 = 1'h0; 1: mux_2654 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2655;
  function [0:0] mux_2655(input [0:0] sel);
    case (sel) 0: mux_2655 = 1'h0; 1: mux_2655 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2656;
  wire [0:0] v_2657;
  function [0:0] mux_2657(input [0:0] sel);
    case (sel) 0: mux_2657 = 1'h0; 1: mux_2657 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2658;
  function [0:0] mux_2658(input [0:0] sel);
    case (sel) 0: mux_2658 = 1'h0; 1: mux_2658 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2659;
  wire [0:0] v_2660;
  wire [0:0] v_2661;
  wire [0:0] v_2662;
  wire [0:0] v_2663;
  wire [0:0] v_2664;
  wire [0:0] v_2665;
  wire [0:0] v_2667;
  wire [0:0] v_2668;
  reg [31:0] v_2669 = 32'h0;
  wire [31:0] v_2670;
  wire [0:0] v_2672;
  wire [0:0] v_2673;
  wire [0:0] v_2675;
  wire [0:0] v_2676;
  function [0:0] mux_2676(input [0:0] sel);
    case (sel) 0: mux_2676 = 1'h0; 1: mux_2676 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2677;
  function [0:0] mux_2677(input [0:0] sel);
    case (sel) 0: mux_2677 = 1'h0; 1: mux_2677 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2678;
  reg [7:0] v_2681 = 8'h0;
  wire [7:0] v_2682;
  wire [7:0] v_2683;
  function [7:0] mux_2683(input [0:0] sel);
    case (sel) 0: mux_2683 = 8'h0; 1: mux_2683 = v_2684;
    endcase
  endfunction
  wire [7:0] v_2684;
  wire [7:0] v_2685;
  function [7:0] mux_2685(input [0:0] sel);
    case (sel) 0: mux_2685 = 8'h0; 1: mux_2685 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_2686;
  // Instances
  //////////////////////////////////////////////////////////////////////////////
  assign v_1 = v_2 & 1'h1;
  assign v_2 = v_3 & act_35;
  assign v_3 = v_4 | v_2652;
  assign v_4 = v_5 | v_2649;
  assign v_5 = v_6 | v_2648;
  assign v_6 = mux_6(v_7);
  assign v_7 = v_8 & v_2646;
  assign v_9 = v_10 | v_2636;
  assign v_10 = v_11 | v_25;
  assign v_11 = 1'h1 & v_12;
  assign v_12 = v_13 | v_2635;
  assign v_14 = v_15 | v_16;
  assign v_15 = v_11 & v_13;
  assign v_16 = v_17 & 1'h1;
  assign v_17 = v_18 & v_2631;
  assign v_18 = v_19 | v_2629;
  assign v_19 = mux_19(1'h1);
  assign v_20 = v_21 | v_2628;
  assign v_23 = v_24 | v_2626;
  assign v_24 = mux_24(v_25);
  assign v_25 = v_26 & v_419;
  assign v_26 = v_27 & v_411;
  assign v_27 = v_28 | 1'h0;
  assign v_30 = v_31 | v_2620;
  assign v_31 = v_32 & v_33;
  assign v_32 = ~v_3;
  assign v_33 = 1'h1 & v_34;
  assign v_34 = ~act_35;
  assign act_35 = v_36 | v_2618;
  assign v_36 = v_37 | v_2599;
  assign v_37 = v_38 & v_411;
  assign v_38 = v_39 | 1'h0;
  assign v_40 = v_41 & v_2617;
  assign v_41 = v_42 & v_85;
  assign v_42 = v_43 & v_84;
  assign v_43 = v_44 & v_2616;
  assign v_44 = v_45 & v_2615;
  assign v_45 = v_46 & v_2614;
  assign v_46 = v_47 & v_79;
  assign v_47 = v_48 & v_2613;
  assign v_48 = v_49 & v_137;
  assign v_49 = 1'h1 & v_50;
  assign v_50 = v_51[1:1];
  BlockRAM# (.INIT_FILE("prog.mif"), .ADDR_WIDTH(9), .DATA_WIDTH(32))
    ram52
      (.CLK(clock),
       .ADDR(v_53),
       .DI(v_2604),
       .WE(v_2606),
       .RE(v_2608),
       .DO(v_52));
  assign v_53 = v_54 | v_2602;
  assign v_54 = mux_54(1'h1);
  assign v_55 = v_56[8:0];
  assign v_56 = v_57[31:2];
  assign v_57 = mux_57(act_35);
  assign v_58 = v_59 + 32'h4;
  assign v_60 = 1'h1 & v_61;
  assign v_61 = ~v_3;
  assign v_62 = v_63 | v_2589;
  assign v_63 = v_64 | v_2587;
  assign v_64 = mux_64(v_65);
  assign v_65 = v_66 & v_411;
  assign v_66 = v_67 | v_2523;
  assign v_67 = v_68 | v_2517;
  assign v_68 = v_69 & v_90;
  assign v_69 = v_70 | 1'h0;
  assign v_71 = v_72 & v_88;
  assign v_72 = v_73 & v_86;
  assign v_73 = v_74 & v_85;
  assign v_74 = v_75 & v_84;
  assign v_75 = v_76 & v_82;
  assign v_76 = v_77 & v_80;
  assign v_77 = v_47 & v_78;
  assign v_78 = ~v_79;
  assign v_79 = v_51[2:2];
  assign v_80 = ~v_81;
  assign v_81 = v_51[14:14];
  assign v_82 = ~v_83;
  assign v_83 = v_51[13:13];
  assign v_84 = v_51[6:6];
  assign v_85 = v_51[5:5];
  assign v_86 = ~v_87;
  assign v_87 = v_51[12:12];
  assign v_88 = ~v_89;
  assign v_89 = v_51[4:4];
  assign v_90 = v_91 == v_115;
  assign v_92 = v_93 & 1'h1;
  assign v_93 = ~v_3;
  assign v_94 = mux_94(v_95);
  assign v_95 = act_96 & v_2418;
  assign act_96 = v_97 | v_2411;
  assign v_97 = v_98 | v_2408;
  assign v_98 = v_99 | v_2407;
  assign v_99 = v_100 | v_1067;
  assign v_100 = v_101 & v_112;
  assign v_101 = v_102 != 5'h0;
  assign v_102 = {v_103, v_105};
  assign v_103 = v_104[11:11];
  assign v_105 = {v_106, v_107};
  assign v_106 = v_104[10:10];
  assign v_107 = {v_108, v_109};
  assign v_108 = v_104[9:9];
  assign v_109 = {v_110, v_111};
  assign v_110 = v_104[8:8];
  assign v_111 = v_104[7:7];
  assign v_112 = v_113 & v_408;
  assign v_113 = v_114 == 12'h805;
  assign v_114 = v_115[11:0];
  assign v_116 = mux_116(v_117);
  assign v_117 = v_118 | v_205;
  assign v_118 = v_119 | v_151;
  assign v_119 = v_120 | v_138;
  assign v_120 = v_121 | v_123;
  assign v_121 = v_122 & v_89;
  assign v_122 = v_73 & v_87;
  assign v_123 = v_124 & v_137;
  assign v_124 = v_125 & v_50;
  assign v_125 = v_126 & v_136;
  assign v_126 = v_127 & v_134;
  assign v_127 = v_128 & v_133;
  assign v_128 = v_129 & v_85;
  assign v_129 = v_130 & v_132;
  assign v_130 = 1'h1 & v_131;
  assign v_131 = ~v_81;
  assign v_132 = ~v_84;
  assign v_133 = ~v_89;
  assign v_134 = ~v_135;
  assign v_135 = v_51[3:3];
  assign v_136 = ~v_79;
  assign v_137 = v_51[0:0];
  assign v_138 = v_139 | v_40;
  assign v_139 = v_140 & v_150;
  assign v_140 = v_141 & v_149;
  assign v_141 = v_142 & v_148;
  assign v_142 = v_143 & v_147;
  assign v_143 = v_144 & v_146;
  assign v_144 = v_145 & v_137;
  assign v_145 = 1'h1 & v_50;
  assign v_146 = ~v_84;
  assign v_147 = ~v_135;
  assign v_148 = ~v_85;
  assign v_149 = ~v_89;
  assign v_150 = ~v_79;
  assign v_151 = v_152 | v_194;
  assign v_152 = v_153 | v_159;
  assign v_153 = v_154 & v_79;
  assign v_154 = v_155 & v_135;
  assign v_155 = v_156 & v_158;
  assign v_156 = v_157 & v_85;
  assign v_157 = v_144 & v_84;
  assign v_158 = ~v_89;
  assign v_159 = v_160 & v_193;
  assign v_160 = v_161 & v_87;
  assign v_161 = v_162 & v_81;
  assign v_162 = v_163 & v_192;
  assign v_163 = v_164 & v_191;
  assign v_164 = v_165 & v_137;
  assign v_165 = v_166 & v_50;
  assign v_166 = v_167 & v_190;
  assign v_167 = v_168 & v_189;
  assign v_168 = v_169 & v_89;
  assign v_169 = v_170 & v_188;
  assign v_170 = v_171 & v_186;
  assign v_171 = v_172 & v_184;
  assign v_172 = v_173 & v_182;
  assign v_173 = v_174 & v_180;
  assign v_174 = v_175 & v_178;
  assign v_175 = 1'h1 & v_176;
  assign v_176 = ~v_177;
  assign v_177 = v_51[31:31];
  assign v_178 = ~v_179;
  assign v_179 = v_51[29:29];
  assign v_180 = ~v_181;
  assign v_181 = v_51[28:28];
  assign v_182 = ~v_183;
  assign v_183 = v_51[27:27];
  assign v_184 = ~v_185;
  assign v_185 = v_51[26:26];
  assign v_186 = ~v_187;
  assign v_187 = v_51[25:25];
  assign v_188 = ~v_84;
  assign v_189 = ~v_135;
  assign v_190 = ~v_79;
  assign v_191 = v_51[30:30];
  assign v_192 = ~v_83;
  assign v_193 = ~v_85;
  assign v_194 = v_195 | v_203;
  assign v_195 = v_196 & v_81;
  assign v_196 = v_197 & v_87;
  assign v_197 = v_198 & v_202;
  assign v_198 = v_199 & v_201;
  assign v_199 = v_164 & v_200;
  assign v_200 = ~v_191;
  assign v_201 = ~v_85;
  assign v_202 = ~v_83;
  assign v_203 = v_196 & v_204;
  assign v_204 = ~v_81;
  assign v_205 = v_206 | v_240;
  assign v_206 = v_207 | v_226;
  assign v_207 = v_208 | v_218;
  assign v_208 = v_209 & v_89;
  assign v_209 = v_210 & v_217;
  assign v_210 = v_211 & v_216;
  assign v_211 = v_212 & v_215;
  assign v_212 = v_213 & v_214;
  assign v_213 = v_77 & v_81;
  assign v_214 = ~v_83;
  assign v_215 = ~v_87;
  assign v_216 = ~v_84;
  assign v_217 = ~v_85;
  assign v_218 = v_219 & v_89;
  assign v_219 = v_220 & v_225;
  assign v_220 = v_221 & v_224;
  assign v_221 = v_222 & v_223;
  assign v_222 = v_213 & v_83;
  assign v_223 = ~v_87;
  assign v_224 = ~v_84;
  assign v_225 = ~v_85;
  assign v_226 = v_227 | v_233;
  assign v_227 = v_228 & v_89;
  assign v_228 = v_229 & v_232;
  assign v_229 = v_230 & v_231;
  assign v_230 = v_222 & v_87;
  assign v_231 = ~v_84;
  assign v_232 = ~v_85;
  assign v_233 = v_234 & v_87;
  assign v_234 = v_235 & v_89;
  assign v_235 = v_236 & v_239;
  assign v_236 = v_237 & v_238;
  assign v_237 = v_76 & v_83;
  assign v_238 = ~v_84;
  assign v_239 = ~v_85;
  assign v_240 = v_241 | v_251;
  assign v_241 = v_242 | v_244;
  assign v_242 = v_234 & v_243;
  assign v_243 = ~v_87;
  assign v_244 = v_245 & v_89;
  assign v_245 = v_246 & v_250;
  assign v_246 = v_247 & v_249;
  assign v_247 = v_75 & v_248;
  assign v_248 = ~v_84;
  assign v_249 = ~v_87;
  assign v_250 = ~v_85;
  assign v_251 = v_252 | v_254;
  assign v_252 = v_253 & v_79;
  assign v_253 = v_141 & v_89;
  assign v_254 = v_255 & v_79;
  assign v_255 = v_256 & v_89;
  assign v_256 = v_142 & v_85;
  assign v_257 = mux_257(v_258);
  assign v_258 = act_96 & v_259;
  assign v_259 = v_260 == v_269;
  assign v_260 = {v_261, v_262};
  assign v_261 = v_104[11:11];
  assign v_262 = {v_263, v_264};
  assign v_263 = v_104[10:10];
  assign v_264 = {v_265, v_266};
  assign v_265 = v_104[9:9];
  assign v_266 = {v_267, v_268};
  assign v_267 = v_104[8:8];
  assign v_268 = v_104[7:7];
  assign v_269 = {v_270, v_271};
  assign v_270 = v_51[24:24];
  assign v_271 = {v_272, v_273};
  assign v_272 = v_51[23:23];
  assign v_273 = {v_274, v_275};
  assign v_274 = v_51[22:22];
  assign v_275 = {v_276, v_277};
  assign v_276 = v_51[21:21];
  assign v_277 = v_51[20:20];
  assign v_278 = mux_278(v_279);
  assign v_279 = act_280 & v_309;
  assign act_280 = v_281 | v_308;
  assign v_281 = v_282 & 1'h1;
  assign v_282 = v_283 & v_307;
  assign v_283 = ~act_284;
  assign act_284 = v_285 & v_11;
  assign v_285 = v_286 != 5'h0;
  assign v_286 = {v_287, v_300};
  assign v_287 = v_288[11:11];
  assign v_289 = v_290 & 1'h1;
  assign v_291 = v_292 | v_294;
  assign v_292 = 1'h1 & v_293;
  assign v_293 = ~act_35;
  assign v_294 = 1'h1 & act_35;
  assign v_295 = v_296 | v_299;
  assign v_296 = mux_296(v_292);
  assign v_297 = v_29 & v_298;
  assign v_298 = ~v_3;
  assign v_299 = mux_299(v_294);
  assign v_300 = {v_301, v_302};
  assign v_301 = v_288[10:10];
  assign v_302 = {v_303, v_304};
  assign v_303 = v_288[9:9];
  assign v_304 = {v_305, v_306};
  assign v_305 = v_288[8:8];
  assign v_306 = v_288[7:7];
  assign v_308 = act_284 & 1'h1;
  assign v_309 = v_310 == v_319;
  assign v_310 = {v_311, v_312};
  assign v_311 = v_288[11:11];
  assign v_312 = {v_313, v_314};
  assign v_313 = v_288[10:10];
  assign v_314 = {v_315, v_316};
  assign v_315 = v_288[9:9];
  assign v_316 = {v_317, v_318};
  assign v_317 = v_288[8:8];
  assign v_318 = v_288[7:7];
  assign v_319 = {v_320, v_321};
  assign v_320 = v_51[24:24];
  assign v_321 = {v_322, v_323};
  assign v_322 = v_51[23:23];
  assign v_323 = {v_324, v_325};
  assign v_324 = v_51[22:22];
  assign v_325 = {v_326, v_327};
  assign v_326 = v_51[21:21];
  assign v_327 = v_51[20:20];
  assign v_328 = mux_328(v_329);
  assign v_329 = v_330 & v_334;
  assign v_330 = v_331 & v_332;
  assign act_333 = act_280 & 1'h1;
  assign v_334 = v_335 == v_359;
  assign v_336 = v_337 | v_357;
  assign v_337 = mux_337(1'h1);
  assign v_338 = mux_338(v_3);
  assign v_339 = {v_340, v_341};
  assign v_340 = v_52[24:24];
  assign v_341 = {v_342, v_343};
  assign v_342 = v_52[23:23];
  assign v_343 = {v_344, v_345};
  assign v_344 = v_52[22:22];
  assign v_345 = {v_346, v_347};
  assign v_346 = v_52[21:21];
  assign v_347 = v_52[20:20];
  assign v_348 = {v_349, v_350};
  assign v_349 = v_51[24:24];
  assign v_350 = {v_351, v_352};
  assign v_351 = v_51[23:23];
  assign v_352 = {v_353, v_354};
  assign v_353 = v_51[22:22];
  assign v_354 = {v_355, v_356};
  assign v_355 = v_51[21:21];
  assign v_356 = v_51[20:20];
  assign v_357 = mux_357(v_358);
  assign v_358 = ~1'h1;
  assign v_360 = v_361 | v_371;
  assign v_361 = mux_361(act_333);
  assign v_362 = {v_363, v_364};
  assign v_363 = v_288[11:11];
  assign v_364 = {v_365, v_366};
  assign v_365 = v_288[10:10];
  assign v_366 = {v_367, v_368};
  assign v_367 = v_288[9:9];
  assign v_368 = {v_369, v_370};
  assign v_369 = v_288[8:8];
  assign v_370 = v_288[7:7];
  assign v_371 = mux_371(v_372);
  assign v_372 = ~act_333;
  BlockRAMDual#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(5), .DATA_WIDTH(32))
    ram373
      (.CLK(clock),
       .RD_ADDR(v_374),
       .WR_ADDR(v_378),
       .DI(v_382),
       .WE(v_1363),
       .RE(v_1367),
       .DO(v_373));
  assign v_374 = v_375 | v_376;
  assign v_375 = mux_375(1'h1);
  assign v_376 = mux_376(v_377);
  assign v_377 = ~1'h1;
  assign v_378 = v_379 | v_380;
  assign v_379 = mux_379(act_333);
  assign v_380 = mux_380(v_381);
  assign v_381 = ~act_333;
  assign v_382 = v_383 | v_1361;
  assign v_383 = mux_383(act_333);
  assign v_384 = v_385 | v_387;
  assign v_385 = mux_385(v_386);
  assign v_386 = ~act_280;
  assign v_387 = v_388 | v_1082;
  assign v_388 = mux_388(v_281);
  assign v_390 = v_391 | v_905;
  assign v_391 = v_392 | v_812;
  assign v_392 = v_393 | v_777;
  assign v_393 = v_394 | v_700;
  assign v_394 = mux_394(v_395);
  assign v_395 = v_396 & v_406;
  assign v_396 = v_397 != 5'h0;
  assign v_397 = {v_398, v_399};
  assign v_398 = v_104[11:11];
  assign v_399 = {v_400, v_401};
  assign v_400 = v_104[10:10];
  assign v_401 = {v_402, v_403};
  assign v_402 = v_104[9:9];
  assign v_403 = {v_404, v_405};
  assign v_404 = v_104[8:8];
  assign v_405 = v_104[7:7];
  assign v_406 = v_407 & v_408;
  assign v_407 = v_114 == 12'h802;
  assign v_408 = v_409 & v_411;
  assign v_409 = v_410 | 1'h0;
  assign v_411 = v_412 & 1'h1;
  assign v_412 = v_290 | v_413;
  assign v_414 = v_415 | v_669;
  assign v_415 = v_416 | v_666;
  assign v_416 = mux_416(v_417);
  assign v_417 = v_26 & v_418;
  assign v_418 = ~v_419;
  assign v_419 = ~v_420;
  assign v_421 = v_422 | v_634;
  assign v_422 = v_423 & v_425;
  assign v_423 = v_11 & v_424;
  assign v_424 = ~v_13;
  assign v_425 = ~v_426;
  assign v_427 = v_428 | v_435;
  assign v_428 = v_426 & v_429;
  assign v_429 = ~v_430;
  assign v_430 = v_431 | v_433;
  assign v_431 = mux_431(v_432);
  assign v_432 = v_423 & v_426;
  assign v_433 = mux_433(v_434);
  assign v_434 = ~v_432;
  assign v_435 = act_436 & v_443;
  assign act_436 = v_437 & v_442;
  assign v_437 = v_438 & v_411;
  assign v_438 = v_439 | v_440;
  assign v_440 = v_441 | 1'h0;
  assign v_442 = ~v_428;
  assign v_443 = ~v_444;
  assign v_444 = v_445[32:32];
  assign v_445 = v_446[32:0];
  assign v_446 = v_447[77:39];
  assign v_447 = {v_448, v_624};
  assign v_448 = {v_449, v_620};
  assign v_449 = v_450[38:33];
  assign v_450 = v_451[77:39];
  assign v_451 = v_452 | v_564;
  assign v_452 = {v_453, v_554};
  assign v_453 = {v_454, v_550};
  assign v_454 = v_455[38:33];
  assign v_455 = v_456[77:39];
  assign v_456 = mux_456(act_436);
  assign v_457 = {v_458, v_465};
  assign v_458 = {v_459, v_461};
  assign v_459 = v_460[38:33];
  assign v_460 = 39'h0;
  assign v_461 = {v_462, v_464};
  assign v_462 = v_463[32:32];
  assign v_463 = v_460[32:0];
  assign v_464 = v_463[31:0];
  assign v_465 = {v_466, v_471};
  assign v_466 = {v_467, v_470};
  assign v_467 = v_468[35:32];
  assign v_468 = v_469[38:3];
  assign v_469 = 39'h0;
  assign v_470 = v_468[31:0];
  assign v_471 = {v_472, v_474};
  assign v_472 = v_473[2:1];
  assign v_473 = v_469[2:0];
  assign v_474 = v_473[0:0];
  assign v_475 = {v_476, v_540};
  assign v_476 = {v_477, v_536};
  assign v_477 = v_478[38:33];
  assign v_478 = v_479[77:39];
  assign v_479 = {v_480, v_484};
  assign v_480 = {6'bxxxxxx, v_481};
  assign v_481 = {v_482, v_483};
  assign v_482 = v_441 | 1'h0;
  assign v_483 = v_91 + v_115;
  assign v_484 = {v_485, v_534};
  assign v_485 = {v_486, v_512};
  assign v_486 = v_487 | v_500;
  assign v_487 = mux_487(v_488);
  assign v_488 = v_489 == 2'h0;
  assign v_489 = {v_490, v_491};
  assign v_492 = {v_493, v_495};
  assign v_493 = v_494 == 2'h3;
  assign v_494 = v_483[1:0];
  assign v_495 = {v_496, v_497};
  assign v_496 = v_494 == 2'h2;
  assign v_497 = {v_498, v_499};
  assign v_498 = v_494 == 2'h1;
  assign v_499 = v_494 == 2'h0;
  assign v_500 = v_501 | v_503;
  assign v_501 = mux_501(v_502);
  assign v_502 = v_489 == 2'h2;
  assign v_503 = mux_503(v_504);
  assign v_504 = v_489 == 2'h1;
  assign v_505 = {v_506, v_507};
  assign v_506 = v_494 == 2'h2;
  assign v_507 = {v_508, v_509};
  assign v_508 = v_494 == 2'h2;
  assign v_509 = {v_510, v_511};
  assign v_510 = v_494 == 2'h0;
  assign v_511 = v_494 == 2'h0;
  assign v_512 = v_513 | v_520;
  assign v_513 = mux_513(v_514);
  assign v_514 = v_489 == 2'h0;
  assign v_515 = {v_516, v_518};
  assign v_516 = v_517[7:0];
  assign v_518 = {v_516, v_519};
  assign v_519 = {v_516, v_516};
  assign v_520 = v_521 | v_529;
  assign v_521 = mux_521(v_522);
  assign v_522 = v_489 == 2'h2;
  assign v_523 = {v_524, v_525};
  assign v_524 = v_517[31:24];
  assign v_525 = {v_526, v_527};
  assign v_526 = v_517[23:16];
  assign v_527 = {v_528, v_516};
  assign v_528 = v_517[15:8];
  assign v_529 = mux_529(v_530);
  assign v_530 = v_489 == 2'h1;
  assign v_531 = {v_528, v_532};
  assign v_532 = {v_516, v_533};
  assign v_533 = {v_528, v_516};
  assign v_534 = {v_489, v_535};
  assign v_536 = {v_537, v_539};
  assign v_537 = v_538[32:32];
  assign v_538 = v_478[32:0];
  assign v_539 = v_538[31:0];
  assign v_540 = {v_541, v_546};
  assign v_541 = {v_542, v_545};
  assign v_542 = v_543[35:32];
  assign v_543 = v_544[38:3];
  assign v_544 = v_479[38:0];
  assign v_545 = v_543[31:0];
  assign v_546 = {v_547, v_549};
  assign v_547 = v_548[2:1];
  assign v_548 = v_544[2:0];
  assign v_549 = v_548[0:0];
  assign v_550 = {v_551, v_553};
  assign v_551 = v_552[32:32];
  assign v_552 = v_455[32:0];
  assign v_553 = v_552[31:0];
  assign v_554 = {v_555, v_560};
  assign v_555 = {v_556, v_559};
  assign v_556 = v_557[35:32];
  assign v_557 = v_558[38:3];
  assign v_558 = v_456[38:0];
  assign v_559 = v_557[31:0];
  assign v_560 = {v_561, v_563};
  assign v_561 = v_562[2:1];
  assign v_562 = v_558[2:0];
  assign v_563 = v_562[0:0];
  assign v_564 = {v_565, v_610};
  assign v_565 = {v_566, v_606};
  assign v_566 = v_567[38:33];
  assign v_567 = v_568[77:39];
  assign v_568 = mux_568(v_569);
  assign v_569 = ~act_436;
  assign v_570 = {v_571, v_578};
  assign v_571 = {v_572, v_574};
  assign v_572 = v_573[38:33];
  assign v_573 = 39'h0;
  assign v_574 = {v_575, v_577};
  assign v_575 = v_576[32:32];
  assign v_576 = v_573[32:0];
  assign v_577 = v_576[31:0];
  assign v_578 = {v_579, v_584};
  assign v_579 = {v_580, v_583};
  assign v_580 = v_581[35:32];
  assign v_581 = v_582[38:3];
  assign v_582 = 39'h0;
  assign v_583 = v_581[31:0];
  assign v_584 = {v_585, v_587};
  assign v_585 = v_586[2:1];
  assign v_586 = v_582[2:0];
  assign v_587 = v_586[0:0];
  assign v_588 = {v_589, v_596};
  assign v_589 = {v_590, v_592};
  assign v_590 = v_591[38:33];
  assign v_591 = 39'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  assign v_592 = {v_593, v_595};
  assign v_593 = v_594[32:32];
  assign v_594 = v_591[32:0];
  assign v_595 = v_594[31:0];
  assign v_596 = {v_597, v_602};
  assign v_597 = {v_598, v_601};
  assign v_598 = v_599[35:32];
  assign v_599 = v_600[38:3];
  assign v_600 = 39'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  assign v_601 = v_599[31:0];
  assign v_602 = {v_603, v_605};
  assign v_603 = v_604[2:1];
  assign v_604 = v_600[2:0];
  assign v_605 = v_604[0:0];
  assign v_606 = {v_607, v_609};
  assign v_607 = v_608[32:32];
  assign v_608 = v_567[32:0];
  assign v_609 = v_608[31:0];
  assign v_610 = {v_611, v_616};
  assign v_611 = {v_612, v_615};
  assign v_612 = v_613[35:32];
  assign v_613 = v_614[38:3];
  assign v_614 = v_568[38:0];
  assign v_615 = v_613[31:0];
  assign v_616 = {v_617, v_619};
  assign v_617 = v_618[2:1];
  assign v_618 = v_614[2:0];
  assign v_619 = v_618[0:0];
  assign v_620 = {v_621, v_623};
  assign v_621 = v_622[32:32];
  assign v_622 = v_450[32:0];
  assign v_623 = v_622[31:0];
  assign v_624 = {v_625, v_630};
  assign v_625 = {v_626, v_629};
  assign v_626 = v_627[35:32];
  assign v_627 = v_628[38:3];
  assign v_628 = v_451[38:0];
  assign v_629 = v_627[31:0];
  assign v_630 = {v_631, v_633};
  assign v_631 = v_632[2:1];
  assign v_632 = v_628[2:0];
  assign v_633 = v_632[0:0];
  assign v_634 = v_635 & v_419;
  assign v_635 = v_636 & v_411;
  assign v_636 = v_637 | 1'h0;
  assign v_638 = v_639 & v_662;
  assign v_639 = v_640 & v_137;
  assign v_640 = v_641 & v_50;
  assign v_641 = v_642 & v_661;
  assign v_642 = v_643 & v_660;
  assign v_643 = v_644 & v_89;
  assign v_644 = v_645 & v_85;
  assign v_645 = v_646 & v_659;
  assign v_646 = v_647 & v_187;
  assign v_647 = v_648 & v_658;
  assign v_648 = v_649 & v_657;
  assign v_649 = v_650 & v_656;
  assign v_650 = v_651 & v_655;
  assign v_651 = v_652 & v_654;
  assign v_652 = 1'h1 & v_653;
  assign v_653 = ~v_177;
  assign v_654 = ~v_191;
  assign v_655 = ~v_179;
  assign v_656 = ~v_181;
  assign v_657 = ~v_183;
  assign v_658 = ~v_185;
  assign v_659 = ~v_84;
  assign v_660 = ~v_135;
  assign v_661 = ~v_79;
  assign v_662 = ~v_81;
  assign v_663 = v_664 | v_665;
  assign v_664 = mux_664(v_422);
  assign v_665 = mux_665(v_634);
  assign v_666 = mux_666(v_667);
  assign v_667 = v_635 & v_668;
  assign v_668 = ~v_419;
  assign v_669 = v_670 | v_673;
  assign v_670 = mux_670(v_671);
  assign v_671 = v_437 & v_672;
  assign v_672 = ~v_442;
  assign v_673 = mux_673(v_674);
  assign v_674 = ~v_675;
  assign v_675 = v_671 | v_676;
  assign v_676 = v_417 | v_667;
  assign v_677 = {{31{1'b0}}, v_678};
  assign v_678 = v_679 | 1'h0;
  assign v_679 = ~v_680;
  assign v_681 = v_682 | v_686;
  assign v_682 = act_683 & 1'h1;
  assign act_683 = v_684 & v_408;
  assign v_684 = v_685 == 12'h803;
  assign v_685 = v_115[11:0];
  assign v_686 = v_687 & 1'h1;
  assign v_687 = v_688 & v_689;
  assign v_688 = ~act_683;
  assign v_689 = v_690 | v_696;
  assign v_690 = v_691 | v_694;
  assign v_691 = mux_691(v_692);
  assign v_692 = v_693 & 1'h1;
  assign v_693 = out_consume_en;
  assign v_694 = mux_694(v_695);
  assign v_695 = ~v_692;
  assign v_696 = ~v_680;
  assign v_697 = v_698 | v_699;
  assign v_698 = mux_698(v_682);
  assign v_699 = mux_699(v_686);
  assign v_700 = mux_700(v_701);
  assign v_701 = v_702 & v_712;
  assign v_702 = v_703 != 5'h0;
  assign v_703 = {v_704, v_705};
  assign v_704 = v_104[11:11];
  assign v_705 = {v_706, v_707};
  assign v_706 = v_104[10:10];
  assign v_707 = {v_708, v_709};
  assign v_708 = v_104[9:9];
  assign v_709 = {v_710, v_711};
  assign v_710 = v_104[8:8];
  assign v_711 = v_104[7:7];
  assign v_712 = v_713 & v_408;
  assign v_713 = v_114 == 12'h342;
  assign v_715 = v_716 | v_763;
  assign v_716 = v_717 & v_411;
  assign v_717 = v_718 | 1'h0;
  assign v_719 = v_720 & v_761;
  assign v_720 = v_721 & v_137;
  assign v_721 = v_722 & v_50;
  assign v_722 = v_723 & v_760;
  assign v_723 = v_724 & v_759;
  assign v_724 = v_725 & v_89;
  assign v_725 = v_726 & v_85;
  assign v_726 = v_727 & v_84;
  assign v_727 = v_728 & v_758;
  assign v_728 = v_729 & v_757;
  assign v_729 = v_730 & v_756;
  assign v_730 = v_731 & v_754;
  assign v_731 = v_732 & v_752;
  assign v_732 = v_733 & v_750;
  assign v_733 = v_734 & v_748;
  assign v_734 = v_735 & v_747;
  assign v_735 = v_736 & v_746;
  assign v_736 = v_737 & v_745;
  assign v_737 = v_738 & v_744;
  assign v_738 = v_739 & v_743;
  assign v_739 = v_740 & v_742;
  assign v_740 = 1'h1 & v_741;
  assign v_741 = ~v_177;
  assign v_742 = ~v_191;
  assign v_743 = ~v_179;
  assign v_744 = ~v_181;
  assign v_745 = ~v_183;
  assign v_746 = ~v_185;
  assign v_747 = ~v_187;
  assign v_748 = ~v_749;
  assign v_749 = v_51[24:24];
  assign v_750 = ~v_751;
  assign v_751 = v_51[23:23];
  assign v_752 = ~v_753;
  assign v_753 = v_51[22:22];
  assign v_754 = ~v_755;
  assign v_755 = v_51[21:21];
  assign v_756 = ~v_81;
  assign v_757 = ~v_83;
  assign v_758 = ~v_87;
  assign v_759 = ~v_135;
  assign v_760 = ~v_79;
  assign v_761 = ~v_762;
  assign v_762 = v_51[20:20];
  assign v_763 = v_764 | v_766;
  assign v_764 = v_765 & v_408;
  assign v_765 = v_685 == 12'h342;
  assign v_766 = v_767 & v_411;
  assign v_767 = v_768 | 1'h0;
  assign v_769 = v_720 & v_762;
  assign v_770 = v_771 | v_773;
  assign v_771 = mux_771(v_716);
  assign v_772 = {1'h0, 31'h8};
  assign v_773 = v_774 | v_775;
  assign v_774 = mux_774(v_764);
  assign v_775 = mux_775(v_766);
  assign v_776 = {1'h0, 31'h3};
  assign v_777 = v_778 | v_795;
  assign v_778 = mux_778(v_779);
  assign v_779 = v_780 & v_790;
  assign v_780 = v_781 != 5'h0;
  assign v_781 = {v_782, v_783};
  assign v_782 = v_104[11:11];
  assign v_783 = {v_784, v_785};
  assign v_784 = v_104[10:10];
  assign v_785 = {v_786, v_787};
  assign v_786 = v_104[9:9];
  assign v_787 = {v_788, v_789};
  assign v_788 = v_104[8:8];
  assign v_789 = v_104[7:7];
  assign v_790 = v_791 & v_408;
  assign v_791 = v_114 == 12'h341;
  assign v_793 = v_794 & v_408;
  assign v_794 = v_685 == 12'h341;
  assign v_795 = mux_795(v_796);
  assign v_796 = v_797 & v_807;
  assign v_797 = v_798 != 5'h0;
  assign v_798 = {v_799, v_800};
  assign v_799 = v_104[11:11];
  assign v_800 = {v_801, v_802};
  assign v_801 = v_104[10:10];
  assign v_802 = {v_803, v_804};
  assign v_803 = v_104[9:9];
  assign v_804 = {v_805, v_806};
  assign v_805 = v_104[8:8];
  assign v_806 = v_104[7:7];
  assign v_807 = v_808 & v_408;
  assign v_808 = v_114 == 12'h300;
  assign v_810 = v_811 & v_408;
  assign v_811 = v_685 == 12'h300;
  assign v_812 = v_813 | v_865;
  assign v_813 = v_814 | v_833;
  assign v_814 = mux_814(v_815);
  assign v_815 = v_816 & v_826;
  assign v_816 = v_817 != 5'h0;
  assign v_817 = {v_818, v_819};
  assign v_818 = v_104[11:11];
  assign v_819 = {v_820, v_821};
  assign v_820 = v_104[10:10];
  assign v_821 = {v_822, v_823};
  assign v_822 = v_104[9:9];
  assign v_823 = {v_824, v_825};
  assign v_824 = v_104[8:8];
  assign v_825 = v_104[7:7];
  assign v_826 = v_827 & v_411;
  assign v_827 = v_828 | v_829;
  assign v_829 = v_39 | 1'h0;
  assign v_830 = v_831 + 32'h4;
  assign v_833 = mux_833(v_834);
  assign v_834 = v_835 & v_845;
  assign v_835 = v_836 != 5'h0;
  assign v_836 = {v_837, v_838};
  assign v_837 = v_104[11:11];
  assign v_838 = {v_839, v_840};
  assign v_839 = v_104[10:10];
  assign v_840 = {v_841, v_842};
  assign v_841 = v_104[9:9];
  assign v_842 = {v_843, v_844};
  assign v_843 = v_104[8:8];
  assign v_844 = v_104[7:7];
  assign v_845 = v_846 & v_411;
  assign v_846 = v_847 | v_854;
  assign v_848 = v_849 | v_195;
  assign v_849 = v_850 & v_87;
  assign v_850 = v_851 & v_853;
  assign v_851 = v_852 & v_81;
  assign v_852 = v_199 & v_85;
  assign v_853 = ~v_83;
  assign v_854 = v_855 | 1'h0;
  assign v_856 = v_857 | v_159;
  assign v_857 = v_160 & v_85;
  assign v_858 = v_859[31:0];
  assign v_859 = $signed(v_860) >>> v_864;
  assign v_860 = {v_861, v_91};
  assign v_861 = mux_861(v_862);
  assign v_862 = v_855 | 1'h0;
  assign v_863 = v_91[31:31];
  assign v_864 = v_115[4:0];
  assign v_865 = v_866 | v_889;
  assign v_866 = mux_866(v_867);
  assign v_867 = v_868 & v_878;
  assign v_868 = v_869 != 5'h0;
  assign v_869 = {v_870, v_871};
  assign v_870 = v_104[11:11];
  assign v_871 = {v_872, v_873};
  assign v_872 = v_104[10:10];
  assign v_873 = {v_874, v_875};
  assign v_874 = v_104[9:9];
  assign v_875 = {v_876, v_877};
  assign v_876 = v_104[8:8];
  assign v_877 = v_104[7:7];
  assign v_878 = v_879 & v_411;
  assign v_879 = v_880 | 1'h0;
  assign v_881 = v_882 | v_203;
  assign v_882 = v_883 & v_87;
  assign v_883 = v_884 & v_886;
  assign v_884 = v_852 & v_885;
  assign v_885 = ~v_81;
  assign v_886 = ~v_83;
  assign v_887 = v_91 << v_888;
  assign v_888 = v_115[4:0];
  assign v_889 = mux_889(v_890);
  assign v_890 = v_891 & v_901;
  assign v_891 = v_892 != 5'h0;
  assign v_892 = {v_893, v_894};
  assign v_893 = v_104[11:11];
  assign v_894 = {v_895, v_896};
  assign v_895 = v_104[10:10];
  assign v_896 = {v_897, v_898};
  assign v_897 = v_104[9:9];
  assign v_898 = {v_899, v_900};
  assign v_899 = v_104[8:8];
  assign v_900 = v_104[7:7];
  assign v_901 = v_902 & v_411;
  assign v_902 = v_903 | 1'h0;
  assign v_904 = v_831 + v_115;
  assign v_905 = v_906 | v_981;
  assign v_906 = v_907 | v_942;
  assign v_907 = v_908 | v_923;
  assign v_908 = mux_908(v_909);
  assign v_909 = v_910 & v_920;
  assign v_910 = v_911 != 5'h0;
  assign v_911 = {v_912, v_913};
  assign v_912 = v_104[11:11];
  assign v_913 = {v_914, v_915};
  assign v_914 = v_104[10:10];
  assign v_915 = {v_916, v_917};
  assign v_916 = v_104[9:9];
  assign v_917 = {v_918, v_919};
  assign v_918 = v_104[8:8];
  assign v_919 = v_104[7:7];
  assign v_920 = v_921 & v_411;
  assign v_921 = v_922 | 1'h0;
  assign v_923 = mux_923(v_924);
  assign v_924 = v_925 & v_935;
  assign v_925 = v_926 != 5'h0;
  assign v_926 = {v_927, v_928};
  assign v_927 = v_104[11:11];
  assign v_928 = {v_929, v_930};
  assign v_929 = v_104[10:10];
  assign v_930 = {v_931, v_932};
  assign v_931 = v_104[9:9];
  assign v_932 = {v_933, v_934};
  assign v_933 = v_104[8:8];
  assign v_934 = v_104[7:7];
  assign v_935 = v_936 & v_411;
  assign v_936 = v_937 | 1'h0;
  assign v_938 = v_939 | v_208;
  assign v_939 = v_850 & v_940;
  assign v_940 = ~v_87;
  assign v_941 = v_91 ^ v_115;
  assign v_942 = v_943 | v_963;
  assign v_943 = mux_943(v_944);
  assign v_944 = v_945 & v_955;
  assign v_945 = v_946 != 5'h0;
  assign v_946 = {v_947, v_948};
  assign v_947 = v_104[11:11];
  assign v_948 = {v_949, v_950};
  assign v_949 = v_104[10:10];
  assign v_950 = {v_951, v_952};
  assign v_951 = v_104[9:9];
  assign v_952 = {v_953, v_954};
  assign v_953 = v_104[8:8];
  assign v_954 = v_104[7:7];
  assign v_955 = v_956 & v_411;
  assign v_956 = v_957 | 1'h0;
  assign v_958 = v_959 | v_218;
  assign v_959 = v_960 & v_961;
  assign v_960 = v_851 & v_83;
  assign v_961 = ~v_87;
  assign v_962 = v_91 | v_115;
  assign v_963 = mux_963(v_964);
  assign v_964 = v_965 & v_975;
  assign v_965 = v_966 != 5'h0;
  assign v_966 = {v_967, v_968};
  assign v_967 = v_104[11:11];
  assign v_968 = {v_969, v_970};
  assign v_969 = v_104[10:10];
  assign v_970 = {v_971, v_972};
  assign v_971 = v_104[9:9];
  assign v_972 = {v_973, v_974};
  assign v_973 = v_104[8:8];
  assign v_974 = v_104[7:7];
  assign v_975 = v_976 & v_411;
  assign v_976 = v_977 | 1'h0;
  assign v_978 = v_979 | v_227;
  assign v_979 = v_960 & v_87;
  assign v_980 = v_91 & v_115;
  assign v_981 = v_982 | v_1059;
  assign v_982 = v_983 | v_1037;
  assign v_983 = mux_983(v_984);
  assign v_984 = v_985 & v_995;
  assign v_985 = v_986 != 5'h0;
  assign v_986 = {v_987, v_988};
  assign v_987 = v_104[11:11];
  assign v_988 = {v_989, v_990};
  assign v_989 = v_104[10:10];
  assign v_990 = {v_991, v_992};
  assign v_991 = v_104[9:9];
  assign v_992 = {v_993, v_994};
  assign v_993 = v_104[8:8];
  assign v_994 = v_104[7:7];
  assign v_995 = v_996 & v_411;
  assign v_996 = v_997 | v_1002;
  assign v_998 = v_999 | v_242;
  assign v_999 = v_1000 & v_1001;
  assign v_1000 = v_884 & v_83;
  assign v_1001 = ~v_87;
  assign v_1002 = v_1003 | 1'h0;
  assign v_1004 = v_1005 | v_233;
  assign v_1005 = v_1000 & v_87;
  assign v_1006 = {{31{1'b0}}, v_1007};
  assign v_1007 = v_1008[32:32];
  assign v_1008 = v_1009 + v_1036;
  assign v_1009 = v_1010 + v_1026;
  assign v_1010 = {v_1011, v_91};
  assign v_1011 = mux_1011(v_1012);
  assign v_1012 = v_1003 | v_1013;
  assign v_1013 = v_1014 | v_1019;
  assign v_1015 = v_1016 & v_1018;
  assign v_1016 = v_1017 & v_85;
  assign v_1017 = v_221 & v_84;
  assign v_1018 = ~v_89;
  assign v_1019 = v_1020 | 1'h0;
  assign v_1021 = v_1022 & v_1024;
  assign v_1022 = v_1023 & v_85;
  assign v_1023 = v_230 & v_84;
  assign v_1024 = ~v_89;
  assign v_1025 = v_91[31:31];
  assign v_1026 = mux_1026(v_1027);
  assign v_1027 = v_1028 | 1'h0;
  assign v_1029 = v_1030 | v_244;
  assign v_1030 = v_883 & v_1031;
  assign v_1031 = ~v_87;
  assign v_1032 = ~v_1033;
  assign v_1033 = {v_1034, v_115};
  assign v_1034 = mux_1034(v_1012);
  assign v_1035 = v_115[31:31];
  assign v_1036 = mux_1036(v_1027);
  assign v_1037 = mux_1037(v_1038);
  assign v_1038 = v_1039 & v_1049;
  assign v_1039 = v_1040 != 5'h0;
  assign v_1040 = {v_1041, v_1042};
  assign v_1041 = v_104[11:11];
  assign v_1042 = {v_1043, v_1044};
  assign v_1043 = v_104[10:10];
  assign v_1044 = {v_1045, v_1046};
  assign v_1045 = v_104[9:9];
  assign v_1046 = {v_1047, v_1048};
  assign v_1047 = v_104[8:8];
  assign v_1048 = v_104[7:7];
  assign v_1049 = v_1050 & v_411;
  assign v_1050 = v_1028 | v_1051;
  assign v_1051 = v_1052 | 1'h0;
  assign v_1053 = v_1054 & v_85;
  assign v_1054 = v_1055 & v_1057;
  assign v_1055 = v_162 & v_1056;
  assign v_1056 = ~v_81;
  assign v_1057 = ~v_87;
  assign v_1058 = v_1008[31:0];
  assign v_1059 = v_1060 | v_1062;
  assign v_1060 = mux_1060(v_1061);
  assign v_1061 = ~act_96;
  assign v_1062 = v_1063 | v_1066;
  assign v_1063 = mux_1063(v_100);
  assign v_1064 = {{24{1'b0}}, v_1065};
  assign v_1065 = in0_peek;
  assign v_1066 = mux_1066(v_1067);
  assign v_1067 = v_1068 & v_1078;
  assign v_1068 = v_1069 != 5'h0;
  assign v_1069 = {v_1070, v_1071};
  assign v_1070 = v_104[11:11];
  assign v_1071 = {v_1072, v_1073};
  assign v_1072 = v_104[10:10];
  assign v_1073 = {v_1074, v_1075};
  assign v_1074 = v_104[9:9];
  assign v_1075 = {v_1076, v_1077};
  assign v_1076 = v_104[8:8];
  assign v_1077 = v_104[7:7];
  assign v_1078 = v_1079 & v_408;
  assign v_1079 = v_114 == 12'h804;
  assign v_1080 = {{31{1'b0}}, v_1081};
  assign v_1081 = in0_canPeek;
  assign v_1082 = mux_1082(v_308);
  assign v_1083 = v_1084 | v_1359;
  assign v_1084 = mux_1084(act_284);
  assign v_1085 = v_1086[31:0];
  assign v_1086 = mux_1086(v_13);
  assign v_1087 = {v_1088, v_1281};
  assign v_1088 = v_1089[37:32];
  assign v_1089 = mux_1089(v_426);
  assign v_1090 = {v_1091, v_1135};
  assign v_1091 = v_1092[69:64];
  assign v_1092 = v_1093[72:3];
  assign v_1093 = {v_1094, v_1128};
  assign v_1094 = {v_1095, v_1124};
  assign v_1095 = v_1096[69:64];
  assign v_1096 = v_1097[72:3];
  assign v_1098 = {v_1099, v_1117};
  assign v_1099 = {v_1100, v_1113};
  assign v_1100 = v_1101[69:64];
  assign v_1101 = v_1102[72:3];
  assign v_1102 = {v_1103, v_1105};
  assign v_1103 = {6'bxxxxxx, v_1104};
  assign v_1104 = {v_91, v_517};
  assign v_1105 = {v_1106, v_1110};
  assign v_1106 = v_1107 == 2'h0;
  assign v_1107 = {v_1108, v_1109};
  assign v_1110 = {v_1111, v_1112};
  assign v_1111 = v_1107 == 2'h3;
  assign v_1112 = v_1107[1:1];
  assign v_1113 = {v_1114, v_1116};
  assign v_1114 = v_1115[63:32];
  assign v_1115 = v_1101[63:0];
  assign v_1116 = v_1115[31:0];
  assign v_1117 = {v_1118, v_1120};
  assign v_1118 = v_1119[2:2];
  assign v_1119 = v_1102[2:0];
  assign v_1120 = {v_1121, v_1123};
  assign v_1121 = v_1122[1:1];
  assign v_1122 = v_1119[1:0];
  assign v_1123 = v_1122[0:0];
  assign v_1124 = {v_1125, v_1127};
  assign v_1125 = v_1126[63:32];
  assign v_1126 = v_1096[63:0];
  assign v_1127 = v_1126[31:0];
  assign v_1128 = {v_1129, v_1131};
  assign v_1129 = v_1130[2:2];
  assign v_1130 = v_1097[2:0];
  assign v_1131 = {v_1132, v_1134};
  assign v_1132 = v_1133[1:1];
  assign v_1133 = v_1130[1:0];
  assign v_1134 = v_1133[0:0];
  assign v_1135 = mux_1135(v_1136);
  assign v_1136 = v_1137[2:2];
  assign v_1137 = v_1093[2:0];
  assign v_1138 = v_1139[63:32];
  assign v_1140 = v_1141[63:0];
  assign v_1141 = $signed(v_1142)*$signed(v_1145);
  assign v_1142 = {v_1143, v_91};
  assign v_1143 = mux_1143(v_1111);
  assign v_1144 = v_91[31:31];
  assign v_1145 = {v_1146, v_517};
  assign v_1146 = mux_1146(v_1112);
  assign v_1147 = v_517[31:31];
  assign v_1148 = v_1139[31:0];
  assign v_1149 = {v_1150, v_1205};
  assign v_1150 = v_1151[38:33];
  assign v_1151 = v_1152[77:39];
  assign v_1152 = {v_1153, v_1195};
  assign v_1153 = {v_1154, v_1191};
  assign v_1154 = v_1155[38:33];
  assign v_1155 = v_1156[77:39];
  assign v_1157 = act_436 & 1'h1;
  assign v_1158 = {v_1159, v_1181};
  assign v_1159 = {v_1160, v_1177};
  assign v_1160 = v_1161[38:33];
  assign v_1161 = v_1162[77:39];
  assign v_1162 = {v_1163, v_1167};
  assign v_1163 = {v_1164, v_1165};
  assign v_1164 = v_446[38:33];
  assign v_1165 = {v_444, v_1166};
  assign v_1166 = v_445[31:0];
  assign v_1167 = {v_1168, v_1173};
  assign v_1168 = {v_1169, v_1172};
  assign v_1169 = v_1170[35:32];
  assign v_1170 = v_1171[38:3];
  assign v_1171 = v_447[38:0];
  assign v_1172 = v_1170[31:0];
  assign v_1173 = {v_1174, v_1176};
  assign v_1174 = v_1175[2:1];
  assign v_1175 = v_1171[2:0];
  assign v_1176 = v_1175[0:0];
  assign v_1177 = {v_1178, v_1180};
  assign v_1178 = v_1179[32:32];
  assign v_1179 = v_1161[32:0];
  assign v_1180 = v_1179[31:0];
  assign v_1181 = {v_1182, v_1187};
  assign v_1182 = {v_1183, v_1186};
  assign v_1183 = v_1184[35:32];
  assign v_1184 = v_1185[38:3];
  assign v_1185 = v_1162[38:0];
  assign v_1186 = v_1184[31:0];
  assign v_1187 = {v_1188, v_1190};
  assign v_1188 = v_1189[2:1];
  assign v_1189 = v_1185[2:0];
  assign v_1190 = v_1189[0:0];
  assign v_1191 = {v_1192, v_1194};
  assign v_1192 = v_1193[32:32];
  assign v_1193 = v_1155[32:0];
  assign v_1194 = v_1193[31:0];
  assign v_1195 = {v_1196, v_1201};
  assign v_1196 = {v_1197, v_1200};
  assign v_1197 = v_1198[35:32];
  assign v_1198 = v_1199[38:3];
  assign v_1199 = v_1156[38:0];
  assign v_1200 = v_1198[31:0];
  assign v_1201 = {v_1202, v_1204};
  assign v_1202 = v_1203[2:1];
  assign v_1203 = v_1199[2:0];
  assign v_1204 = v_1203[0:0];
  assign v_1205 = v_1206 | v_1264;
  assign v_1206 = mux_1206(v_1207);
  assign v_1207 = v_1208 == 2'h0;
  assign v_1208 = v_1209[2:1];
  assign v_1209 = v_1210[2:0];
  assign v_1210 = v_1152[38:0];
  assign v_1211 = {v_1212, v_1216};
  assign v_1212 = mux_1212(v_1213);
  assign v_1213 = v_1209[0:0];
  assign v_1214 = {{23{v_1215[0]}}, v_1215};
  assign v_1215 = v_1216[7:7];
  assign v_1216 = v_1217 | v_1257;
  assign v_1217 = v_1218 | v_1254;
  assign v_1218 = mux_1218(v_1219);
  assign v_1219 = v_1220 == 2'h0;
  assign v_1220 = v_1221[1:0];
  assign v_1221 = v_1222[31:0];
  assign v_1222 = v_1151[32:0];
  assign v_1223 = v_1224[7:0];
  BlockRAMBE#
    (.INIT_FILE("data.mif"), .ADDR_WIDTH(9), .DATA_WIDTH(32))
    ram1224
      (.CLK(clock),
       .ADDR(v_1225),
       .DI(v_1237),
       .WE(v_1241),
       .RE(v_1245),
       .BE(v_1250),
       .DO(v_1224));
  assign v_1225 = v_1226 | v_1232;
  assign v_1226 = mux_1226(v_1227);
  assign v_1227 = ~v_1228;
  assign v_1228 = v_1229 | v_1231;
  assign v_1229 = v_1157 & v_1230;
  assign v_1230 = ~v_444;
  assign v_1231 = v_1157 & v_444;
  assign v_1232 = v_1233 | v_1236;
  assign v_1233 = mux_1233(v_1229);
  assign v_1234 = v_1235[8:0];
  assign v_1235 = v_1166[31:2];
  assign v_1236 = mux_1236(v_1231);
  assign v_1237 = v_1238 | v_1239;
  assign v_1238 = mux_1238(v_1231);
  assign v_1239 = mux_1239(v_1240);
  assign v_1240 = ~v_1231;
  assign v_1241 = v_1242 | v_1243;
  assign v_1242 = mux_1242(v_1231);
  assign v_1243 = mux_1243(v_1244);
  assign v_1244 = ~v_1231;
  assign v_1245 = v_1246 | v_1248;
  assign v_1246 = mux_1246(v_1247);
  assign v_1247 = v_428 & 1'h1;
  assign v_1248 = mux_1248(v_1249);
  assign v_1249 = ~v_1247;
  assign v_1250 = v_1251 | v_1252;
  assign v_1251 = mux_1251(v_1231);
  assign v_1252 = mux_1252(v_1253);
  assign v_1253 = ~v_1231;
  assign v_1254 = mux_1254(v_1255);
  assign v_1255 = v_1220 == 2'h1;
  assign v_1256 = v_1224[15:8];
  assign v_1257 = v_1258 | v_1261;
  assign v_1258 = mux_1258(v_1259);
  assign v_1259 = v_1220 == 2'h2;
  assign v_1260 = v_1224[23:16];
  assign v_1261 = mux_1261(v_1262);
  assign v_1262 = v_1220 == 2'h3;
  assign v_1263 = v_1224[31:24];
  assign v_1264 = v_1265 | v_1270;
  assign v_1265 = mux_1265(v_1266);
  assign v_1266 = v_1208 == 2'h2;
  assign v_1267 = {v_1263, v_1268};
  assign v_1268 = {v_1260, v_1269};
  assign v_1269 = {v_1256, v_1223};
  assign v_1270 = mux_1270(v_1271);
  assign v_1271 = v_1208 == 2'h1;
  assign v_1272 = {v_1273, v_1276};
  assign v_1273 = mux_1273(v_1213);
  assign v_1274 = {{15{v_1275[0]}}, v_1275};
  assign v_1275 = v_1276[15:15];
  assign v_1276 = mux_1276(v_1277);
  assign v_1277 = v_1278 == 1'h0;
  assign v_1278 = v_1220[1:1];
  assign v_1279 = {v_1263, v_1260};
  assign v_1280 = {v_1256, v_1223};
  assign v_1281 = v_1089[31:0];
  assign v_1282 = {v_1283, v_1284};
  assign v_1285 = mux_1285(v_1286);
  assign v_1287 = v_22 & 1'h1;
  assign v_1288 = v_1289 & v_1310;
  assign v_1289 = v_1290 & v_1296;
  assign v_1291 = v_1292[0:0];
  assign v_1292 = ~v_1293;
  assign v_1293 = {v_1294, v_1295};
  assign v_1296 = ~v_1297;
  assign v_1297 = v_1298 == 32'h0;
  assign v_1299 = v_25 | v_1300;
  assign v_1300 = v_1301 & v_1302;
  assign v_1301 = v_1298[31:31];
  assign v_1302 = v_1303 & v_1287;
  assign v_1303 = v_1290 & v_1304;
  assign v_1304 = ~v_1297;
  assign v_1305 = v_1306 | v_1307;
  assign v_1306 = mux_1306(v_25);
  assign v_1307 = mux_1307(v_1300);
  assign v_1308 = v_1309 + 32'h1;
  assign v_1309 = ~v_1298;
  assign v_1310 = mux_1310(v_1311);
  assign v_1312 = v_1293[1:1];
  assign v_1313 = v_1314 ^ v_1301;
  assign v_1314 = v_1315[31:31];
  assign v_1316 = v_1317 | v_1318;
  assign v_1317 = v_1314 & v_1302;
  assign v_1318 = v_25 | v_1319;
  assign v_1319 = v_1320 & 1'h1;
  assign v_1320 = v_18 & v_1321;
  assign v_1321 = v_1322 != 6'h0;
  assign v_1323 = v_1319 | v_1287;
  assign v_1324 = v_1325 | v_1327;
  assign v_1325 = mux_1325(v_1319);
  assign v_1326 = v_1322 - 6'h1;
  assign v_1327 = mux_1327(v_1287);
  assign v_1328 = v_1329 | v_1332;
  assign v_1329 = mux_1329(v_1317);
  assign v_1330 = v_1331 + 32'h1;
  assign v_1331 = ~v_1315;
  assign v_1332 = v_1333 | v_1334;
  assign v_1333 = mux_1333(v_25);
  assign v_1334 = mux_1334(v_1319);
  assign v_1335 = v_1315 << 1'h1;
  assign v_1336 = mux_1336(v_1311);
  assign v_1338 = v_1319 | v_1287;
  assign v_1339 = v_1340 | v_1356;
  assign v_1340 = mux_1340(v_1319);
  assign v_1341 = v_1342 | v_1343;
  assign v_1342 = v_1337 << 1'h1;
  assign v_1343 = mux_1343(v_1344);
  assign v_1344 = v_1298 <= v_1345;
  assign v_1345 = v_1346 | v_1354;
  assign v_1346 = v_1347 << 1'h1;
  assign v_1348 = v_1319 | v_1287;
  assign v_1349 = v_1350 | v_1353;
  assign v_1350 = mux_1350(v_1319);
  assign v_1351 = v_1345 - v_1352;
  assign v_1352 = mux_1352(v_1344);
  assign v_1353 = mux_1353(v_1287);
  assign v_1354 = {{31{1'b0}}, v_1355};
  assign v_1355 = v_1315[31:31];
  assign v_1356 = mux_1356(v_1287);
  assign v_1357 = v_1358 + 32'h1;
  assign v_1358 = ~v_1336;
  assign v_1359 = mux_1359(v_1360);
  assign v_1360 = ~act_284;
  assign v_1361 = mux_1361(v_1362);
  assign v_1362 = ~act_333;
  assign v_1363 = v_1364 | v_1365;
  assign v_1364 = mux_1364(act_333);
  assign v_1365 = mux_1365(v_1366);
  assign v_1366 = ~act_333;
  assign v_1367 = mux_1367(v_1368);
  assign v_1368 = ~1'h0;
  assign v_1370 = v_1371 | v_1372;
  assign v_1371 = mux_1371(act_333);
  assign v_1372 = mux_1372(v_1373);
  assign v_1373 = ~act_333;
  assign v_1374 = {v_1375, v_1406};
  assign v_1375 = v_1376 | v_1391;
  assign v_1376 = v_1377 | v_1384;
  assign v_1377 = v_1378 | v_1381;
  assign v_1378 = v_1379 | v_1380;
  assign v_1379 = v_121 & v_177;
  assign v_1380 = v_123 & v_177;
  assign v_1381 = v_1382 | v_1383;
  assign v_1382 = v_139 & v_177;
  assign v_1383 = v_40 & v_177;
  assign v_1384 = v_1385 | v_1388;
  assign v_1385 = v_1386 | v_1387;
  assign v_1386 = v_153 & v_177;
  assign v_1387 = v_159 & v_749;
  assign v_1388 = v_1389 | v_1390;
  assign v_1389 = v_195 & v_749;
  assign v_1390 = v_203 & v_749;
  assign v_1391 = v_1392 | v_1399;
  assign v_1392 = v_1393 | v_1396;
  assign v_1393 = v_1394 | v_1395;
  assign v_1394 = v_208 & v_177;
  assign v_1395 = v_218 & v_177;
  assign v_1396 = v_1397 | v_1398;
  assign v_1397 = v_227 & v_177;
  assign v_1398 = v_233 & v_177;
  assign v_1399 = v_1400 | v_1403;
  assign v_1400 = v_1401 | v_1402;
  assign v_1401 = v_242 & v_177;
  assign v_1402 = v_244 & v_177;
  assign v_1403 = v_1404 | v_1405;
  assign v_1404 = v_252 & v_177;
  assign v_1405 = v_254 & v_177;
  assign v_1406 = {v_1407, v_1438};
  assign v_1407 = v_1408 | v_1423;
  assign v_1408 = v_1409 | v_1416;
  assign v_1409 = v_1410 | v_1413;
  assign v_1410 = v_1411 | v_1412;
  assign v_1411 = v_121 & v_177;
  assign v_1412 = v_123 & v_177;
  assign v_1413 = v_1414 | v_1415;
  assign v_1414 = v_139 & v_177;
  assign v_1415 = v_40 & v_177;
  assign v_1416 = v_1417 | v_1420;
  assign v_1417 = v_1418 | v_1419;
  assign v_1418 = v_153 & v_177;
  assign v_1419 = v_159 & v_749;
  assign v_1420 = v_1421 | v_1422;
  assign v_1421 = v_195 & v_749;
  assign v_1422 = v_203 & v_749;
  assign v_1423 = v_1424 | v_1431;
  assign v_1424 = v_1425 | v_1428;
  assign v_1425 = v_1426 | v_1427;
  assign v_1426 = v_208 & v_177;
  assign v_1427 = v_218 & v_177;
  assign v_1428 = v_1429 | v_1430;
  assign v_1429 = v_227 & v_177;
  assign v_1430 = v_233 & v_177;
  assign v_1431 = v_1432 | v_1435;
  assign v_1432 = v_1433 | v_1434;
  assign v_1433 = v_242 & v_177;
  assign v_1434 = v_244 & v_177;
  assign v_1435 = v_1436 | v_1437;
  assign v_1436 = v_252 & v_191;
  assign v_1437 = v_254 & v_191;
  assign v_1438 = {v_1439, v_1470};
  assign v_1439 = v_1440 | v_1455;
  assign v_1440 = v_1441 | v_1448;
  assign v_1441 = v_1442 | v_1445;
  assign v_1442 = v_1443 | v_1444;
  assign v_1443 = v_121 & v_177;
  assign v_1444 = v_123 & v_177;
  assign v_1445 = v_1446 | v_1447;
  assign v_1446 = v_139 & v_177;
  assign v_1447 = v_40 & v_177;
  assign v_1448 = v_1449 | v_1452;
  assign v_1449 = v_1450 | v_1451;
  assign v_1450 = v_153 & v_177;
  assign v_1451 = v_159 & v_749;
  assign v_1452 = v_1453 | v_1454;
  assign v_1453 = v_195 & v_749;
  assign v_1454 = v_203 & v_749;
  assign v_1455 = v_1456 | v_1463;
  assign v_1456 = v_1457 | v_1460;
  assign v_1457 = v_1458 | v_1459;
  assign v_1458 = v_208 & v_177;
  assign v_1459 = v_218 & v_177;
  assign v_1460 = v_1461 | v_1462;
  assign v_1461 = v_227 & v_177;
  assign v_1462 = v_233 & v_177;
  assign v_1463 = v_1464 | v_1467;
  assign v_1464 = v_1465 | v_1466;
  assign v_1465 = v_242 & v_177;
  assign v_1466 = v_244 & v_177;
  assign v_1467 = v_1468 | v_1469;
  assign v_1468 = v_252 & v_179;
  assign v_1469 = v_254 & v_179;
  assign v_1470 = {v_1471, v_1502};
  assign v_1471 = v_1472 | v_1487;
  assign v_1472 = v_1473 | v_1480;
  assign v_1473 = v_1474 | v_1477;
  assign v_1474 = v_1475 | v_1476;
  assign v_1475 = v_121 & v_177;
  assign v_1476 = v_123 & v_177;
  assign v_1477 = v_1478 | v_1479;
  assign v_1478 = v_139 & v_177;
  assign v_1479 = v_40 & v_177;
  assign v_1480 = v_1481 | v_1484;
  assign v_1481 = v_1482 | v_1483;
  assign v_1482 = v_153 & v_177;
  assign v_1483 = v_159 & v_749;
  assign v_1484 = v_1485 | v_1486;
  assign v_1485 = v_195 & v_749;
  assign v_1486 = v_203 & v_749;
  assign v_1487 = v_1488 | v_1495;
  assign v_1488 = v_1489 | v_1492;
  assign v_1489 = v_1490 | v_1491;
  assign v_1490 = v_208 & v_177;
  assign v_1491 = v_218 & v_177;
  assign v_1492 = v_1493 | v_1494;
  assign v_1493 = v_227 & v_177;
  assign v_1494 = v_233 & v_177;
  assign v_1495 = v_1496 | v_1499;
  assign v_1496 = v_1497 | v_1498;
  assign v_1497 = v_242 & v_177;
  assign v_1498 = v_244 & v_177;
  assign v_1499 = v_1500 | v_1501;
  assign v_1500 = v_252 & v_181;
  assign v_1501 = v_254 & v_181;
  assign v_1502 = {v_1503, v_1534};
  assign v_1503 = v_1504 | v_1519;
  assign v_1504 = v_1505 | v_1512;
  assign v_1505 = v_1506 | v_1509;
  assign v_1506 = v_1507 | v_1508;
  assign v_1507 = v_121 & v_177;
  assign v_1508 = v_123 & v_177;
  assign v_1509 = v_1510 | v_1511;
  assign v_1510 = v_139 & v_177;
  assign v_1511 = v_40 & v_177;
  assign v_1512 = v_1513 | v_1516;
  assign v_1513 = v_1514 | v_1515;
  assign v_1514 = v_153 & v_177;
  assign v_1515 = v_159 & v_749;
  assign v_1516 = v_1517 | v_1518;
  assign v_1517 = v_195 & v_749;
  assign v_1518 = v_203 & v_749;
  assign v_1519 = v_1520 | v_1527;
  assign v_1520 = v_1521 | v_1524;
  assign v_1521 = v_1522 | v_1523;
  assign v_1522 = v_208 & v_177;
  assign v_1523 = v_218 & v_177;
  assign v_1524 = v_1525 | v_1526;
  assign v_1525 = v_227 & v_177;
  assign v_1526 = v_233 & v_177;
  assign v_1527 = v_1528 | v_1531;
  assign v_1528 = v_1529 | v_1530;
  assign v_1529 = v_242 & v_177;
  assign v_1530 = v_244 & v_177;
  assign v_1531 = v_1532 | v_1533;
  assign v_1532 = v_252 & v_183;
  assign v_1533 = v_254 & v_183;
  assign v_1534 = {v_1535, v_1566};
  assign v_1535 = v_1536 | v_1551;
  assign v_1536 = v_1537 | v_1544;
  assign v_1537 = v_1538 | v_1541;
  assign v_1538 = v_1539 | v_1540;
  assign v_1539 = v_121 & v_177;
  assign v_1540 = v_123 & v_177;
  assign v_1541 = v_1542 | v_1543;
  assign v_1542 = v_139 & v_177;
  assign v_1543 = v_40 & v_177;
  assign v_1544 = v_1545 | v_1548;
  assign v_1545 = v_1546 | v_1547;
  assign v_1546 = v_153 & v_177;
  assign v_1547 = v_159 & v_749;
  assign v_1548 = v_1549 | v_1550;
  assign v_1549 = v_195 & v_749;
  assign v_1550 = v_203 & v_749;
  assign v_1551 = v_1552 | v_1559;
  assign v_1552 = v_1553 | v_1556;
  assign v_1553 = v_1554 | v_1555;
  assign v_1554 = v_208 & v_177;
  assign v_1555 = v_218 & v_177;
  assign v_1556 = v_1557 | v_1558;
  assign v_1557 = v_227 & v_177;
  assign v_1558 = v_233 & v_177;
  assign v_1559 = v_1560 | v_1563;
  assign v_1560 = v_1561 | v_1562;
  assign v_1561 = v_242 & v_177;
  assign v_1562 = v_244 & v_177;
  assign v_1563 = v_1564 | v_1565;
  assign v_1564 = v_252 & v_185;
  assign v_1565 = v_254 & v_185;
  assign v_1566 = {v_1567, v_1598};
  assign v_1567 = v_1568 | v_1583;
  assign v_1568 = v_1569 | v_1576;
  assign v_1569 = v_1570 | v_1573;
  assign v_1570 = v_1571 | v_1572;
  assign v_1571 = v_121 & v_177;
  assign v_1572 = v_123 & v_177;
  assign v_1573 = v_1574 | v_1575;
  assign v_1574 = v_139 & v_177;
  assign v_1575 = v_40 & v_177;
  assign v_1576 = v_1577 | v_1580;
  assign v_1577 = v_1578 | v_1579;
  assign v_1578 = v_153 & v_177;
  assign v_1579 = v_159 & v_749;
  assign v_1580 = v_1581 | v_1582;
  assign v_1581 = v_195 & v_749;
  assign v_1582 = v_203 & v_749;
  assign v_1583 = v_1584 | v_1591;
  assign v_1584 = v_1585 | v_1588;
  assign v_1585 = v_1586 | v_1587;
  assign v_1586 = v_208 & v_177;
  assign v_1587 = v_218 & v_177;
  assign v_1588 = v_1589 | v_1590;
  assign v_1589 = v_227 & v_177;
  assign v_1590 = v_233 & v_177;
  assign v_1591 = v_1592 | v_1595;
  assign v_1592 = v_1593 | v_1594;
  assign v_1593 = v_242 & v_177;
  assign v_1594 = v_244 & v_177;
  assign v_1595 = v_1596 | v_1597;
  assign v_1596 = v_252 & v_187;
  assign v_1597 = v_254 & v_187;
  assign v_1598 = {v_1599, v_1630};
  assign v_1599 = v_1600 | v_1615;
  assign v_1600 = v_1601 | v_1608;
  assign v_1601 = v_1602 | v_1605;
  assign v_1602 = v_1603 | v_1604;
  assign v_1603 = v_121 & v_177;
  assign v_1604 = v_123 & v_177;
  assign v_1605 = v_1606 | v_1607;
  assign v_1606 = v_139 & v_177;
  assign v_1607 = v_40 & v_177;
  assign v_1608 = v_1609 | v_1612;
  assign v_1609 = v_1610 | v_1611;
  assign v_1610 = v_153 & v_177;
  assign v_1611 = v_159 & v_749;
  assign v_1612 = v_1613 | v_1614;
  assign v_1613 = v_195 & v_749;
  assign v_1614 = v_203 & v_749;
  assign v_1615 = v_1616 | v_1623;
  assign v_1616 = v_1617 | v_1620;
  assign v_1617 = v_1618 | v_1619;
  assign v_1618 = v_208 & v_177;
  assign v_1619 = v_218 & v_177;
  assign v_1620 = v_1621 | v_1622;
  assign v_1621 = v_227 & v_177;
  assign v_1622 = v_233 & v_177;
  assign v_1623 = v_1624 | v_1627;
  assign v_1624 = v_1625 | v_1626;
  assign v_1625 = v_242 & v_177;
  assign v_1626 = v_244 & v_177;
  assign v_1627 = v_1628 | v_1629;
  assign v_1628 = v_252 & v_749;
  assign v_1629 = v_254 & v_749;
  assign v_1630 = {v_1631, v_1662};
  assign v_1631 = v_1632 | v_1647;
  assign v_1632 = v_1633 | v_1640;
  assign v_1633 = v_1634 | v_1637;
  assign v_1634 = v_1635 | v_1636;
  assign v_1635 = v_121 & v_177;
  assign v_1636 = v_123 & v_177;
  assign v_1637 = v_1638 | v_1639;
  assign v_1638 = v_139 & v_177;
  assign v_1639 = v_40 & v_177;
  assign v_1640 = v_1641 | v_1644;
  assign v_1641 = v_1642 | v_1643;
  assign v_1642 = v_153 & v_177;
  assign v_1643 = v_159 & v_749;
  assign v_1644 = v_1645 | v_1646;
  assign v_1645 = v_195 & v_749;
  assign v_1646 = v_203 & v_749;
  assign v_1647 = v_1648 | v_1655;
  assign v_1648 = v_1649 | v_1652;
  assign v_1649 = v_1650 | v_1651;
  assign v_1650 = v_208 & v_177;
  assign v_1651 = v_218 & v_177;
  assign v_1652 = v_1653 | v_1654;
  assign v_1653 = v_227 & v_177;
  assign v_1654 = v_233 & v_177;
  assign v_1655 = v_1656 | v_1659;
  assign v_1656 = v_1657 | v_1658;
  assign v_1657 = v_242 & v_177;
  assign v_1658 = v_244 & v_177;
  assign v_1659 = v_1660 | v_1661;
  assign v_1660 = v_252 & v_751;
  assign v_1661 = v_254 & v_751;
  assign v_1662 = {v_1663, v_1694};
  assign v_1663 = v_1664 | v_1679;
  assign v_1664 = v_1665 | v_1672;
  assign v_1665 = v_1666 | v_1669;
  assign v_1666 = v_1667 | v_1668;
  assign v_1667 = v_121 & v_177;
  assign v_1668 = v_123 & v_177;
  assign v_1669 = v_1670 | v_1671;
  assign v_1670 = v_139 & v_177;
  assign v_1671 = v_40 & v_177;
  assign v_1672 = v_1673 | v_1676;
  assign v_1673 = v_1674 | v_1675;
  assign v_1674 = v_153 & v_177;
  assign v_1675 = v_159 & v_749;
  assign v_1676 = v_1677 | v_1678;
  assign v_1677 = v_195 & v_749;
  assign v_1678 = v_203 & v_749;
  assign v_1679 = v_1680 | v_1687;
  assign v_1680 = v_1681 | v_1684;
  assign v_1681 = v_1682 | v_1683;
  assign v_1682 = v_208 & v_177;
  assign v_1683 = v_218 & v_177;
  assign v_1684 = v_1685 | v_1686;
  assign v_1685 = v_227 & v_177;
  assign v_1686 = v_233 & v_177;
  assign v_1687 = v_1688 | v_1691;
  assign v_1688 = v_1689 | v_1690;
  assign v_1689 = v_242 & v_177;
  assign v_1690 = v_244 & v_177;
  assign v_1691 = v_1692 | v_1693;
  assign v_1692 = v_252 & v_753;
  assign v_1693 = v_254 & v_753;
  assign v_1694 = {v_1695, v_1726};
  assign v_1695 = v_1696 | v_1711;
  assign v_1696 = v_1697 | v_1704;
  assign v_1697 = v_1698 | v_1701;
  assign v_1698 = v_1699 | v_1700;
  assign v_1699 = v_121 & v_177;
  assign v_1700 = v_123 & v_177;
  assign v_1701 = v_1702 | v_1703;
  assign v_1702 = v_139 & v_177;
  assign v_1703 = v_40 & v_177;
  assign v_1704 = v_1705 | v_1708;
  assign v_1705 = v_1706 | v_1707;
  assign v_1706 = v_153 & v_177;
  assign v_1707 = v_159 & v_749;
  assign v_1708 = v_1709 | v_1710;
  assign v_1709 = v_195 & v_749;
  assign v_1710 = v_203 & v_749;
  assign v_1711 = v_1712 | v_1719;
  assign v_1712 = v_1713 | v_1716;
  assign v_1713 = v_1714 | v_1715;
  assign v_1714 = v_208 & v_177;
  assign v_1715 = v_218 & v_177;
  assign v_1716 = v_1717 | v_1718;
  assign v_1717 = v_227 & v_177;
  assign v_1718 = v_233 & v_177;
  assign v_1719 = v_1720 | v_1723;
  assign v_1720 = v_1721 | v_1722;
  assign v_1721 = v_242 & v_177;
  assign v_1722 = v_244 & v_177;
  assign v_1723 = v_1724 | v_1725;
  assign v_1724 = v_252 & v_755;
  assign v_1725 = v_254 & v_755;
  assign v_1726 = {v_1727, v_1758};
  assign v_1727 = v_1728 | v_1743;
  assign v_1728 = v_1729 | v_1736;
  assign v_1729 = v_1730 | v_1733;
  assign v_1730 = v_1731 | v_1732;
  assign v_1731 = v_121 & v_177;
  assign v_1732 = v_123 & v_177;
  assign v_1733 = v_1734 | v_1735;
  assign v_1734 = v_139 & v_177;
  assign v_1735 = v_40 & v_177;
  assign v_1736 = v_1737 | v_1740;
  assign v_1737 = v_1738 | v_1739;
  assign v_1738 = v_153 & v_177;
  assign v_1739 = v_159 & v_749;
  assign v_1740 = v_1741 | v_1742;
  assign v_1741 = v_195 & v_749;
  assign v_1742 = v_203 & v_749;
  assign v_1743 = v_1744 | v_1751;
  assign v_1744 = v_1745 | v_1748;
  assign v_1745 = v_1746 | v_1747;
  assign v_1746 = v_208 & v_177;
  assign v_1747 = v_218 & v_177;
  assign v_1748 = v_1749 | v_1750;
  assign v_1749 = v_227 & v_177;
  assign v_1750 = v_233 & v_177;
  assign v_1751 = v_1752 | v_1755;
  assign v_1752 = v_1753 | v_1754;
  assign v_1753 = v_242 & v_177;
  assign v_1754 = v_244 & v_177;
  assign v_1755 = v_1756 | v_1757;
  assign v_1756 = v_252 & v_762;
  assign v_1757 = v_254 & v_762;
  assign v_1758 = {v_1759, v_1791};
  assign v_1759 = v_1760 | v_1776;
  assign v_1760 = v_1761 | v_1768;
  assign v_1761 = v_1762 | v_1765;
  assign v_1762 = v_1763 | v_1764;
  assign v_1763 = v_121 & v_177;
  assign v_1764 = v_123 & v_177;
  assign v_1765 = v_1766 | v_1767;
  assign v_1766 = v_139 & v_177;
  assign v_1767 = v_40 & v_177;
  assign v_1768 = v_1769 | v_1773;
  assign v_1769 = v_1770 | v_1772;
  assign v_1770 = v_153 & v_1771;
  assign v_1771 = v_51[19:19];
  assign v_1772 = v_159 & v_749;
  assign v_1773 = v_1774 | v_1775;
  assign v_1774 = v_195 & v_749;
  assign v_1775 = v_203 & v_749;
  assign v_1776 = v_1777 | v_1784;
  assign v_1777 = v_1778 | v_1781;
  assign v_1778 = v_1779 | v_1780;
  assign v_1779 = v_208 & v_177;
  assign v_1780 = v_218 & v_177;
  assign v_1781 = v_1782 | v_1783;
  assign v_1782 = v_227 & v_177;
  assign v_1783 = v_233 & v_177;
  assign v_1784 = v_1785 | v_1788;
  assign v_1785 = v_1786 | v_1787;
  assign v_1786 = v_242 & v_177;
  assign v_1787 = v_244 & v_177;
  assign v_1788 = v_1789 | v_1790;
  assign v_1789 = v_252 & v_1771;
  assign v_1790 = v_254 & v_1771;
  assign v_1791 = {v_1792, v_1824};
  assign v_1792 = v_1793 | v_1809;
  assign v_1793 = v_1794 | v_1801;
  assign v_1794 = v_1795 | v_1798;
  assign v_1795 = v_1796 | v_1797;
  assign v_1796 = v_121 & v_177;
  assign v_1797 = v_123 & v_177;
  assign v_1798 = v_1799 | v_1800;
  assign v_1799 = v_139 & v_177;
  assign v_1800 = v_40 & v_177;
  assign v_1801 = v_1802 | v_1806;
  assign v_1802 = v_1803 | v_1805;
  assign v_1803 = v_153 & v_1804;
  assign v_1804 = v_51[18:18];
  assign v_1805 = v_159 & v_749;
  assign v_1806 = v_1807 | v_1808;
  assign v_1807 = v_195 & v_749;
  assign v_1808 = v_203 & v_749;
  assign v_1809 = v_1810 | v_1817;
  assign v_1810 = v_1811 | v_1814;
  assign v_1811 = v_1812 | v_1813;
  assign v_1812 = v_208 & v_177;
  assign v_1813 = v_218 & v_177;
  assign v_1814 = v_1815 | v_1816;
  assign v_1815 = v_227 & v_177;
  assign v_1816 = v_233 & v_177;
  assign v_1817 = v_1818 | v_1821;
  assign v_1818 = v_1819 | v_1820;
  assign v_1819 = v_242 & v_177;
  assign v_1820 = v_244 & v_177;
  assign v_1821 = v_1822 | v_1823;
  assign v_1822 = v_252 & v_1804;
  assign v_1823 = v_254 & v_1804;
  assign v_1824 = {v_1825, v_1857};
  assign v_1825 = v_1826 | v_1842;
  assign v_1826 = v_1827 | v_1834;
  assign v_1827 = v_1828 | v_1831;
  assign v_1828 = v_1829 | v_1830;
  assign v_1829 = v_121 & v_177;
  assign v_1830 = v_123 & v_177;
  assign v_1831 = v_1832 | v_1833;
  assign v_1832 = v_139 & v_177;
  assign v_1833 = v_40 & v_177;
  assign v_1834 = v_1835 | v_1839;
  assign v_1835 = v_1836 | v_1838;
  assign v_1836 = v_153 & v_1837;
  assign v_1837 = v_51[17:17];
  assign v_1838 = v_159 & v_749;
  assign v_1839 = v_1840 | v_1841;
  assign v_1840 = v_195 & v_749;
  assign v_1841 = v_203 & v_749;
  assign v_1842 = v_1843 | v_1850;
  assign v_1843 = v_1844 | v_1847;
  assign v_1844 = v_1845 | v_1846;
  assign v_1845 = v_208 & v_177;
  assign v_1846 = v_218 & v_177;
  assign v_1847 = v_1848 | v_1849;
  assign v_1848 = v_227 & v_177;
  assign v_1849 = v_233 & v_177;
  assign v_1850 = v_1851 | v_1854;
  assign v_1851 = v_1852 | v_1853;
  assign v_1852 = v_242 & v_177;
  assign v_1853 = v_244 & v_177;
  assign v_1854 = v_1855 | v_1856;
  assign v_1855 = v_252 & v_1837;
  assign v_1856 = v_254 & v_1837;
  assign v_1857 = {v_1858, v_1890};
  assign v_1858 = v_1859 | v_1875;
  assign v_1859 = v_1860 | v_1867;
  assign v_1860 = v_1861 | v_1864;
  assign v_1861 = v_1862 | v_1863;
  assign v_1862 = v_121 & v_177;
  assign v_1863 = v_123 & v_177;
  assign v_1864 = v_1865 | v_1866;
  assign v_1865 = v_139 & v_177;
  assign v_1866 = v_40 & v_177;
  assign v_1867 = v_1868 | v_1872;
  assign v_1868 = v_1869 | v_1871;
  assign v_1869 = v_153 & v_1870;
  assign v_1870 = v_51[16:16];
  assign v_1871 = v_159 & v_749;
  assign v_1872 = v_1873 | v_1874;
  assign v_1873 = v_195 & v_749;
  assign v_1874 = v_203 & v_749;
  assign v_1875 = v_1876 | v_1883;
  assign v_1876 = v_1877 | v_1880;
  assign v_1877 = v_1878 | v_1879;
  assign v_1878 = v_208 & v_177;
  assign v_1879 = v_218 & v_177;
  assign v_1880 = v_1881 | v_1882;
  assign v_1881 = v_227 & v_177;
  assign v_1882 = v_233 & v_177;
  assign v_1883 = v_1884 | v_1887;
  assign v_1884 = v_1885 | v_1886;
  assign v_1885 = v_242 & v_177;
  assign v_1886 = v_244 & v_177;
  assign v_1887 = v_1888 | v_1889;
  assign v_1888 = v_252 & v_1870;
  assign v_1889 = v_254 & v_1870;
  assign v_1890 = {v_1891, v_1923};
  assign v_1891 = v_1892 | v_1908;
  assign v_1892 = v_1893 | v_1900;
  assign v_1893 = v_1894 | v_1897;
  assign v_1894 = v_1895 | v_1896;
  assign v_1895 = v_121 & v_177;
  assign v_1896 = v_123 & v_177;
  assign v_1897 = v_1898 | v_1899;
  assign v_1898 = v_139 & v_177;
  assign v_1899 = v_40 & v_177;
  assign v_1900 = v_1901 | v_1905;
  assign v_1901 = v_1902 | v_1904;
  assign v_1902 = v_153 & v_1903;
  assign v_1903 = v_51[15:15];
  assign v_1904 = v_159 & v_749;
  assign v_1905 = v_1906 | v_1907;
  assign v_1906 = v_195 & v_749;
  assign v_1907 = v_203 & v_749;
  assign v_1908 = v_1909 | v_1916;
  assign v_1909 = v_1910 | v_1913;
  assign v_1910 = v_1911 | v_1912;
  assign v_1911 = v_208 & v_177;
  assign v_1912 = v_218 & v_177;
  assign v_1913 = v_1914 | v_1915;
  assign v_1914 = v_227 & v_177;
  assign v_1915 = v_233 & v_177;
  assign v_1916 = v_1917 | v_1920;
  assign v_1917 = v_1918 | v_1919;
  assign v_1918 = v_242 & v_177;
  assign v_1919 = v_244 & v_177;
  assign v_1920 = v_1921 | v_1922;
  assign v_1921 = v_252 & v_1903;
  assign v_1922 = v_254 & v_1903;
  assign v_1923 = {v_1924, v_1955};
  assign v_1924 = v_1925 | v_1940;
  assign v_1925 = v_1926 | v_1933;
  assign v_1926 = v_1927 | v_1930;
  assign v_1927 = v_1928 | v_1929;
  assign v_1928 = v_121 & v_177;
  assign v_1929 = v_123 & v_177;
  assign v_1930 = v_1931 | v_1932;
  assign v_1931 = v_139 & v_177;
  assign v_1932 = v_40 & v_177;
  assign v_1933 = v_1934 | v_1937;
  assign v_1934 = v_1935 | v_1936;
  assign v_1935 = v_153 & v_81;
  assign v_1936 = v_159 & v_749;
  assign v_1937 = v_1938 | v_1939;
  assign v_1938 = v_195 & v_749;
  assign v_1939 = v_203 & v_749;
  assign v_1940 = v_1941 | v_1948;
  assign v_1941 = v_1942 | v_1945;
  assign v_1942 = v_1943 | v_1944;
  assign v_1943 = v_208 & v_177;
  assign v_1944 = v_218 & v_177;
  assign v_1945 = v_1946 | v_1947;
  assign v_1946 = v_227 & v_177;
  assign v_1947 = v_233 & v_177;
  assign v_1948 = v_1949 | v_1952;
  assign v_1949 = v_1950 | v_1951;
  assign v_1950 = v_242 & v_177;
  assign v_1951 = v_244 & v_177;
  assign v_1952 = v_1953 | v_1954;
  assign v_1953 = v_252 & v_81;
  assign v_1954 = v_254 & v_81;
  assign v_1955 = {v_1956, v_1987};
  assign v_1956 = v_1957 | v_1972;
  assign v_1957 = v_1958 | v_1965;
  assign v_1958 = v_1959 | v_1962;
  assign v_1959 = v_1960 | v_1961;
  assign v_1960 = v_121 & v_177;
  assign v_1961 = v_123 & v_177;
  assign v_1962 = v_1963 | v_1964;
  assign v_1963 = v_139 & v_177;
  assign v_1964 = v_40 & v_177;
  assign v_1965 = v_1966 | v_1969;
  assign v_1966 = v_1967 | v_1968;
  assign v_1967 = v_153 & v_83;
  assign v_1968 = v_159 & v_749;
  assign v_1969 = v_1970 | v_1971;
  assign v_1970 = v_195 & v_749;
  assign v_1971 = v_203 & v_749;
  assign v_1972 = v_1973 | v_1980;
  assign v_1973 = v_1974 | v_1977;
  assign v_1974 = v_1975 | v_1976;
  assign v_1975 = v_208 & v_177;
  assign v_1976 = v_218 & v_177;
  assign v_1977 = v_1978 | v_1979;
  assign v_1978 = v_227 & v_177;
  assign v_1979 = v_233 & v_177;
  assign v_1980 = v_1981 | v_1984;
  assign v_1981 = v_1982 | v_1983;
  assign v_1982 = v_242 & v_177;
  assign v_1983 = v_244 & v_177;
  assign v_1984 = v_1985 | v_1986;
  assign v_1985 = v_252 & v_83;
  assign v_1986 = v_254 & v_83;
  assign v_1987 = {v_1988, v_2019};
  assign v_1988 = v_1989 | v_2004;
  assign v_1989 = v_1990 | v_1997;
  assign v_1990 = v_1991 | v_1994;
  assign v_1991 = v_1992 | v_1993;
  assign v_1992 = v_121 & v_177;
  assign v_1993 = v_123 & v_177;
  assign v_1994 = v_1995 | v_1996;
  assign v_1995 = v_139 & v_177;
  assign v_1996 = v_40 & v_177;
  assign v_1997 = v_1998 | v_2001;
  assign v_1998 = v_1999 | v_2000;
  assign v_1999 = v_153 & v_87;
  assign v_2000 = v_159 & v_749;
  assign v_2001 = v_2002 | v_2003;
  assign v_2002 = v_195 & v_749;
  assign v_2003 = v_203 & v_749;
  assign v_2004 = v_2005 | v_2012;
  assign v_2005 = v_2006 | v_2009;
  assign v_2006 = v_2007 | v_2008;
  assign v_2007 = v_208 & v_177;
  assign v_2008 = v_218 & v_177;
  assign v_2009 = v_2010 | v_2011;
  assign v_2010 = v_227 & v_177;
  assign v_2011 = v_233 & v_177;
  assign v_2012 = v_2013 | v_2016;
  assign v_2013 = v_2014 | v_2015;
  assign v_2014 = v_242 & v_177;
  assign v_2015 = v_244 & v_177;
  assign v_2016 = v_2017 | v_2018;
  assign v_2017 = v_252 & v_87;
  assign v_2018 = v_254 & v_87;
  assign v_2019 = {v_2020, v_2051};
  assign v_2020 = v_2021 | v_2036;
  assign v_2021 = v_2022 | v_2029;
  assign v_2022 = v_2023 | v_2026;
  assign v_2023 = v_2024 | v_2025;
  assign v_2024 = v_121 & v_177;
  assign v_2025 = v_123 & v_177;
  assign v_2026 = v_2027 | v_2028;
  assign v_2027 = v_139 & v_177;
  assign v_2028 = v_40 & v_177;
  assign v_2029 = v_2030 | v_2033;
  assign v_2030 = v_2031 | v_2032;
  assign v_2031 = v_153 & v_762;
  assign v_2032 = v_159 & v_749;
  assign v_2033 = v_2034 | v_2035;
  assign v_2034 = v_195 & v_749;
  assign v_2035 = v_203 & v_749;
  assign v_2036 = v_2037 | v_2044;
  assign v_2037 = v_2038 | v_2041;
  assign v_2038 = v_2039 | v_2040;
  assign v_2039 = v_208 & v_177;
  assign v_2040 = v_218 & v_177;
  assign v_2041 = v_2042 | v_2043;
  assign v_2042 = v_227 & v_177;
  assign v_2043 = v_233 & v_177;
  assign v_2044 = v_2045 | v_2048;
  assign v_2045 = v_2046 | v_2047;
  assign v_2046 = v_242 & v_177;
  assign v_2047 = v_244 & v_177;
  assign v_2048 = v_2049 | v_2050;
  assign v_2049 = v_252 & 1'h0;
  assign v_2050 = v_254 & 1'h0;
  assign v_2051 = {v_2052, v_2083};
  assign v_2052 = v_2053 | v_2068;
  assign v_2053 = v_2054 | v_2061;
  assign v_2054 = v_2055 | v_2058;
  assign v_2055 = v_2056 | v_2057;
  assign v_2056 = v_121 & v_191;
  assign v_2057 = v_123 & v_191;
  assign v_2058 = v_2059 | v_2060;
  assign v_2059 = v_139 & v_191;
  assign v_2060 = v_40 & v_191;
  assign v_2061 = v_2062 | v_2065;
  assign v_2062 = v_2063 | v_2064;
  assign v_2063 = v_153 & v_191;
  assign v_2064 = v_159 & v_749;
  assign v_2065 = v_2066 | v_2067;
  assign v_2066 = v_195 & v_749;
  assign v_2067 = v_203 & v_749;
  assign v_2068 = v_2069 | v_2076;
  assign v_2069 = v_2070 | v_2073;
  assign v_2070 = v_2071 | v_2072;
  assign v_2071 = v_208 & v_191;
  assign v_2072 = v_218 & v_191;
  assign v_2073 = v_2074 | v_2075;
  assign v_2074 = v_227 & v_191;
  assign v_2075 = v_233 & v_191;
  assign v_2076 = v_2077 | v_2080;
  assign v_2077 = v_2078 | v_2079;
  assign v_2078 = v_242 & v_191;
  assign v_2079 = v_244 & v_191;
  assign v_2080 = v_2081 | v_2082;
  assign v_2081 = v_252 & 1'h0;
  assign v_2082 = v_254 & 1'h0;
  assign v_2083 = {v_2084, v_2115};
  assign v_2084 = v_2085 | v_2100;
  assign v_2085 = v_2086 | v_2093;
  assign v_2086 = v_2087 | v_2090;
  assign v_2087 = v_2088 | v_2089;
  assign v_2088 = v_121 & v_179;
  assign v_2089 = v_123 & v_179;
  assign v_2090 = v_2091 | v_2092;
  assign v_2091 = v_139 & v_179;
  assign v_2092 = v_40 & v_179;
  assign v_2093 = v_2094 | v_2097;
  assign v_2094 = v_2095 | v_2096;
  assign v_2095 = v_153 & v_179;
  assign v_2096 = v_159 & v_749;
  assign v_2097 = v_2098 | v_2099;
  assign v_2098 = v_195 & v_749;
  assign v_2099 = v_203 & v_749;
  assign v_2100 = v_2101 | v_2108;
  assign v_2101 = v_2102 | v_2105;
  assign v_2102 = v_2103 | v_2104;
  assign v_2103 = v_208 & v_179;
  assign v_2104 = v_218 & v_179;
  assign v_2105 = v_2106 | v_2107;
  assign v_2106 = v_227 & v_179;
  assign v_2107 = v_233 & v_179;
  assign v_2108 = v_2109 | v_2112;
  assign v_2109 = v_2110 | v_2111;
  assign v_2110 = v_242 & v_179;
  assign v_2111 = v_244 & v_179;
  assign v_2112 = v_2113 | v_2114;
  assign v_2113 = v_252 & 1'h0;
  assign v_2114 = v_254 & 1'h0;
  assign v_2115 = {v_2116, v_2147};
  assign v_2116 = v_2117 | v_2132;
  assign v_2117 = v_2118 | v_2125;
  assign v_2118 = v_2119 | v_2122;
  assign v_2119 = v_2120 | v_2121;
  assign v_2120 = v_121 & v_181;
  assign v_2121 = v_123 & v_181;
  assign v_2122 = v_2123 | v_2124;
  assign v_2123 = v_139 & v_181;
  assign v_2124 = v_40 & v_181;
  assign v_2125 = v_2126 | v_2129;
  assign v_2126 = v_2127 | v_2128;
  assign v_2127 = v_153 & v_181;
  assign v_2128 = v_159 & v_749;
  assign v_2129 = v_2130 | v_2131;
  assign v_2130 = v_195 & v_749;
  assign v_2131 = v_203 & v_749;
  assign v_2132 = v_2133 | v_2140;
  assign v_2133 = v_2134 | v_2137;
  assign v_2134 = v_2135 | v_2136;
  assign v_2135 = v_208 & v_181;
  assign v_2136 = v_218 & v_181;
  assign v_2137 = v_2138 | v_2139;
  assign v_2138 = v_227 & v_181;
  assign v_2139 = v_233 & v_181;
  assign v_2140 = v_2141 | v_2144;
  assign v_2141 = v_2142 | v_2143;
  assign v_2142 = v_242 & v_181;
  assign v_2143 = v_244 & v_181;
  assign v_2144 = v_2145 | v_2146;
  assign v_2145 = v_252 & 1'h0;
  assign v_2146 = v_254 & 1'h0;
  assign v_2147 = {v_2148, v_2179};
  assign v_2148 = v_2149 | v_2164;
  assign v_2149 = v_2150 | v_2157;
  assign v_2150 = v_2151 | v_2154;
  assign v_2151 = v_2152 | v_2153;
  assign v_2152 = v_121 & v_183;
  assign v_2153 = v_123 & v_183;
  assign v_2154 = v_2155 | v_2156;
  assign v_2155 = v_139 & v_183;
  assign v_2156 = v_40 & v_183;
  assign v_2157 = v_2158 | v_2161;
  assign v_2158 = v_2159 | v_2160;
  assign v_2159 = v_153 & v_183;
  assign v_2160 = v_159 & v_749;
  assign v_2161 = v_2162 | v_2163;
  assign v_2162 = v_195 & v_749;
  assign v_2163 = v_203 & v_749;
  assign v_2164 = v_2165 | v_2172;
  assign v_2165 = v_2166 | v_2169;
  assign v_2166 = v_2167 | v_2168;
  assign v_2167 = v_208 & v_183;
  assign v_2168 = v_218 & v_183;
  assign v_2169 = v_2170 | v_2171;
  assign v_2170 = v_227 & v_183;
  assign v_2171 = v_233 & v_183;
  assign v_2172 = v_2173 | v_2176;
  assign v_2173 = v_2174 | v_2175;
  assign v_2174 = v_242 & v_183;
  assign v_2175 = v_244 & v_183;
  assign v_2176 = v_2177 | v_2178;
  assign v_2177 = v_252 & 1'h0;
  assign v_2178 = v_254 & 1'h0;
  assign v_2179 = {v_2180, v_2211};
  assign v_2180 = v_2181 | v_2196;
  assign v_2181 = v_2182 | v_2189;
  assign v_2182 = v_2183 | v_2186;
  assign v_2183 = v_2184 | v_2185;
  assign v_2184 = v_121 & v_185;
  assign v_2185 = v_123 & v_185;
  assign v_2186 = v_2187 | v_2188;
  assign v_2187 = v_139 & v_185;
  assign v_2188 = v_40 & v_185;
  assign v_2189 = v_2190 | v_2193;
  assign v_2190 = v_2191 | v_2192;
  assign v_2191 = v_153 & v_185;
  assign v_2192 = v_159 & v_749;
  assign v_2193 = v_2194 | v_2195;
  assign v_2194 = v_195 & v_749;
  assign v_2195 = v_203 & v_749;
  assign v_2196 = v_2197 | v_2204;
  assign v_2197 = v_2198 | v_2201;
  assign v_2198 = v_2199 | v_2200;
  assign v_2199 = v_208 & v_185;
  assign v_2200 = v_218 & v_185;
  assign v_2201 = v_2202 | v_2203;
  assign v_2202 = v_227 & v_185;
  assign v_2203 = v_233 & v_185;
  assign v_2204 = v_2205 | v_2208;
  assign v_2205 = v_2206 | v_2207;
  assign v_2206 = v_242 & v_185;
  assign v_2207 = v_244 & v_185;
  assign v_2208 = v_2209 | v_2210;
  assign v_2209 = v_252 & 1'h0;
  assign v_2210 = v_254 & 1'h0;
  assign v_2211 = {v_2212, v_2243};
  assign v_2212 = v_2213 | v_2228;
  assign v_2213 = v_2214 | v_2221;
  assign v_2214 = v_2215 | v_2218;
  assign v_2215 = v_2216 | v_2217;
  assign v_2216 = v_121 & v_187;
  assign v_2217 = v_123 & v_187;
  assign v_2218 = v_2219 | v_2220;
  assign v_2219 = v_139 & v_187;
  assign v_2220 = v_40 & v_187;
  assign v_2221 = v_2222 | v_2225;
  assign v_2222 = v_2223 | v_2224;
  assign v_2223 = v_153 & v_187;
  assign v_2224 = v_159 & v_749;
  assign v_2225 = v_2226 | v_2227;
  assign v_2226 = v_195 & v_749;
  assign v_2227 = v_203 & v_749;
  assign v_2228 = v_2229 | v_2236;
  assign v_2229 = v_2230 | v_2233;
  assign v_2230 = v_2231 | v_2232;
  assign v_2231 = v_208 & v_187;
  assign v_2232 = v_218 & v_187;
  assign v_2233 = v_2234 | v_2235;
  assign v_2234 = v_227 & v_187;
  assign v_2235 = v_233 & v_187;
  assign v_2236 = v_2237 | v_2240;
  assign v_2237 = v_2238 | v_2239;
  assign v_2238 = v_242 & v_187;
  assign v_2239 = v_244 & v_187;
  assign v_2240 = v_2241 | v_2242;
  assign v_2241 = v_252 & 1'h0;
  assign v_2242 = v_254 & 1'h0;
  assign v_2243 = {v_2244, v_2276};
  assign v_2244 = v_2245 | v_2261;
  assign v_2245 = v_2246 | v_2254;
  assign v_2246 = v_2247 | v_2251;
  assign v_2247 = v_2248 | v_2249;
  assign v_2248 = v_121 & v_749;
  assign v_2249 = v_123 & v_2250;
  assign v_2250 = v_51[11:11];
  assign v_2251 = v_2252 | v_2253;
  assign v_2252 = v_139 & v_749;
  assign v_2253 = v_40 & v_749;
  assign v_2254 = v_2255 | v_2258;
  assign v_2255 = v_2256 | v_2257;
  assign v_2256 = v_153 & v_749;
  assign v_2257 = v_159 & v_749;
  assign v_2258 = v_2259 | v_2260;
  assign v_2259 = v_195 & v_749;
  assign v_2260 = v_203 & v_749;
  assign v_2261 = v_2262 | v_2269;
  assign v_2262 = v_2263 | v_2266;
  assign v_2263 = v_2264 | v_2265;
  assign v_2264 = v_208 & v_749;
  assign v_2265 = v_218 & v_749;
  assign v_2266 = v_2267 | v_2268;
  assign v_2267 = v_227 & v_749;
  assign v_2268 = v_233 & v_749;
  assign v_2269 = v_2270 | v_2273;
  assign v_2270 = v_2271 | v_2272;
  assign v_2271 = v_242 & v_749;
  assign v_2272 = v_244 & v_749;
  assign v_2273 = v_2274 | v_2275;
  assign v_2274 = v_252 & 1'h0;
  assign v_2275 = v_254 & 1'h0;
  assign v_2276 = {v_2277, v_2309};
  assign v_2277 = v_2278 | v_2294;
  assign v_2278 = v_2279 | v_2287;
  assign v_2279 = v_2280 | v_2284;
  assign v_2280 = v_2281 | v_2282;
  assign v_2281 = v_121 & v_751;
  assign v_2282 = v_123 & v_2283;
  assign v_2283 = v_51[10:10];
  assign v_2284 = v_2285 | v_2286;
  assign v_2285 = v_139 & v_751;
  assign v_2286 = v_40 & v_751;
  assign v_2287 = v_2288 | v_2291;
  assign v_2288 = v_2289 | v_2290;
  assign v_2289 = v_153 & v_751;
  assign v_2290 = v_159 & v_751;
  assign v_2291 = v_2292 | v_2293;
  assign v_2292 = v_195 & v_751;
  assign v_2293 = v_203 & v_751;
  assign v_2294 = v_2295 | v_2302;
  assign v_2295 = v_2296 | v_2299;
  assign v_2296 = v_2297 | v_2298;
  assign v_2297 = v_208 & v_751;
  assign v_2298 = v_218 & v_751;
  assign v_2299 = v_2300 | v_2301;
  assign v_2300 = v_227 & v_751;
  assign v_2301 = v_233 & v_751;
  assign v_2302 = v_2303 | v_2306;
  assign v_2303 = v_2304 | v_2305;
  assign v_2304 = v_242 & v_751;
  assign v_2305 = v_244 & v_751;
  assign v_2306 = v_2307 | v_2308;
  assign v_2307 = v_252 & 1'h0;
  assign v_2308 = v_254 & 1'h0;
  assign v_2309 = {v_2310, v_2342};
  assign v_2310 = v_2311 | v_2327;
  assign v_2311 = v_2312 | v_2320;
  assign v_2312 = v_2313 | v_2317;
  assign v_2313 = v_2314 | v_2315;
  assign v_2314 = v_121 & v_753;
  assign v_2315 = v_123 & v_2316;
  assign v_2316 = v_51[9:9];
  assign v_2317 = v_2318 | v_2319;
  assign v_2318 = v_139 & v_753;
  assign v_2319 = v_40 & v_753;
  assign v_2320 = v_2321 | v_2324;
  assign v_2321 = v_2322 | v_2323;
  assign v_2322 = v_153 & v_753;
  assign v_2323 = v_159 & v_753;
  assign v_2324 = v_2325 | v_2326;
  assign v_2325 = v_195 & v_753;
  assign v_2326 = v_203 & v_753;
  assign v_2327 = v_2328 | v_2335;
  assign v_2328 = v_2329 | v_2332;
  assign v_2329 = v_2330 | v_2331;
  assign v_2330 = v_208 & v_753;
  assign v_2331 = v_218 & v_753;
  assign v_2332 = v_2333 | v_2334;
  assign v_2333 = v_227 & v_753;
  assign v_2334 = v_233 & v_753;
  assign v_2335 = v_2336 | v_2339;
  assign v_2336 = v_2337 | v_2338;
  assign v_2337 = v_242 & v_753;
  assign v_2338 = v_244 & v_753;
  assign v_2339 = v_2340 | v_2341;
  assign v_2340 = v_252 & 1'h0;
  assign v_2341 = v_254 & 1'h0;
  assign v_2342 = {v_2343, v_2375};
  assign v_2343 = v_2344 | v_2360;
  assign v_2344 = v_2345 | v_2353;
  assign v_2345 = v_2346 | v_2350;
  assign v_2346 = v_2347 | v_2348;
  assign v_2347 = v_121 & v_755;
  assign v_2348 = v_123 & v_2349;
  assign v_2349 = v_51[8:8];
  assign v_2350 = v_2351 | v_2352;
  assign v_2351 = v_139 & v_755;
  assign v_2352 = v_40 & v_755;
  assign v_2353 = v_2354 | v_2357;
  assign v_2354 = v_2355 | v_2356;
  assign v_2355 = v_153 & v_755;
  assign v_2356 = v_159 & v_755;
  assign v_2357 = v_2358 | v_2359;
  assign v_2358 = v_195 & v_755;
  assign v_2359 = v_203 & v_755;
  assign v_2360 = v_2361 | v_2368;
  assign v_2361 = v_2362 | v_2365;
  assign v_2362 = v_2363 | v_2364;
  assign v_2363 = v_208 & v_755;
  assign v_2364 = v_218 & v_755;
  assign v_2365 = v_2366 | v_2367;
  assign v_2366 = v_227 & v_755;
  assign v_2367 = v_233 & v_755;
  assign v_2368 = v_2369 | v_2372;
  assign v_2369 = v_2370 | v_2371;
  assign v_2370 = v_242 & v_755;
  assign v_2371 = v_244 & v_755;
  assign v_2372 = v_2373 | v_2374;
  assign v_2373 = v_252 & 1'h0;
  assign v_2374 = v_254 & 1'h0;
  assign v_2375 = v_2376 | v_2392;
  assign v_2376 = v_2377 | v_2385;
  assign v_2377 = v_2378 | v_2382;
  assign v_2378 = v_2379 | v_2380;
  assign v_2379 = v_121 & v_762;
  assign v_2380 = v_123 & v_2381;
  assign v_2381 = v_51[7:7];
  assign v_2382 = v_2383 | v_2384;
  assign v_2383 = v_139 & v_762;
  assign v_2384 = v_40 & v_762;
  assign v_2385 = v_2386 | v_2389;
  assign v_2386 = v_2387 | v_2388;
  assign v_2387 = v_153 & 1'h0;
  assign v_2388 = v_159 & v_762;
  assign v_2389 = v_2390 | v_2391;
  assign v_2390 = v_195 & v_762;
  assign v_2391 = v_203 & v_762;
  assign v_2392 = v_2393 | v_2400;
  assign v_2393 = v_2394 | v_2397;
  assign v_2394 = v_2395 | v_2396;
  assign v_2395 = v_208 & v_762;
  assign v_2396 = v_218 & v_762;
  assign v_2397 = v_2398 | v_2399;
  assign v_2398 = v_227 & v_762;
  assign v_2399 = v_233 & v_762;
  assign v_2400 = v_2401 | v_2404;
  assign v_2401 = v_2402 | v_2403;
  assign v_2402 = v_242 & v_762;
  assign v_2403 = v_244 & v_762;
  assign v_2404 = v_2405 | v_2406;
  assign v_2405 = v_252 & 1'h0;
  assign v_2406 = v_254 & 1'h0;
  assign v_2407 = v_395 | v_701;
  assign v_2408 = v_2409 | v_2410;
  assign v_2409 = v_779 | v_796;
  assign v_2410 = v_815 | v_834;
  assign v_2411 = v_2412 | v_2415;
  assign v_2412 = v_2413 | v_2414;
  assign v_2413 = v_867 | v_890;
  assign v_2414 = v_909 | v_924;
  assign v_2415 = v_2416 | v_2417;
  assign v_2416 = v_944 | v_964;
  assign v_2417 = v_984 | v_1038;
  assign v_2418 = v_2419 == v_2428;
  assign v_2419 = {v_2420, v_2421};
  assign v_2420 = v_104[11:11];
  assign v_2421 = {v_2422, v_2423};
  assign v_2422 = v_104[10:10];
  assign v_2423 = {v_2424, v_2425};
  assign v_2424 = v_104[9:9];
  assign v_2425 = {v_2426, v_2427};
  assign v_2426 = v_104[8:8];
  assign v_2427 = v_104[7:7];
  assign v_2428 = {v_2429, v_2430};
  assign v_2429 = v_51[19:19];
  assign v_2430 = {v_2431, v_2432};
  assign v_2431 = v_51[18:18];
  assign v_2432 = {v_2433, v_2434};
  assign v_2433 = v_51[17:17];
  assign v_2434 = {v_2435, v_2436};
  assign v_2435 = v_51[16:16];
  assign v_2436 = v_51[15:15];
  assign v_2437 = mux_2437(v_2438);
  assign v_2438 = act_280 & v_2439;
  assign v_2439 = v_2440 == v_2449;
  assign v_2440 = {v_2441, v_2442};
  assign v_2441 = v_288[11:11];
  assign v_2442 = {v_2443, v_2444};
  assign v_2443 = v_288[10:10];
  assign v_2444 = {v_2445, v_2446};
  assign v_2445 = v_288[9:9];
  assign v_2446 = {v_2447, v_2448};
  assign v_2447 = v_288[8:8];
  assign v_2448 = v_288[7:7];
  assign v_2449 = {v_2450, v_2451};
  assign v_2450 = v_51[19:19];
  assign v_2451 = {v_2452, v_2453};
  assign v_2452 = v_51[18:18];
  assign v_2453 = {v_2454, v_2455};
  assign v_2454 = v_51[17:17];
  assign v_2455 = {v_2456, v_2457};
  assign v_2456 = v_51[16:16];
  assign v_2457 = v_51[15:15];
  assign v_2458 = mux_2458(v_2459);
  assign v_2459 = v_2460 & v_2463;
  assign v_2460 = v_2461 & v_2462;
  assign v_2463 = v_2464 == v_2488;
  assign v_2465 = v_2466 | v_2486;
  assign v_2466 = mux_2466(1'h1);
  assign v_2467 = mux_2467(v_3);
  assign v_2468 = {v_2469, v_2470};
  assign v_2469 = v_52[19:19];
  assign v_2470 = {v_2471, v_2472};
  assign v_2471 = v_52[18:18];
  assign v_2472 = {v_2473, v_2474};
  assign v_2473 = v_52[17:17];
  assign v_2474 = {v_2475, v_2476};
  assign v_2475 = v_52[16:16];
  assign v_2476 = v_52[15:15];
  assign v_2477 = {v_2478, v_2479};
  assign v_2478 = v_51[19:19];
  assign v_2479 = {v_2480, v_2481};
  assign v_2480 = v_51[18:18];
  assign v_2481 = {v_2482, v_2483};
  assign v_2482 = v_51[17:17];
  assign v_2483 = {v_2484, v_2485};
  assign v_2484 = v_51[16:16];
  assign v_2485 = v_51[15:15];
  assign v_2486 = mux_2486(v_2487);
  assign v_2487 = ~1'h1;
  assign v_2489 = v_2490 | v_2491;
  assign v_2490 = mux_2490(act_333);
  assign v_2491 = mux_2491(v_2492);
  assign v_2492 = ~act_333;
  BlockRAMDual#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(5), .DATA_WIDTH(32))
    ram2493
      (.CLK(clock),
       .RD_ADDR(v_2494),
       .WR_ADDR(v_2498),
       .DI(v_2502),
       .WE(v_2506),
       .RE(v_2510),
       .DO(v_2493));
  assign v_2494 = v_2495 | v_2496;
  assign v_2495 = mux_2495(1'h1);
  assign v_2496 = mux_2496(v_2497);
  assign v_2497 = ~1'h1;
  assign v_2498 = v_2499 | v_2500;
  assign v_2499 = mux_2499(act_333);
  assign v_2500 = mux_2500(v_2501);
  assign v_2501 = ~act_333;
  assign v_2502 = v_2503 | v_2504;
  assign v_2503 = mux_2503(act_333);
  assign v_2504 = mux_2504(v_2505);
  assign v_2505 = ~act_333;
  assign v_2506 = v_2507 | v_2508;
  assign v_2507 = mux_2507(act_333);
  assign v_2508 = mux_2508(v_2509);
  assign v_2509 = ~act_333;
  assign v_2510 = mux_2510(v_2511);
  assign v_2511 = ~1'h0;
  assign v_2513 = v_2514 | v_2515;
  assign v_2514 = mux_2514(act_333);
  assign v_2515 = mux_2515(v_2516);
  assign v_2516 = ~act_333;
  assign v_2517 = v_2518 & v_2522;
  assign v_2518 = v_2519 | 1'h0;
  assign v_2520 = v_122 & v_2521;
  assign v_2521 = ~v_89;
  assign v_2522 = ~v_90;
  assign v_2523 = v_2524 | v_2532;
  assign v_2524 = v_2525 & v_1007;
  assign v_2525 = v_2526 | v_2531;
  assign v_2527 = v_2528 & v_2530;
  assign v_2528 = v_2529 & v_85;
  assign v_2529 = v_211 & v_84;
  assign v_2530 = ~v_89;
  assign v_2531 = v_1014 | 1'h0;
  assign v_2532 = v_2533 & v_2541;
  assign v_2533 = v_2534 | v_2540;
  assign v_2535 = v_2536 & v_2539;
  assign v_2536 = v_2537 & v_85;
  assign v_2537 = v_2538 & v_84;
  assign v_2538 = v_212 & v_87;
  assign v_2539 = ~v_89;
  assign v_2540 = v_1020 | 1'h0;
  assign v_2541 = ~v_1007;
  assign v_2542 = v_831 + v_2543;
  assign v_2543 = {v_2544, v_2545};
  assign v_2545 = {v_2544, v_2546};
  assign v_2546 = {v_2544, v_2547};
  assign v_2547 = {v_2544, v_2548};
  assign v_2548 = {v_2544, v_2549};
  assign v_2549 = {v_2544, v_2550};
  assign v_2550 = {v_2544, v_2551};
  assign v_2551 = {v_2544, v_2552};
  assign v_2552 = {v_2544, v_2553};
  assign v_2553 = {v_2544, v_2554};
  assign v_2554 = {v_2544, v_2555};
  assign v_2555 = {v_2544, v_2556};
  assign v_2556 = {v_2544, v_2557};
  assign v_2557 = {v_2544, v_2558};
  assign v_2558 = {v_2544, v_2559};
  assign v_2559 = {v_2544, v_2560};
  assign v_2560 = {v_2544, v_2561};
  assign v_2561 = {v_2544, v_2562};
  assign v_2562 = {v_2544, v_2563};
  assign v_2563 = {v_2544, v_2564};
  assign v_2564 = {v_2565, v_2566};
  assign v_2566 = {v_2567, v_2568};
  assign v_2568 = {v_2569, v_2570};
  assign v_2570 = {v_2571, v_2572};
  assign v_2572 = {v_2573, v_2574};
  assign v_2574 = {v_2575, v_2576};
  assign v_2576 = {v_2577, v_2578};
  assign v_2578 = {v_2579, v_2580};
  assign v_2580 = {v_2581, v_2582};
  assign v_2582 = {v_2583, v_2584};
  assign v_2584 = {v_2585, v_2586};
  assign v_2587 = mux_2587(v_2588);
  assign v_2588 = ~act_35;
  assign v_2589 = v_2590 | v_2593;
  assign v_2590 = v_2591 | v_2592;
  assign v_2591 = mux_2591(v_766);
  assign v_2592 = mux_2592(v_716);
  assign v_2593 = v_2594 | v_2598;
  assign v_2594 = mux_2594(v_37);
  assign v_2595 = {v_2596, 1'h0};
  assign v_2596 = v_2597[31:1];
  assign v_2597 = v_91 + v_115;
  assign v_2598 = mux_2598(v_2599);
  assign v_2599 = v_2600 & v_411;
  assign v_2600 = v_828 | 1'h0;
  assign v_2601 = v_831 + v_115;
  assign v_2602 = mux_2602(v_2603);
  assign v_2603 = ~1'h1;
  assign v_2604 = mux_2604(v_2605);
  assign v_2605 = ~1'h0;
  assign v_2606 = mux_2606(v_2607);
  assign v_2607 = ~1'h0;
  assign v_2608 = v_2609 | v_2611;
  assign v_2609 = mux_2609(v_2610);
  assign v_2610 = 1'h1 & v_3;
  assign v_2611 = mux_2611(v_2612);
  assign v_2612 = ~v_2610;
  assign v_2613 = ~v_135;
  assign v_2614 = ~v_81;
  assign v_2615 = ~v_83;
  assign v_2616 = ~v_87;
  assign v_2617 = ~v_89;
  assign v_2618 = v_65 | v_2619;
  assign v_2619 = v_766 | v_716;
  assign v_2620 = 1'h1 & act_35;
  assign v_2621 = v_2622 | v_2624;
  assign v_2622 = mux_2622(v_31);
  assign v_2624 = mux_2624(v_2620);
  assign v_2625 = v_639 & v_81;
  assign v_2626 = mux_2626(v_2627);
  assign v_2627 = ~v_25;
  assign v_2629 = mux_2629(v_2630);
  assign v_2630 = ~1'h1;
  assign v_2631 = ~v_1321;
  assign v_2632 = v_2633 | v_2634;
  assign v_2633 = mux_2633(v_15);
  assign v_2634 = mux_2634(v_16);
  assign v_2635 = v_426 | v_420;
  assign v_2636 = v_634 | v_2637;
  assign v_2637 = v_2638 & act_436;
  assign v_2638 = ~v_482;
  assign v_2639 = v_2640 | v_2643;
  assign v_2640 = v_2641 | v_2642;
  assign v_2641 = mux_2641(v_11);
  assign v_2642 = mux_2642(v_25);
  assign v_2643 = v_2644 | v_2645;
  assign v_2644 = mux_2644(v_634);
  assign v_2645 = mux_2645(v_2637);
  assign v_2646 = 1'h1 & v_2647;
  assign v_2647 = ~v_12;
  assign v_2648 = mux_2648(v_417);
  assign v_2649 = v_2650 | v_2651;
  assign v_2650 = mux_2650(v_25);
  assign v_2651 = mux_2651(v_667);
  assign v_2652 = v_2653 | v_2656;
  assign v_2653 = v_2654 | v_2655;
  assign v_2654 = mux_2654(v_634);
  assign v_2655 = mux_2655(v_671);
  assign v_2656 = v_2657 | v_2658;
  assign v_2657 = mux_2657(v_2637);
  assign v_2658 = mux_2658(v_2659);
  assign v_2659 = ~v_2660;
  assign v_2660 = v_2661 | v_2663;
  assign v_2661 = v_2637 | v_2662;
  assign v_2662 = v_7 | v_417;
  assign v_2663 = v_2664 | v_2665;
  assign v_2664 = v_25 | v_667;
  assign v_2665 = v_634 | v_671;
  assign v_2667 = v_2668 & v_408;
  assign v_2668 = v_685 == 12'h800;
  assign v_2670 = v_2669 + 32'h1;
  assign v_2672 = v_2673 & v_408;
  assign v_2673 = v_685 == 12'h801;
  assign in0_consume_en = v_2675;
  assign v_2675 = v_2676 | v_2677;
  assign v_2676 = mux_2676(v_112);
  assign v_2677 = mux_2677(v_2678);
  assign v_2678 = ~v_112;
  assign out_canPeek = v_680;
  assign out_peek = v_2681;
  assign v_2682 = v_2683 | v_2685;
  assign v_2683 = mux_2683(act_683);
  assign v_2684 = v_91[7:0];
  assign v_2685 = mux_2685(v_2686);
  assign v_2686 = ~act_683;
  // Always block
  //////////////////////////////////////////////////////////////////////////////
  always @(posedge clock) begin
    if (reset) begin
      v_8 <= 1'h0;
      v_13 <= 1'h0;
      v_21 <= 1'h0;
      v_22 <= 1'h0;
      v_28 <= 1'h0;
      v_29 <= 1'h0;
      v_39 <= 1'h0;
      v_51 <= 32'h0;
      v_59 <= 32'hfffffffc;
      v_70 <= 1'h0;
      v_91 <= 32'h0;
      v_104 <= 32'h0;
      v_115 <= 32'h0;
      v_288 <= 32'h0;
      v_290 <= 1'h0;
      v_307 <= 1'h0;
      v_331 <= 1'h0;
      v_332 <= 1'h0;
      v_335 <= 5'h0;
      v_359 <= 5'h0;
      v_389 <= 32'h0;
      v_410 <= 1'h0;
      v_413 <= 1'h0;
      v_420 <= 1'h0;
      v_426 <= 1'h0;
      v_439 <= 1'h0;
      v_441 <= 1'h0;
      v_490 <= 1'h0;
      v_491 <= 1'h0;
      v_517 <= 32'h0;
      v_535 <= 1'h0;
      v_637 <= 1'h0;
      v_680 <= 1'h0;
      v_714 <= 32'h0;
      v_718 <= 1'h0;
      v_768 <= 1'h0;
      v_792 <= 32'h0;
      v_809 <= 32'h0;
      v_828 <= 1'h0;
      v_831 <= 32'h0;
      v_832 <= 32'h0;
      v_847 <= 1'h0;
      v_855 <= 1'h0;
      v_880 <= 1'h0;
      v_903 <= 1'h0;
      v_922 <= 1'h0;
      v_937 <= 1'h0;
      v_957 <= 1'h0;
      v_977 <= 1'h0;
      v_997 <= 1'h0;
      v_1003 <= 1'h0;
      v_1014 <= 1'h0;
      v_1020 <= 1'h0;
      v_1028 <= 1'h0;
      v_1052 <= 1'h0;
      v_1097 <= 73'h0;
      v_1108 <= 1'h0;
      v_1109 <= 1'h0;
      v_1139 <= 64'h0;
      v_1156 <= 78'h0;
      v_1283 <= 6'h0;
      v_1284 <= 32'h0;
      v_1286 <= 1'h0;
      v_1290 <= 1'h0;
      v_1294 <= 1'h0;
      v_1295 <= 1'h0;
      v_1298 <= 32'h0;
      v_1311 <= 1'h0;
      v_1315 <= 32'h0;
      v_1322 <= 6'h0;
      v_1337 <= 32'h0;
      v_1347 <= 32'h0;
      v_1369 <= 32'h0;
      v_2461 <= 1'h0;
      v_2462 <= 1'h0;
      v_2464 <= 5'h0;
      v_2488 <= 5'h0;
      v_2512 <= 32'h0;
      v_2519 <= 1'h0;
      v_2526 <= 1'h0;
      v_2534 <= 1'h0;
      v_2544 <= 1'h0;
      v_2565 <= 1'h0;
      v_2567 <= 1'h0;
      v_2569 <= 1'h0;
      v_2571 <= 1'h0;
      v_2573 <= 1'h0;
      v_2575 <= 1'h0;
      v_2577 <= 1'h0;
      v_2579 <= 1'h0;
      v_2581 <= 1'h0;
      v_2583 <= 1'h0;
      v_2585 <= 1'h0;
      v_2586 <= 1'h0;
      v_2623 <= 1'h0;
      v_2628 <= 1'h0;
      v_2669 <= 32'h0;
      v_2681 <= 8'h0;
    end else begin
      if (v_1 == 1) $write
        ("Pipeline assertion failed: simultaneous stall and flush", "\n");
      if (v_9 == 1) v_8 <= v_2639;
      if (v_14 == 1) v_13 <= v_2632;
      v_21 <= v_22;
      if (1'h1 == 1) v_22 <= v_23;
      if (v_29 == 1) v_28 <= v_2625;
      if (v_30 == 1) v_29 <= v_2621;
      if (v_29 == 1) v_39 <= v_40;
      if (v_31 == 1) v_51 <= v_52;
      if (v_60 == 1) v_59 <= v_57;
      if (v_29 == 1) v_70 <= v_71;
      if (v_92 == 1) v_91 <= v_94;
      if (v_92 == 1) v_104 <= v_51;
      if (v_92 == 1) v_115 <= v_116;
      if (v_289 == 1) v_288 <= v_104;
      if (v_291 == 1) v_290 <= v_295;
      v_307 <= act_96;
      v_331 <= 1'h1;
      v_332 <= act_333;
      v_335 <= v_336;
      v_359 <= v_360;
      v_389 <= v_390;
      if (v_29 == 1) v_410 <= v_121;
      if (1'h1 == 1) v_413 <= v_414;
      if (v_421 == 1) v_420 <= v_663;
      if (1'h1 == 1) v_426 <= v_427;
      if (v_29 == 1) v_439 <= v_139;
      if (v_29 == 1) v_441 <= v_123;
      if (v_29 == 1) v_490 <= v_83;
      if (v_29 == 1) v_491 <= v_87;
      if (v_92 == 1) v_517 <= v_257;
      if (v_29 == 1) v_535 <= v_81;
      if (v_29 == 1) v_637 <= v_638;
      if (v_681 == 1) v_680 <= v_697;
      if (v_715 == 1) v_714 <= v_770;
      if (v_29 == 1) v_718 <= v_719;
      if (v_29 == 1) v_768 <= v_769;
      if (v_793 == 1) v_792 <= v_91;
      if (v_810 == 1) v_809 <= v_91;
      if (v_29 == 1) v_828 <= v_153;
      if (v_92 == 1) v_831 <= v_832;
      if (v_31 == 1) v_832 <= v_59;
      if (v_29 == 1) v_847 <= v_848;
      if (v_29 == 1) v_855 <= v_856;
      if (v_29 == 1) v_880 <= v_881;
      if (v_29 == 1) v_903 <= v_252;
      if (v_29 == 1) v_922 <= v_254;
      if (v_29 == 1) v_937 <= v_938;
      if (v_29 == 1) v_957 <= v_958;
      if (v_29 == 1) v_977 <= v_978;
      if (v_29 == 1) v_997 <= v_998;
      if (v_29 == 1) v_1003 <= v_1004;
      if (v_29 == 1) v_1014 <= v_1015;
      if (v_29 == 1) v_1020 <= v_1021;
      if (v_29 == 1) v_1028 <= v_1029;
      if (v_29 == 1) v_1052 <= v_1053;
      if (v_634 == 1) v_1097 <= v_1098;
      if (v_29 == 1) v_1108 <= v_83;
      if (v_29 == 1) v_1109 <= v_87;
      if (v_634 == 1) v_1139 <= v_1140;
      if (v_1157 == 1) v_1156 <= v_1158;
      if (v_25 == 1) v_1283 <= 6'bxxxxxx;
      if (v_16 == 1) v_1284 <= v_1285;
      if (v_1287 == 1) v_1286 <= v_1288;
      if (v_25 == 1) v_1290 <= v_1291;
      if (v_29 == 1) v_1294 <= v_83;
      if (v_29 == 1) v_1295 <= v_87;
      if (v_1299 == 1) v_1298 <= v_1305;
      if (v_25 == 1) v_1311 <= v_1312;
      if (v_1316 == 1) v_1315 <= v_1328;
      if (v_1323 == 1) v_1322 <= v_1324;
      if (v_1338 == 1) v_1337 <= v_1339;
      if (v_1348 == 1) v_1347 <= v_1349;
      v_1369 <= v_1370;
      v_2461 <= 1'h1;
      v_2462 <= act_333;
      v_2464 <= v_2465;
      v_2488 <= v_2489;
      v_2512 <= v_2513;
      if (v_29 == 1) v_2519 <= v_2520;
      if (v_29 == 1) v_2526 <= v_2527;
      if (v_29 == 1) v_2534 <= v_2535;
      if (v_29 == 1) v_2544 <= v_177;
      if (v_29 == 1) v_2565 <= v_2381;
      if (v_29 == 1) v_2567 <= v_191;
      if (v_29 == 1) v_2569 <= v_179;
      if (v_29 == 1) v_2571 <= v_181;
      if (v_29 == 1) v_2573 <= v_183;
      if (v_29 == 1) v_2575 <= v_185;
      if (v_29 == 1) v_2577 <= v_187;
      if (v_29 == 1) v_2579 <= v_2250;
      if (v_29 == 1) v_2581 <= v_2283;
      if (v_29 == 1) v_2583 <= v_2316;
      if (v_29 == 1) v_2585 <= v_2349;
      if (v_29 == 1) v_2586 <= 1'h0;
      v_2623 <= 1'h1;
      v_2628 <= v_1320;
      if (v_2667 == 1) $write (v_2669, ": 0x%08x", v_91, "\n");
      if (1'h1 == 1) v_2669 <= v_2670;
      if (v_2672 == 1) $finish;
      if (v_682 == 1) v_2681 <= v_2682;
    end
  end
endmodule