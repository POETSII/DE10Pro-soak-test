module Pebbles
  (input wire clock,
   input wire reset,
   input wire [0:0] out_consume_en,
   input wire [0:0] in0_canPeek,
   input wire [7:0] in0_peek,
   output wire [0:0] in0_consume_en,
   output wire [0:0] out_canPeek,
   output wire [7:0] out_peek);
  // Declarations
  //////////////////////////////////////////////////////////////////////////////
  wire [0:0] v_0;
  wire [0:0] v_1;
  function [0:0] mux_1(input [0:0] sel);
    case (sel) 0: mux_1 = 1'h0; 1: mux_1 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2;
  wire [0:0] vin0_consume_en_3;
  wire [0:0] vout_canPeek_3;
  wire [7:0] vout_peek_3;
  wire [0:0] v_4;
  function [0:0] mux_4(input [0:0] sel);
    case (sel) 0: mux_4 = 1'h0; 1: mux_4 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5;
  wire [0:0] v_6;
  wire [0:0] v_7;
  function [0:0] mux_7(input [0:0] sel);
    case (sel) 0: mux_7 = 1'h0; 1: mux_7 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8;
  wire [0:0] v_9;
  wire [0:0] v_10;
  wire [0:0] vin0_consume_en_11;
  wire [0:0] vout_canPeek_11;
  wire [7:0] vout_peek_11;
  wire [0:0] v_12;
  function [0:0] mux_12(input [0:0] sel);
    case (sel) 0: mux_12 = 1'h0; 1: mux_12 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13;
  wire [0:0] v_14;
  wire [0:0] v_15;
  function [0:0] mux_15(input [0:0] sel);
    case (sel) 0: mux_15 = 1'h0; 1: mux_15 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16;
  wire [0:0] vin0_consume_en_17;
  wire [0:0] vout_canPeek_17;
  wire [7:0] vout_peek_17;
  wire [0:0] v_18;
  function [0:0] mux_18(input [0:0] sel);
    case (sel) 0: mux_18 = 1'h0; 1: mux_18 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19;
  wire [0:0] v_20;
  wire [0:0] v_21;
  function [0:0] mux_21(input [0:0] sel);
    case (sel) 0: mux_21 = 1'h0; 1: mux_21 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22;
  wire [0:0] v_23;
  wire [0:0] v_24;
  wire [0:0] vin0_consume_en_25;
  wire [0:0] vout_canPeek_25;
  wire [7:0] vout_peek_25;
  wire [0:0] v_26;
  function [0:0] mux_26(input [0:0] sel);
    case (sel) 0: mux_26 = 1'h0; 1: mux_26 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_27;
  wire [0:0] v_28;
  wire [0:0] v_29;
  function [0:0] mux_29(input [0:0] sel);
    case (sel) 0: mux_29 = 1'h0; 1: mux_29 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_30;
  wire [0:0] vin0_consume_en_31;
  wire [0:0] vout_canPeek_31;
  wire [7:0] vout_peek_31;
  wire [0:0] v_32;
  function [0:0] mux_32(input [0:0] sel);
    case (sel) 0: mux_32 = 1'h0; 1: mux_32 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_33;
  wire [0:0] v_34;
  wire [0:0] v_35;
  function [0:0] mux_35(input [0:0] sel);
    case (sel) 0: mux_35 = 1'h0; 1: mux_35 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_36;
  wire [0:0] v_37;
  wire [0:0] v_38;
  wire [0:0] vin0_consume_en_39;
  wire [0:0] vout_canPeek_39;
  wire [7:0] vout_peek_39;
  wire [0:0] v_40;
  function [0:0] mux_40(input [0:0] sel);
    case (sel) 0: mux_40 = 1'h0; 1: mux_40 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_41;
  wire [0:0] v_42;
  wire [0:0] v_43;
  function [0:0] mux_43(input [0:0] sel);
    case (sel) 0: mux_43 = 1'h0; 1: mux_43 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_44;
  wire [0:0] vin0_consume_en_45;
  wire [0:0] vout_canPeek_45;
  wire [7:0] vout_peek_45;
  wire [0:0] v_46;
  function [0:0] mux_46(input [0:0] sel);
    case (sel) 0: mux_46 = 1'h0; 1: mux_46 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_47;
  wire [0:0] v_48;
  wire [0:0] v_49;
  function [0:0] mux_49(input [0:0] sel);
    case (sel) 0: mux_49 = 1'h0; 1: mux_49 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_50;
  wire [0:0] v_51;
  wire [0:0] v_52;
  wire [0:0] vin0_consume_en_53;
  wire [0:0] vout_canPeek_53;
  wire [7:0] vout_peek_53;
  wire [0:0] v_54;
  function [0:0] mux_54(input [0:0] sel);
    case (sel) 0: mux_54 = 1'h0; 1: mux_54 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_55;
  wire [0:0] v_56;
  wire [0:0] v_57;
  function [0:0] mux_57(input [0:0] sel);
    case (sel) 0: mux_57 = 1'h0; 1: mux_57 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_58;
  wire [0:0] vin0_consume_en_59;
  wire [0:0] vout_canPeek_59;
  wire [7:0] vout_peek_59;
  wire [0:0] v_60;
  function [0:0] mux_60(input [0:0] sel);
    case (sel) 0: mux_60 = 1'h0; 1: mux_60 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_61;
  wire [0:0] v_62;
  wire [0:0] v_63;
  function [0:0] mux_63(input [0:0] sel);
    case (sel) 0: mux_63 = 1'h0; 1: mux_63 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_64;
  wire [0:0] v_65;
  wire [0:0] v_66;
  wire [0:0] vin0_consume_en_67;
  wire [0:0] vout_canPeek_67;
  wire [7:0] vout_peek_67;
  wire [0:0] v_68;
  function [0:0] mux_68(input [0:0] sel);
    case (sel) 0: mux_68 = 1'h0; 1: mux_68 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_69;
  wire [0:0] v_71;
  function [0:0] mux_71(input [0:0] sel);
    case (sel) 0: mux_71 = 1'h0; 1: mux_71 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_72;
  reg [0:0] v_74 = 1'h0;
  wire [0:0] v_75;
  wire [0:0] v_76;
  wire [0:0] act_77;
  wire [0:0] v_78;
  wire [0:0] v_79;
  wire [0:0] v_80;
  reg [0:0] v_81 = 1'h0;
  wire [0:0] v_82;
  wire [0:0] v_83;
  wire [0:0] act_84;
  wire [0:0] v_85;
  wire [0:0] v_86;
  wire [0:0] v_87;
  reg [0:0] v_88 = 1'h0;
  wire [0:0] v_89;
  wire [0:0] v_90;
  wire [0:0] act_91;
  wire [0:0] v_92;
  wire [0:0] v_93;
  wire [0:0] v_94;
  wire [0:0] v_95;
  wire [0:0] v_96;
  wire [0:0] v_97;
  function [0:0] mux_97(input [0:0] sel);
    case (sel) 0: mux_97 = 1'h0; 1: mux_97 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_98;
  wire [0:0] v_99;
  function [0:0] mux_99(input [0:0] sel);
    case (sel) 0: mux_99 = 1'h0; 1: mux_99 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_100;
  wire [0:0] v_101;
  wire [0:0] v_102;
  wire [0:0] v_103;
  function [0:0] mux_103(input [0:0] sel);
    case (sel) 0: mux_103 = 1'h0; 1: mux_103 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_104;
  function [0:0] mux_104(input [0:0] sel);
    case (sel) 0: mux_104 = 1'h0; 1: mux_104 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_105 = 1'h0;
  wire [0:0] v_106;
  wire [0:0] v_107;
  wire [0:0] act_108;
  wire [0:0] v_109;
  wire [0:0] v_110;
  wire [0:0] v_111;
  wire [0:0] v_112;
  wire [0:0] v_113;
  wire [0:0] v_114;
  function [0:0] mux_114(input [0:0] sel);
    case (sel) 0: mux_114 = 1'h0; 1: mux_114 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_115;
  function [0:0] mux_115(input [0:0] sel);
    case (sel) 0: mux_115 = 1'h0; 1: mux_115 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_116;
  wire [0:0] v_117;
  wire [0:0] v_118;
  wire [0:0] v_119;
  function [0:0] mux_119(input [0:0] sel);
    case (sel) 0: mux_119 = 1'h0; 1: mux_119 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_120;
  function [0:0] mux_120(input [0:0] sel);
    case (sel) 0: mux_120 = 1'h0; 1: mux_120 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_121;
  wire [0:0] v_122;
  wire [0:0] v_123;
  wire [0:0] v_124;
  wire [0:0] v_125;
  wire [0:0] v_126;
  function [0:0] mux_126(input [0:0] sel);
    case (sel) 0: mux_126 = 1'h0; 1: mux_126 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_127;
  wire [0:0] v_128;
  function [0:0] mux_128(input [0:0] sel);
    case (sel) 0: mux_128 = 1'h0; 1: mux_128 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_129;
  wire [0:0] v_130;
  wire [0:0] v_131;
  wire [0:0] v_132;
  function [0:0] mux_132(input [0:0] sel);
    case (sel) 0: mux_132 = 1'h0; 1: mux_132 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_133;
  function [0:0] mux_133(input [0:0] sel);
    case (sel) 0: mux_133 = 1'h0; 1: mux_133 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_134 = 1'h0;
  wire [0:0] v_135;
  wire [0:0] v_136;
  wire [0:0] act_137;
  wire [0:0] v_138;
  wire [0:0] v_139;
  wire [0:0] v_140;
  reg [0:0] v_141 = 1'h0;
  wire [0:0] v_142;
  wire [0:0] v_143;
  wire [0:0] act_144;
  wire [0:0] v_145;
  wire [0:0] v_146;
  wire [0:0] v_147;
  wire [0:0] v_148;
  wire [0:0] v_149;
  wire [0:0] v_150;
  function [0:0] mux_150(input [0:0] sel);
    case (sel) 0: mux_150 = 1'h0; 1: mux_150 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_151;
  wire [0:0] v_152;
  function [0:0] mux_152(input [0:0] sel);
    case (sel) 0: mux_152 = 1'h0; 1: mux_152 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_153;
  wire [0:0] v_154;
  wire [0:0] v_155;
  wire [0:0] v_156;
  function [0:0] mux_156(input [0:0] sel);
    case (sel) 0: mux_156 = 1'h0; 1: mux_156 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_157;
  function [0:0] mux_157(input [0:0] sel);
    case (sel) 0: mux_157 = 1'h0; 1: mux_157 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_158 = 1'h0;
  wire [0:0] v_159;
  wire [0:0] v_160;
  wire [0:0] act_161;
  wire [0:0] v_162;
  wire [0:0] v_163;
  wire [0:0] v_164;
  reg [0:0] v_165 = 1'h0;
  wire [0:0] v_166;
  wire [0:0] v_167;
  wire [0:0] act_168;
  wire [0:0] v_169;
  wire [0:0] v_170;
  wire [0:0] v_171;
  wire [0:0] v_172;
  wire [0:0] v_173;
  wire [0:0] v_174;
  function [0:0] mux_174(input [0:0] sel);
    case (sel) 0: mux_174 = 1'h0; 1: mux_174 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_175;
  wire [0:0] v_176;
  function [0:0] mux_176(input [0:0] sel);
    case (sel) 0: mux_176 = 1'h0; 1: mux_176 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_177;
  wire [0:0] v_178;
  wire [0:0] v_179;
  wire [0:0] v_180;
  function [0:0] mux_180(input [0:0] sel);
    case (sel) 0: mux_180 = 1'h0; 1: mux_180 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_181;
  function [0:0] mux_181(input [0:0] sel);
    case (sel) 0: mux_181 = 1'h0; 1: mux_181 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_182 = 1'h0;
  wire [0:0] v_183;
  wire [0:0] v_184;
  wire [0:0] act_185;
  wire [0:0] v_186;
  wire [0:0] v_187;
  wire [0:0] v_188;
  wire [0:0] v_189;
  wire [0:0] v_190;
  wire [0:0] v_191;
  function [0:0] mux_191(input [0:0] sel);
    case (sel) 0: mux_191 = 1'h0; 1: mux_191 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_192;
  function [0:0] mux_192(input [0:0] sel);
    case (sel) 0: mux_192 = 1'h0; 1: mux_192 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_193;
  wire [0:0] v_194;
  wire [0:0] v_195;
  wire [0:0] v_196;
  function [0:0] mux_196(input [0:0] sel);
    case (sel) 0: mux_196 = 1'h0; 1: mux_196 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_197;
  function [0:0] mux_197(input [0:0] sel);
    case (sel) 0: mux_197 = 1'h0; 1: mux_197 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_198;
  wire [0:0] v_199;
  wire [0:0] v_200;
  wire [0:0] v_201;
  wire [0:0] v_202;
  wire [0:0] v_203;
  function [0:0] mux_203(input [0:0] sel);
    case (sel) 0: mux_203 = 1'h0; 1: mux_203 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_204;
  function [0:0] mux_204(input [0:0] sel);
    case (sel) 0: mux_204 = 1'h0; 1: mux_204 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_205;
  wire [0:0] v_206;
  wire [0:0] v_207;
  wire [0:0] v_208;
  function [0:0] mux_208(input [0:0] sel);
    case (sel) 0: mux_208 = 1'h0; 1: mux_208 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_209;
  function [0:0] mux_209(input [0:0] sel);
    case (sel) 0: mux_209 = 1'h0; 1: mux_209 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_210;
  wire [0:0] v_211;
  wire [0:0] v_212;
  wire [0:0] v_213;
  wire [0:0] v_214;
  wire [0:0] v_215;
  function [0:0] mux_215(input [0:0] sel);
    case (sel) 0: mux_215 = 1'h0; 1: mux_215 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_216;
  function [0:0] mux_216(input [0:0] sel);
    case (sel) 0: mux_216 = 1'h0; 1: mux_216 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_217;
  wire [0:0] v_218;
  wire [0:0] v_219;
  wire [0:0] v_220;
  function [0:0] mux_220(input [0:0] sel);
    case (sel) 0: mux_220 = 1'h0; 1: mux_220 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_221;
  function [0:0] mux_221(input [0:0] sel);
    case (sel) 0: mux_221 = 1'h0; 1: mux_221 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_222;
  wire [0:0] v_223;
  wire [0:0] v_224;
  wire [0:0] v_225;
  wire [0:0] v_226;
  wire [0:0] v_227;
  function [0:0] mux_227(input [0:0] sel);
    case (sel) 0: mux_227 = 1'h0; 1: mux_227 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_228;
  wire [0:0] v_229;
  wire [0:0] v_230;
  function [0:0] mux_230(input [0:0] sel);
    case (sel) 0: mux_230 = 1'h0; 1: mux_230 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_231;
  wire [0:0] v_232;
  wire [0:0] v_233;
  wire [0:0] v_234;
  function [0:0] mux_234(input [0:0] sel);
    case (sel) 0: mux_234 = 1'h0; 1: mux_234 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_235;
  function [0:0] mux_235(input [0:0] sel);
    case (sel) 0: mux_235 = 1'h0; 1: mux_235 = 1'h0;
    endcase
  endfunction
  reg [7:0] v_237 = 8'h0;
  wire [7:0] v_238;
  wire [7:0] v_239;
  function [7:0] mux_239(input [0:0] sel);
    case (sel) 0: mux_239 = 8'h0; 1: mux_239 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_240;
  wire [7:0] v_241;
  wire [7:0] v_242;
  function [7:0] mux_242(input [0:0] sel);
    case (sel) 0: mux_242 = 8'h0; 1: mux_242 = v_243;
    endcase
  endfunction
  reg [7:0] v_243 = 8'h0;
  wire [7:0] v_244;
  wire [7:0] v_245;
  function [7:0] mux_245(input [0:0] sel);
    case (sel) 0: mux_245 = 8'h0; 1: mux_245 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_246;
  wire [7:0] v_247;
  wire [7:0] v_248;
  function [7:0] mux_248(input [0:0] sel);
    case (sel) 0: mux_248 = 8'h0; 1: mux_248 = v_249;
    endcase
  endfunction
  reg [7:0] v_249 = 8'h0;
  wire [7:0] v_250;
  wire [7:0] v_251;
  function [7:0] mux_251(input [0:0] sel);
    case (sel) 0: mux_251 = 8'h0; 1: mux_251 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_252;
  wire [7:0] v_253;
  wire [7:0] v_254;
  function [7:0] mux_254(input [0:0] sel);
    case (sel) 0: mux_254 = 8'h0; 1: mux_254 = v_255;
    endcase
  endfunction
  reg [7:0] v_255 = 8'h0;
  wire [7:0] v_256;
  wire [7:0] v_257;
  function [7:0] mux_257(input [0:0] sel);
    case (sel) 0: mux_257 = 8'h0; 1: mux_257 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_258;
  wire [7:0] v_259;
  wire [7:0] v_260;
  function [7:0] mux_260(input [0:0] sel);
    case (sel) 0: mux_260 = 8'h0; 1: mux_260 = vout_peek_25;
    endcase
  endfunction
  wire [7:0] v_261;
  function [7:0] mux_261(input [0:0] sel);
    case (sel) 0: mux_261 = 8'h0; 1: mux_261 = vout_peek_17;
    endcase
  endfunction
  wire [7:0] v_262;
  function [7:0] mux_262(input [0:0] sel);
    case (sel) 0: mux_262 = 8'h0; 1: mux_262 = v_263;
    endcase
  endfunction
  reg [7:0] v_263 = 8'h0;
  wire [7:0] v_264;
  wire [7:0] v_265;
  function [7:0] mux_265(input [0:0] sel);
    case (sel) 0: mux_265 = 8'h0; 1: mux_265 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_266;
  wire [7:0] v_267;
  wire [7:0] v_268;
  function [7:0] mux_268(input [0:0] sel);
    case (sel) 0: mux_268 = 8'h0; 1: mux_268 = vout_peek_11;
    endcase
  endfunction
  wire [7:0] v_269;
  function [7:0] mux_269(input [0:0] sel);
    case (sel) 0: mux_269 = 8'h0; 1: mux_269 = vout_peek_3;
    endcase
  endfunction
  wire [7:0] v_270;
  function [7:0] mux_270(input [0:0] sel);
    case (sel) 0: mux_270 = 8'h0; 1: mux_270 = v_271;
    endcase
  endfunction
  reg [7:0] v_271 = 8'h0;
  wire [7:0] v_272;
  wire [7:0] v_273;
  function [7:0] mux_273(input [0:0] sel);
    case (sel) 0: mux_273 = 8'h0; 1: mux_273 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_274;
  wire [7:0] v_275;
  wire [7:0] v_276;
  function [7:0] mux_276(input [0:0] sel);
    case (sel) 0: mux_276 = 8'h0; 1: mux_276 = vout_peek_67;
    endcase
  endfunction
  wire [7:0] v_277;
  function [7:0] mux_277(input [0:0] sel);
    case (sel) 0: mux_277 = 8'h0; 1: mux_277 = vout_peek_59;
    endcase
  endfunction
  wire [7:0] v_278;
  function [7:0] mux_278(input [0:0] sel);
    case (sel) 0: mux_278 = 8'h0; 1: mux_278 = v_279;
    endcase
  endfunction
  reg [7:0] v_279 = 8'h0;
  wire [7:0] v_280;
  wire [7:0] v_281;
  function [7:0] mux_281(input [0:0] sel);
    case (sel) 0: mux_281 = 8'h0; 1: mux_281 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_282;
  wire [7:0] v_283;
  wire [7:0] v_284;
  function [7:0] mux_284(input [0:0] sel);
    case (sel) 0: mux_284 = 8'h0; 1: mux_284 = v_285;
    endcase
  endfunction
  reg [7:0] v_285 = 8'h0;
  wire [7:0] v_286;
  wire [7:0] v_287;
  function [7:0] mux_287(input [0:0] sel);
    case (sel) 0: mux_287 = 8'h0; 1: mux_287 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_288;
  wire [7:0] v_289;
  wire [7:0] v_290;
  function [7:0] mux_290(input [0:0] sel);
    case (sel) 0: mux_290 = 8'h0; 1: mux_290 = vout_peek_53;
    endcase
  endfunction
  wire [7:0] v_291;
  function [7:0] mux_291(input [0:0] sel);
    case (sel) 0: mux_291 = 8'h0; 1: mux_291 = vout_peek_45;
    endcase
  endfunction
  wire [7:0] v_292;
  function [7:0] mux_292(input [0:0] sel);
    case (sel) 0: mux_292 = 8'h0; 1: mux_292 = v_293;
    endcase
  endfunction
  reg [7:0] v_293 = 8'h0;
  wire [7:0] v_294;
  wire [7:0] v_295;
  function [7:0] mux_295(input [0:0] sel);
    case (sel) 0: mux_295 = 8'h0; 1: mux_295 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_296;
  wire [7:0] v_297;
  wire [7:0] v_298;
  function [7:0] mux_298(input [0:0] sel);
    case (sel) 0: mux_298 = 8'h0; 1: mux_298 = vout_peek_39;
    endcase
  endfunction
  wire [7:0] v_299;
  function [7:0] mux_299(input [0:0] sel);
    case (sel) 0: mux_299 = 8'h0; 1: mux_299 = vout_peek_31;
    endcase
  endfunction
  wire [0:0] v_300;
  wire [7:0] v_301;
  // Instances
  //////////////////////////////////////////////////////////////////////////////
  assign v_0 = v_1 | v_4;
  assign v_1 = mux_1(v_2);
  assign v_2 = vout_canPeek_3 & 1'h1;
  pebbles_core
    pebbles_core_3
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_0),
       .in0_consume_en(vin0_consume_en_3),
       .out_canPeek(vout_canPeek_3),
       .out_peek(vout_peek_3));
  assign v_4 = mux_4(v_5);
  assign v_5 = ~v_2;
  assign v_6 = v_7 | v_12;
  assign v_7 = mux_7(v_8);
  assign v_8 = v_9 & 1'h1;
  assign v_9 = v_10 & vout_canPeek_11;
  assign v_10 = ~vout_canPeek_3;
  pebbles_core
    pebbles_core_11
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6),
       .in0_consume_en(vin0_consume_en_11),
       .out_canPeek(vout_canPeek_11),
       .out_peek(vout_peek_11));
  assign v_12 = mux_12(v_13);
  assign v_13 = ~v_8;
  assign v_14 = v_15 | v_18;
  assign v_15 = mux_15(v_16);
  assign v_16 = vout_canPeek_17 & 1'h1;
  pebbles_core
    pebbles_core_17
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14),
       .in0_consume_en(vin0_consume_en_17),
       .out_canPeek(vout_canPeek_17),
       .out_peek(vout_peek_17));
  assign v_18 = mux_18(v_19);
  assign v_19 = ~v_16;
  assign v_20 = v_21 | v_26;
  assign v_21 = mux_21(v_22);
  assign v_22 = v_23 & 1'h1;
  assign v_23 = v_24 & vout_canPeek_25;
  assign v_24 = ~vout_canPeek_17;
  pebbles_core
    pebbles_core_25
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20),
       .in0_consume_en(vin0_consume_en_25),
       .out_canPeek(vout_canPeek_25),
       .out_peek(vout_peek_25));
  assign v_26 = mux_26(v_27);
  assign v_27 = ~v_22;
  assign v_28 = v_29 | v_32;
  assign v_29 = mux_29(v_30);
  assign v_30 = vout_canPeek_31 & 1'h1;
  pebbles_core
    pebbles_core_31
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_28),
       .in0_consume_en(vin0_consume_en_31),
       .out_canPeek(vout_canPeek_31),
       .out_peek(vout_peek_31));
  assign v_32 = mux_32(v_33);
  assign v_33 = ~v_30;
  assign v_34 = v_35 | v_40;
  assign v_35 = mux_35(v_36);
  assign v_36 = v_37 & 1'h1;
  assign v_37 = v_38 & vout_canPeek_39;
  assign v_38 = ~vout_canPeek_31;
  pebbles_core
    pebbles_core_39
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_34),
       .in0_consume_en(vin0_consume_en_39),
       .out_canPeek(vout_canPeek_39),
       .out_peek(vout_peek_39));
  assign v_40 = mux_40(v_41);
  assign v_41 = ~v_36;
  assign v_42 = v_43 | v_46;
  assign v_43 = mux_43(v_44);
  assign v_44 = vout_canPeek_45 & 1'h1;
  pebbles_core
    pebbles_core_45
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_42),
       .in0_consume_en(vin0_consume_en_45),
       .out_canPeek(vout_canPeek_45),
       .out_peek(vout_peek_45));
  assign v_46 = mux_46(v_47);
  assign v_47 = ~v_44;
  assign v_48 = v_49 | v_54;
  assign v_49 = mux_49(v_50);
  assign v_50 = v_51 & 1'h1;
  assign v_51 = v_52 & vout_canPeek_53;
  assign v_52 = ~vout_canPeek_45;
  pebbles_core
    pebbles_core_53
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_48),
       .in0_consume_en(vin0_consume_en_53),
       .out_canPeek(vout_canPeek_53),
       .out_peek(vout_peek_53));
  assign v_54 = mux_54(v_55);
  assign v_55 = ~v_50;
  assign v_56 = v_57 | v_60;
  assign v_57 = mux_57(v_58);
  assign v_58 = vout_canPeek_59 & 1'h1;
  pebbles_core
    pebbles_core_59
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_56),
       .in0_consume_en(vin0_consume_en_59),
       .out_canPeek(vout_canPeek_59),
       .out_peek(vout_peek_59));
  assign v_60 = mux_60(v_61);
  assign v_61 = ~v_58;
  assign v_62 = v_63 | v_68;
  assign v_63 = mux_63(v_64);
  assign v_64 = v_65 & 1'h1;
  assign v_65 = v_66 & vout_canPeek_67;
  assign v_66 = ~vout_canPeek_59;
  pebbles_core
    pebbles_core_67
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_62),
       .in0_consume_en(vin0_consume_en_67),
       .out_canPeek(vout_canPeek_67),
       .out_peek(vout_peek_67));
  assign v_68 = mux_68(v_69);
  assign v_69 = ~v_64;
  assign in0_consume_en = v_71;
  assign v_71 = mux_71(v_72);
  assign v_72 = ~1'h0;
  assign out_canPeek = v_74;
  assign v_75 = v_76 | v_222;
  assign v_76 = act_77 & 1'h1;
  assign act_77 = v_78 | v_127;
  assign v_78 = v_79 & 1'h1;
  assign v_79 = v_80 & v_134;
  assign v_80 = ~v_81;
  assign v_82 = v_83 | v_121;
  assign v_83 = act_84 & 1'h1;
  assign act_84 = v_85 | v_98;
  assign v_85 = v_86 & 1'h1;
  assign v_86 = v_87 & v_105;
  assign v_87 = ~v_88;
  assign v_89 = v_90 | v_92;
  assign v_90 = act_91 & 1'h1;
  assign act_91 = v_36 | v_30;
  assign v_92 = v_93 & 1'h1;
  assign v_93 = v_94 & v_95;
  assign v_94 = ~act_91;
  assign v_95 = v_96 | v_101;
  assign v_96 = v_97 | v_99;
  assign v_97 = mux_97(v_98);
  assign v_98 = v_88 & 1'h1;
  assign v_99 = mux_99(v_100);
  assign v_100 = ~v_98;
  assign v_101 = ~v_88;
  assign v_102 = v_103 | v_104;
  assign v_103 = mux_103(v_90);
  assign v_104 = mux_104(v_92);
  assign v_106 = v_107 | v_109;
  assign v_107 = act_108 & 1'h1;
  assign act_108 = v_50 | v_44;
  assign v_109 = v_110 & 1'h1;
  assign v_110 = v_111 & v_112;
  assign v_111 = ~act_108;
  assign v_112 = v_113 | v_117;
  assign v_113 = v_114 | v_115;
  assign v_114 = mux_114(v_85);
  assign v_115 = mux_115(v_116);
  assign v_116 = ~v_85;
  assign v_117 = ~v_105;
  assign v_118 = v_119 | v_120;
  assign v_119 = mux_119(v_107);
  assign v_120 = mux_120(v_109);
  assign v_121 = v_122 & 1'h1;
  assign v_122 = v_123 & v_124;
  assign v_123 = ~act_84;
  assign v_124 = v_125 | v_130;
  assign v_125 = v_126 | v_128;
  assign v_126 = mux_126(v_127);
  assign v_127 = v_81 & 1'h1;
  assign v_128 = mux_128(v_129);
  assign v_129 = ~v_127;
  assign v_130 = ~v_81;
  assign v_131 = v_132 | v_133;
  assign v_132 = mux_132(v_83);
  assign v_133 = mux_133(v_121);
  assign v_135 = v_136 | v_210;
  assign v_136 = act_137 & 1'h1;
  assign act_137 = v_138 | v_151;
  assign v_138 = v_139 & 1'h1;
  assign v_139 = v_140 & v_158;
  assign v_140 = ~v_141;
  assign v_142 = v_143 | v_145;
  assign v_143 = act_144 & 1'h1;
  assign act_144 = v_64 | v_58;
  assign v_145 = v_146 & 1'h1;
  assign v_146 = v_147 & v_148;
  assign v_147 = ~act_144;
  assign v_148 = v_149 | v_154;
  assign v_149 = v_150 | v_152;
  assign v_150 = mux_150(v_151);
  assign v_151 = v_141 & 1'h1;
  assign v_152 = mux_152(v_153);
  assign v_153 = ~v_151;
  assign v_154 = ~v_141;
  assign v_155 = v_156 | v_157;
  assign v_156 = mux_156(v_143);
  assign v_157 = mux_157(v_145);
  assign v_159 = v_160 | v_198;
  assign v_160 = act_161 & 1'h1;
  assign act_161 = v_162 | v_175;
  assign v_162 = v_163 & 1'h1;
  assign v_163 = v_164 & v_182;
  assign v_164 = ~v_165;
  assign v_166 = v_167 | v_169;
  assign v_167 = act_168 & 1'h1;
  assign act_168 = v_8 | v_2;
  assign v_169 = v_170 & 1'h1;
  assign v_170 = v_171 & v_172;
  assign v_171 = ~act_168;
  assign v_172 = v_173 | v_178;
  assign v_173 = v_174 | v_176;
  assign v_174 = mux_174(v_175);
  assign v_175 = v_165 & 1'h1;
  assign v_176 = mux_176(v_177);
  assign v_177 = ~v_175;
  assign v_178 = ~v_165;
  assign v_179 = v_180 | v_181;
  assign v_180 = mux_180(v_167);
  assign v_181 = mux_181(v_169);
  assign v_183 = v_184 | v_186;
  assign v_184 = act_185 & 1'h1;
  assign act_185 = v_22 | v_16;
  assign v_186 = v_187 & 1'h1;
  assign v_187 = v_188 & v_189;
  assign v_188 = ~act_185;
  assign v_189 = v_190 | v_194;
  assign v_190 = v_191 | v_192;
  assign v_191 = mux_191(v_162);
  assign v_192 = mux_192(v_193);
  assign v_193 = ~v_162;
  assign v_194 = ~v_182;
  assign v_195 = v_196 | v_197;
  assign v_196 = mux_196(v_184);
  assign v_197 = mux_197(v_186);
  assign v_198 = v_199 & 1'h1;
  assign v_199 = v_200 & v_201;
  assign v_200 = ~act_161;
  assign v_201 = v_202 | v_206;
  assign v_202 = v_203 | v_204;
  assign v_203 = mux_203(v_138);
  assign v_204 = mux_204(v_205);
  assign v_205 = ~v_138;
  assign v_206 = ~v_158;
  assign v_207 = v_208 | v_209;
  assign v_208 = mux_208(v_160);
  assign v_209 = mux_209(v_198);
  assign v_210 = v_211 & 1'h1;
  assign v_211 = v_212 & v_213;
  assign v_212 = ~act_137;
  assign v_213 = v_214 | v_218;
  assign v_214 = v_215 | v_216;
  assign v_215 = mux_215(v_78);
  assign v_216 = mux_216(v_217);
  assign v_217 = ~v_78;
  assign v_218 = ~v_134;
  assign v_219 = v_220 | v_221;
  assign v_220 = mux_220(v_136);
  assign v_221 = mux_221(v_210);
  assign v_222 = v_223 & 1'h1;
  assign v_223 = v_224 & v_225;
  assign v_224 = ~act_77;
  assign v_225 = v_226 | v_232;
  assign v_226 = v_227 | v_230;
  assign v_227 = mux_227(v_228);
  assign v_228 = v_229 & 1'h1;
  assign v_229 = out_consume_en;
  assign v_230 = mux_230(v_231);
  assign v_231 = ~v_228;
  assign v_232 = ~v_74;
  assign v_233 = v_234 | v_235;
  assign v_234 = mux_234(v_76);
  assign v_235 = mux_235(v_222);
  assign out_peek = v_237;
  assign v_238 = v_239 | v_241;
  assign v_239 = mux_239(v_240);
  assign v_240 = ~act_77;
  assign v_241 = v_242 | v_278;
  assign v_242 = mux_242(v_78);
  assign v_244 = v_245 | v_247;
  assign v_245 = mux_245(v_246);
  assign v_246 = ~act_137;
  assign v_247 = v_248 | v_270;
  assign v_248 = mux_248(v_138);
  assign v_250 = v_251 | v_253;
  assign v_251 = mux_251(v_252);
  assign v_252 = ~act_161;
  assign v_253 = v_254 | v_262;
  assign v_254 = mux_254(v_162);
  assign v_256 = v_257 | v_259;
  assign v_257 = mux_257(v_258);
  assign v_258 = ~act_185;
  assign v_259 = v_260 | v_261;
  assign v_260 = mux_260(v_22);
  assign v_261 = mux_261(v_16);
  assign v_262 = mux_262(v_175);
  assign v_264 = v_265 | v_267;
  assign v_265 = mux_265(v_266);
  assign v_266 = ~act_168;
  assign v_267 = v_268 | v_269;
  assign v_268 = mux_268(v_8);
  assign v_269 = mux_269(v_2);
  assign v_270 = mux_270(v_151);
  assign v_272 = v_273 | v_275;
  assign v_273 = mux_273(v_274);
  assign v_274 = ~act_144;
  assign v_275 = v_276 | v_277;
  assign v_276 = mux_276(v_64);
  assign v_277 = mux_277(v_58);
  assign v_278 = mux_278(v_127);
  assign v_280 = v_281 | v_283;
  assign v_281 = mux_281(v_282);
  assign v_282 = ~act_84;
  assign v_283 = v_284 | v_292;
  assign v_284 = mux_284(v_85);
  assign v_286 = v_287 | v_289;
  assign v_287 = mux_287(v_288);
  assign v_288 = ~act_108;
  assign v_289 = v_290 | v_291;
  assign v_290 = mux_290(v_50);
  assign v_291 = mux_291(v_44);
  assign v_292 = mux_292(v_98);
  assign v_294 = v_295 | v_297;
  assign v_295 = mux_295(v_296);
  assign v_296 = ~act_91;
  assign v_297 = v_298 | v_299;
  assign v_298 = mux_298(v_36);
  assign v_299 = mux_299(v_30);
  assign v_300 = in0_canPeek;
  assign v_301 = in0_peek;
  // Always block
  //////////////////////////////////////////////////////////////////////////////
  always @(posedge clock) begin
    if (reset) begin
      v_74 <= 1'h0;
      v_81 <= 1'h0;
      v_88 <= 1'h0;
      v_105 <= 1'h0;
      v_134 <= 1'h0;
      v_141 <= 1'h0;
      v_158 <= 1'h0;
      v_165 <= 1'h0;
      v_182 <= 1'h0;
      v_237 <= 8'h0;
      v_243 <= 8'h0;
      v_249 <= 8'h0;
      v_255 <= 8'h0;
      v_263 <= 8'h0;
      v_271 <= 8'h0;
      v_279 <= 8'h0;
      v_285 <= 8'h0;
      v_293 <= 8'h0;
    end else begin
      if (v_75 == 1) v_74 <= v_233;
      if (v_82 == 1) v_81 <= v_131;
      if (v_89 == 1) v_88 <= v_102;
      if (v_106 == 1) v_105 <= v_118;
      if (v_135 == 1) v_134 <= v_219;
      if (v_142 == 1) v_141 <= v_155;
      if (v_159 == 1) v_158 <= v_207;
      if (v_166 == 1) v_165 <= v_179;
      if (v_183 == 1) v_182 <= v_195;
      if (v_76 == 1) v_237 <= v_238;
      if (v_136 == 1) v_243 <= v_244;
      if (v_160 == 1) v_249 <= v_250;
      if (v_184 == 1) v_255 <= v_256;
      if (v_167 == 1) v_263 <= v_264;
      if (v_143 == 1) v_271 <= v_272;
      if (v_83 == 1) v_279 <= v_280;
      if (v_107 == 1) v_285 <= v_286;
      if (v_90 == 1) v_293 <= v_294;
    end
  end
endmodule