module Pebbles
  (input wire clock,
   input wire reset,
   input wire [0:0] out_consume_en,
   input wire [0:0] in0_canPeek,
   input wire [7:0] in0_peek,
   output wire [0:0] in0_consume_en,
   output wire [0:0] out_canPeek,
   output wire [7:0] out_peek);
  // Declarations
  //////////////////////////////////////////////////////////////////////////////
  wire [0:0] v_0;
  wire [0:0] v_1;
  function [0:0] mux_1(input [0:0] sel);
    case (sel) 0: mux_1 = 1'h0; 1: mux_1 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2;
  wire [0:0] vin0_consume_en_3;
  wire [0:0] vout_canPeek_3;
  wire [7:0] vout_peek_3;
  wire [0:0] v_4;
  wire [0:0] v_5;
  wire [0:0] v_6;
  reg [0:0] v_7 = 1'h0;
  wire [0:0] v_8;
  wire [0:0] v_9;
  wire [0:0] act_10;
  wire [0:0] v_11;
  wire [0:0] v_12;
  wire [0:0] v_13;
  wire [0:0] vin0_consume_en_14;
  wire [0:0] vout_canPeek_14;
  wire [7:0] vout_peek_14;
  wire [0:0] v_15;
  wire [0:0] v_16;
  function [0:0] mux_16(input [0:0] sel);
    case (sel) 0: mux_16 = 1'h0; 1: mux_16 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17;
  function [0:0] mux_17(input [0:0] sel);
    case (sel) 0: mux_17 = 1'h0; 1: mux_17 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18;
  wire [0:0] v_19;
  wire [0:0] v_20;
  wire [0:0] v_21;
  wire [0:0] v_22;
  wire [0:0] v_23;
  wire [0:0] v_24;
  function [0:0] mux_24(input [0:0] sel);
    case (sel) 0: mux_24 = 1'h0; 1: mux_24 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_25;
  wire [0:0] v_26;
  wire [0:0] v_27;
  wire [0:0] v_28;
  reg [0:0] v_29 = 1'h0;
  wire [0:0] v_30;
  wire [0:0] v_31;
  wire [0:0] act_32;
  wire [0:0] v_33;
  wire [0:0] v_34;
  wire [0:0] v_35;
  reg [0:0] v_36 = 1'h0;
  wire [0:0] v_37;
  wire [0:0] v_38;
  wire [0:0] act_39;
  wire [0:0] v_40;
  wire [0:0] v_41;
  wire [0:0] v_42;
  wire [0:0] vin0_consume_en_43;
  wire [0:0] vout_canPeek_43;
  wire [7:0] vout_peek_43;
  wire [0:0] v_44;
  wire [0:0] v_45;
  function [0:0] mux_45(input [0:0] sel);
    case (sel) 0: mux_45 = 1'h0; 1: mux_45 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_46;
  wire [0:0] v_47;
  wire [0:0] v_48;
  wire [0:0] v_49;
  wire [0:0] v_50;
  function [0:0] mux_50(input [0:0] sel);
    case (sel) 0: mux_50 = 1'h0; 1: mux_50 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_51;
  wire [0:0] vin0_consume_en_52;
  wire [0:0] vout_canPeek_52;
  wire [7:0] vout_peek_52;
  wire [0:0] v_53;
  wire [0:0] v_54;
  function [0:0] mux_54(input [0:0] sel);
    case (sel) 0: mux_54 = 1'h0; 1: mux_54 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_55;
  function [0:0] mux_55(input [0:0] sel);
    case (sel) 0: mux_55 = 1'h0; 1: mux_55 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_56;
  wire [0:0] v_57;
  wire [0:0] v_58;
  wire [0:0] v_59;
  wire [0:0] v_60;
  wire [0:0] v_61;
  wire [0:0] v_62;
  function [0:0] mux_62(input [0:0] sel);
    case (sel) 0: mux_62 = 1'h0; 1: mux_62 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_63;
  function [0:0] mux_63(input [0:0] sel);
    case (sel) 0: mux_63 = 1'h0; 1: mux_63 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_64;
  wire [0:0] v_65;
  wire [0:0] v_66;
  wire [0:0] v_67;
  function [0:0] mux_67(input [0:0] sel);
    case (sel) 0: mux_67 = 1'h0; 1: mux_67 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_68;
  function [0:0] mux_68(input [0:0] sel);
    case (sel) 0: mux_68 = 1'h0; 1: mux_68 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_69;
  wire [0:0] v_70;
  wire [0:0] v_71;
  wire [0:0] v_72;
  wire [0:0] v_73;
  wire [0:0] v_74;
  function [0:0] mux_74(input [0:0] sel);
    case (sel) 0: mux_74 = 1'h0; 1: mux_74 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_75;
  wire [0:0] v_76;
  wire [0:0] v_77;
  wire [0:0] v_78;
  reg [0:0] v_79 = 1'h0;
  wire [0:0] v_80;
  wire [0:0] v_81;
  wire [0:0] act_82;
  wire [0:0] v_83;
  wire [0:0] v_84;
  wire [0:0] v_85;
  reg [0:0] v_86 = 1'h0;
  wire [0:0] v_87;
  wire [0:0] v_88;
  wire [0:0] act_89;
  wire [0:0] v_90;
  wire [0:0] v_91;
  wire [0:0] v_92;
  reg [0:0] v_93 = 1'h0;
  wire [0:0] v_94;
  wire [0:0] v_95;
  wire [0:0] act_96;
  wire [0:0] v_97;
  wire [0:0] v_98;
  wire [0:0] v_99;
  wire [0:0] vin0_consume_en_100;
  wire [0:0] vout_canPeek_100;
  wire [7:0] vout_peek_100;
  wire [0:0] v_101;
  wire [0:0] v_102;
  function [0:0] mux_102(input [0:0] sel);
    case (sel) 0: mux_102 = 1'h0; 1: mux_102 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_103;
  wire [0:0] v_104;
  wire [0:0] v_105;
  wire [0:0] v_106;
  wire [0:0] v_107;
  function [0:0] mux_107(input [0:0] sel);
    case (sel) 0: mux_107 = 1'h0; 1: mux_107 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_108;
  wire [0:0] vin0_consume_en_109;
  wire [0:0] vout_canPeek_109;
  wire [7:0] vout_peek_109;
  wire [0:0] v_110;
  wire [0:0] v_111;
  function [0:0] mux_111(input [0:0] sel);
    case (sel) 0: mux_111 = 1'h0; 1: mux_111 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_112;
  function [0:0] mux_112(input [0:0] sel);
    case (sel) 0: mux_112 = 1'h0; 1: mux_112 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_113;
  wire [0:0] v_114;
  wire [0:0] v_115;
  wire [0:0] v_116;
  wire [0:0] v_117;
  wire [0:0] v_118;
  wire [0:0] v_119;
  function [0:0] mux_119(input [0:0] sel);
    case (sel) 0: mux_119 = 1'h0; 1: mux_119 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_120;
  wire [0:0] v_121;
  wire [0:0] v_122;
  wire [0:0] v_123;
  wire [0:0] v_124;
  function [0:0] mux_124(input [0:0] sel);
    case (sel) 0: mux_124 = 1'h0; 1: mux_124 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_125;
  wire [0:0] v_126;
  wire [0:0] v_127;
  wire [0:0] v_128;
  function [0:0] mux_128(input [0:0] sel);
    case (sel) 0: mux_128 = 1'h0; 1: mux_128 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_129;
  function [0:0] mux_129(input [0:0] sel);
    case (sel) 0: mux_129 = 1'h0; 1: mux_129 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_130 = 1'h0;
  wire [0:0] v_131;
  wire [0:0] v_132;
  wire [0:0] act_133;
  wire [0:0] v_134;
  wire [0:0] v_135;
  wire [0:0] v_136;
  wire [0:0] vin0_consume_en_137;
  wire [0:0] vout_canPeek_137;
  wire [7:0] vout_peek_137;
  wire [0:0] v_138;
  wire [0:0] v_139;
  function [0:0] mux_139(input [0:0] sel);
    case (sel) 0: mux_139 = 1'h0; 1: mux_139 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_140;
  wire [0:0] v_141;
  wire [0:0] v_142;
  wire [0:0] v_143;
  wire [0:0] v_144;
  function [0:0] mux_144(input [0:0] sel);
    case (sel) 0: mux_144 = 1'h0; 1: mux_144 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_145;
  wire [0:0] vin0_consume_en_146;
  wire [0:0] vout_canPeek_146;
  wire [7:0] vout_peek_146;
  wire [0:0] v_147;
  wire [0:0] v_148;
  function [0:0] mux_148(input [0:0] sel);
    case (sel) 0: mux_148 = 1'h0; 1: mux_148 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_149;
  function [0:0] mux_149(input [0:0] sel);
    case (sel) 0: mux_149 = 1'h0; 1: mux_149 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_150;
  wire [0:0] v_151;
  wire [0:0] v_152;
  wire [0:0] v_153;
  wire [0:0] v_154;
  wire [0:0] v_155;
  wire [0:0] v_156;
  function [0:0] mux_156(input [0:0] sel);
    case (sel) 0: mux_156 = 1'h0; 1: mux_156 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_157;
  function [0:0] mux_157(input [0:0] sel);
    case (sel) 0: mux_157 = 1'h0; 1: mux_157 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_158;
  wire [0:0] v_159;
  wire [0:0] v_160;
  wire [0:0] v_161;
  function [0:0] mux_161(input [0:0] sel);
    case (sel) 0: mux_161 = 1'h0; 1: mux_161 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_162;
  function [0:0] mux_162(input [0:0] sel);
    case (sel) 0: mux_162 = 1'h0; 1: mux_162 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_163;
  wire [0:0] v_164;
  wire [0:0] v_165;
  wire [0:0] v_166;
  wire [0:0] v_167;
  wire [0:0] v_168;
  function [0:0] mux_168(input [0:0] sel);
    case (sel) 0: mux_168 = 1'h0; 1: mux_168 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_169;
  function [0:0] mux_169(input [0:0] sel);
    case (sel) 0: mux_169 = 1'h0; 1: mux_169 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_170;
  wire [0:0] v_171;
  wire [0:0] v_172;
  wire [0:0] v_173;
  function [0:0] mux_173(input [0:0] sel);
    case (sel) 0: mux_173 = 1'h0; 1: mux_173 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_174;
  function [0:0] mux_174(input [0:0] sel);
    case (sel) 0: mux_174 = 1'h0; 1: mux_174 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_175;
  wire [0:0] v_176;
  wire [0:0] v_177;
  wire [0:0] v_178;
  wire [0:0] v_179;
  wire [0:0] v_180;
  function [0:0] mux_180(input [0:0] sel);
    case (sel) 0: mux_180 = 1'h0; 1: mux_180 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_181;
  wire [0:0] v_182;
  wire [0:0] v_183;
  wire [0:0] v_184;
  reg [0:0] v_185 = 1'h0;
  wire [0:0] v_186;
  wire [0:0] v_187;
  wire [0:0] act_188;
  wire [0:0] v_189;
  wire [0:0] v_190;
  wire [0:0] v_191;
  reg [0:0] v_192 = 1'h0;
  wire [0:0] v_193;
  wire [0:0] v_194;
  wire [0:0] act_195;
  wire [0:0] v_196;
  wire [0:0] v_197;
  wire [0:0] v_198;
  reg [0:0] v_199 = 1'h0;
  wire [0:0] v_200;
  wire [0:0] v_201;
  wire [0:0] act_202;
  wire [0:0] v_203;
  wire [0:0] v_204;
  wire [0:0] v_205;
  reg [0:0] v_206 = 1'h0;
  wire [0:0] v_207;
  wire [0:0] v_208;
  wire [0:0] act_209;
  wire [0:0] v_210;
  wire [0:0] v_211;
  wire [0:0] v_212;
  wire [0:0] vin0_consume_en_213;
  wire [0:0] vout_canPeek_213;
  wire [7:0] vout_peek_213;
  wire [0:0] v_214;
  wire [0:0] v_215;
  function [0:0] mux_215(input [0:0] sel);
    case (sel) 0: mux_215 = 1'h0; 1: mux_215 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_216;
  wire [0:0] v_217;
  wire [0:0] v_218;
  wire [0:0] v_219;
  wire [0:0] v_220;
  function [0:0] mux_220(input [0:0] sel);
    case (sel) 0: mux_220 = 1'h0; 1: mux_220 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_221;
  wire [0:0] vin0_consume_en_222;
  wire [0:0] vout_canPeek_222;
  wire [7:0] vout_peek_222;
  wire [0:0] v_223;
  wire [0:0] v_224;
  function [0:0] mux_224(input [0:0] sel);
    case (sel) 0: mux_224 = 1'h0; 1: mux_224 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_225;
  function [0:0] mux_225(input [0:0] sel);
    case (sel) 0: mux_225 = 1'h0; 1: mux_225 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_226;
  wire [0:0] v_227;
  wire [0:0] v_228;
  wire [0:0] v_229;
  wire [0:0] v_230;
  wire [0:0] v_231;
  wire [0:0] v_232;
  function [0:0] mux_232(input [0:0] sel);
    case (sel) 0: mux_232 = 1'h0; 1: mux_232 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_233;
  wire [0:0] v_234;
  wire [0:0] v_235;
  wire [0:0] v_236;
  wire [0:0] v_237;
  function [0:0] mux_237(input [0:0] sel);
    case (sel) 0: mux_237 = 1'h0; 1: mux_237 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_238;
  wire [0:0] v_239;
  wire [0:0] v_240;
  wire [0:0] v_241;
  function [0:0] mux_241(input [0:0] sel);
    case (sel) 0: mux_241 = 1'h0; 1: mux_241 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_242;
  function [0:0] mux_242(input [0:0] sel);
    case (sel) 0: mux_242 = 1'h0; 1: mux_242 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_243 = 1'h0;
  wire [0:0] v_244;
  wire [0:0] v_245;
  wire [0:0] act_246;
  wire [0:0] v_247;
  wire [0:0] v_248;
  wire [0:0] v_249;
  wire [0:0] vin0_consume_en_250;
  wire [0:0] vout_canPeek_250;
  wire [7:0] vout_peek_250;
  wire [0:0] v_251;
  wire [0:0] v_252;
  function [0:0] mux_252(input [0:0] sel);
    case (sel) 0: mux_252 = 1'h0; 1: mux_252 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_253;
  wire [0:0] v_254;
  wire [0:0] v_255;
  wire [0:0] v_256;
  wire [0:0] v_257;
  function [0:0] mux_257(input [0:0] sel);
    case (sel) 0: mux_257 = 1'h0; 1: mux_257 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_258;
  wire [0:0] vin0_consume_en_259;
  wire [0:0] vout_canPeek_259;
  wire [7:0] vout_peek_259;
  wire [0:0] v_260;
  wire [0:0] v_261;
  function [0:0] mux_261(input [0:0] sel);
    case (sel) 0: mux_261 = 1'h0; 1: mux_261 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_262;
  function [0:0] mux_262(input [0:0] sel);
    case (sel) 0: mux_262 = 1'h0; 1: mux_262 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_263;
  wire [0:0] v_264;
  wire [0:0] v_265;
  wire [0:0] v_266;
  wire [0:0] v_267;
  wire [0:0] v_268;
  wire [0:0] v_269;
  function [0:0] mux_269(input [0:0] sel);
    case (sel) 0: mux_269 = 1'h0; 1: mux_269 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_270;
  function [0:0] mux_270(input [0:0] sel);
    case (sel) 0: mux_270 = 1'h0; 1: mux_270 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_271;
  wire [0:0] v_272;
  wire [0:0] v_273;
  wire [0:0] v_274;
  function [0:0] mux_274(input [0:0] sel);
    case (sel) 0: mux_274 = 1'h0; 1: mux_274 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_275;
  function [0:0] mux_275(input [0:0] sel);
    case (sel) 0: mux_275 = 1'h0; 1: mux_275 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_276;
  wire [0:0] v_277;
  wire [0:0] v_278;
  wire [0:0] v_279;
  wire [0:0] v_280;
  wire [0:0] v_281;
  function [0:0] mux_281(input [0:0] sel);
    case (sel) 0: mux_281 = 1'h0; 1: mux_281 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_282;
  wire [0:0] v_283;
  wire [0:0] v_284;
  wire [0:0] v_285;
  wire [0:0] v_286;
  function [0:0] mux_286(input [0:0] sel);
    case (sel) 0: mux_286 = 1'h0; 1: mux_286 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_287;
  wire [0:0] v_288;
  wire [0:0] v_289;
  wire [0:0] v_290;
  function [0:0] mux_290(input [0:0] sel);
    case (sel) 0: mux_290 = 1'h0; 1: mux_290 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_291;
  function [0:0] mux_291(input [0:0] sel);
    case (sel) 0: mux_291 = 1'h0; 1: mux_291 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_292 = 1'h0;
  wire [0:0] v_293;
  wire [0:0] v_294;
  wire [0:0] act_295;
  wire [0:0] v_296;
  wire [0:0] v_297;
  wire [0:0] v_298;
  reg [0:0] v_299 = 1'h0;
  wire [0:0] v_300;
  wire [0:0] v_301;
  wire [0:0] act_302;
  wire [0:0] v_303;
  wire [0:0] v_304;
  wire [0:0] v_305;
  wire [0:0] vin0_consume_en_306;
  wire [0:0] vout_canPeek_306;
  wire [7:0] vout_peek_306;
  wire [0:0] v_307;
  wire [0:0] v_308;
  function [0:0] mux_308(input [0:0] sel);
    case (sel) 0: mux_308 = 1'h0; 1: mux_308 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_309;
  wire [0:0] v_310;
  wire [0:0] v_311;
  wire [0:0] v_312;
  wire [0:0] v_313;
  function [0:0] mux_313(input [0:0] sel);
    case (sel) 0: mux_313 = 1'h0; 1: mux_313 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_314;
  wire [0:0] vin0_consume_en_315;
  wire [0:0] vout_canPeek_315;
  wire [7:0] vout_peek_315;
  wire [0:0] v_316;
  wire [0:0] v_317;
  function [0:0] mux_317(input [0:0] sel);
    case (sel) 0: mux_317 = 1'h0; 1: mux_317 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_318;
  function [0:0] mux_318(input [0:0] sel);
    case (sel) 0: mux_318 = 1'h0; 1: mux_318 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_319;
  wire [0:0] v_320;
  wire [0:0] v_321;
  wire [0:0] v_322;
  wire [0:0] v_323;
  wire [0:0] v_324;
  wire [0:0] v_325;
  function [0:0] mux_325(input [0:0] sel);
    case (sel) 0: mux_325 = 1'h0; 1: mux_325 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_326;
  wire [0:0] v_327;
  wire [0:0] v_328;
  wire [0:0] v_329;
  wire [0:0] v_330;
  function [0:0] mux_330(input [0:0] sel);
    case (sel) 0: mux_330 = 1'h0; 1: mux_330 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_331;
  wire [0:0] v_332;
  wire [0:0] v_333;
  wire [0:0] v_334;
  function [0:0] mux_334(input [0:0] sel);
    case (sel) 0: mux_334 = 1'h0; 1: mux_334 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_335;
  function [0:0] mux_335(input [0:0] sel);
    case (sel) 0: mux_335 = 1'h0; 1: mux_335 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_336 = 1'h0;
  wire [0:0] v_337;
  wire [0:0] v_338;
  wire [0:0] act_339;
  wire [0:0] v_340;
  wire [0:0] v_341;
  wire [0:0] v_342;
  wire [0:0] vin0_consume_en_343;
  wire [0:0] vout_canPeek_343;
  wire [7:0] vout_peek_343;
  wire [0:0] v_344;
  wire [0:0] v_345;
  function [0:0] mux_345(input [0:0] sel);
    case (sel) 0: mux_345 = 1'h0; 1: mux_345 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_346;
  wire [0:0] v_347;
  wire [0:0] v_348;
  wire [0:0] v_349;
  wire [0:0] v_350;
  function [0:0] mux_350(input [0:0] sel);
    case (sel) 0: mux_350 = 1'h0; 1: mux_350 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_351;
  wire [0:0] vin0_consume_en_352;
  wire [0:0] vout_canPeek_352;
  wire [7:0] vout_peek_352;
  wire [0:0] v_353;
  wire [0:0] v_354;
  function [0:0] mux_354(input [0:0] sel);
    case (sel) 0: mux_354 = 1'h0; 1: mux_354 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_355;
  function [0:0] mux_355(input [0:0] sel);
    case (sel) 0: mux_355 = 1'h0; 1: mux_355 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_356;
  wire [0:0] v_357;
  wire [0:0] v_358;
  wire [0:0] v_359;
  wire [0:0] v_360;
  wire [0:0] v_361;
  wire [0:0] v_362;
  function [0:0] mux_362(input [0:0] sel);
    case (sel) 0: mux_362 = 1'h0; 1: mux_362 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_363;
  function [0:0] mux_363(input [0:0] sel);
    case (sel) 0: mux_363 = 1'h0; 1: mux_363 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_364;
  wire [0:0] v_365;
  wire [0:0] v_366;
  wire [0:0] v_367;
  function [0:0] mux_367(input [0:0] sel);
    case (sel) 0: mux_367 = 1'h0; 1: mux_367 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_368;
  function [0:0] mux_368(input [0:0] sel);
    case (sel) 0: mux_368 = 1'h0; 1: mux_368 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_369;
  wire [0:0] v_370;
  wire [0:0] v_371;
  wire [0:0] v_372;
  wire [0:0] v_373;
  wire [0:0] v_374;
  function [0:0] mux_374(input [0:0] sel);
    case (sel) 0: mux_374 = 1'h0; 1: mux_374 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_375;
  function [0:0] mux_375(input [0:0] sel);
    case (sel) 0: mux_375 = 1'h0; 1: mux_375 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_376;
  wire [0:0] v_377;
  wire [0:0] v_378;
  wire [0:0] v_379;
  function [0:0] mux_379(input [0:0] sel);
    case (sel) 0: mux_379 = 1'h0; 1: mux_379 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_380;
  function [0:0] mux_380(input [0:0] sel);
    case (sel) 0: mux_380 = 1'h0; 1: mux_380 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_381;
  wire [0:0] v_382;
  wire [0:0] v_383;
  wire [0:0] v_384;
  wire [0:0] v_385;
  wire [0:0] v_386;
  function [0:0] mux_386(input [0:0] sel);
    case (sel) 0: mux_386 = 1'h0; 1: mux_386 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_387;
  function [0:0] mux_387(input [0:0] sel);
    case (sel) 0: mux_387 = 1'h0; 1: mux_387 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_388;
  wire [0:0] v_389;
  wire [0:0] v_390;
  wire [0:0] v_391;
  function [0:0] mux_391(input [0:0] sel);
    case (sel) 0: mux_391 = 1'h0; 1: mux_391 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_392;
  function [0:0] mux_392(input [0:0] sel);
    case (sel) 0: mux_392 = 1'h0; 1: mux_392 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_393;
  wire [0:0] v_394;
  wire [0:0] v_395;
  wire [0:0] v_396;
  wire [0:0] v_397;
  wire [0:0] v_398;
  function [0:0] mux_398(input [0:0] sel);
    case (sel) 0: mux_398 = 1'h0; 1: mux_398 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_399;
  wire [0:0] v_400;
  wire [0:0] v_401;
  wire [0:0] v_402;
  reg [0:0] v_403 = 1'h0;
  wire [0:0] v_404;
  wire [0:0] v_405;
  wire [0:0] act_406;
  wire [0:0] v_407;
  wire [0:0] v_408;
  wire [0:0] v_409;
  reg [0:0] v_410 = 1'h0;
  wire [0:0] v_411;
  wire [0:0] v_412;
  wire [0:0] act_413;
  wire [0:0] v_414;
  wire [0:0] v_415;
  wire [0:0] v_416;
  reg [0:0] v_417 = 1'h0;
  wire [0:0] v_418;
  wire [0:0] v_419;
  wire [0:0] act_420;
  wire [0:0] v_421;
  wire [0:0] v_422;
  wire [0:0] v_423;
  reg [0:0] v_424 = 1'h0;
  wire [0:0] v_425;
  wire [0:0] v_426;
  wire [0:0] act_427;
  wire [0:0] v_428;
  wire [0:0] v_429;
  wire [0:0] v_430;
  reg [0:0] v_431 = 1'h0;
  wire [0:0] v_432;
  wire [0:0] v_433;
  wire [0:0] act_434;
  wire [0:0] v_435;
  wire [0:0] v_436;
  wire [0:0] v_437;
  wire [0:0] vin0_consume_en_438;
  wire [0:0] vout_canPeek_438;
  wire [7:0] vout_peek_438;
  wire [0:0] v_439;
  wire [0:0] v_440;
  function [0:0] mux_440(input [0:0] sel);
    case (sel) 0: mux_440 = 1'h0; 1: mux_440 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_441;
  wire [0:0] v_442;
  wire [0:0] v_443;
  wire [0:0] v_444;
  wire [0:0] v_445;
  function [0:0] mux_445(input [0:0] sel);
    case (sel) 0: mux_445 = 1'h0; 1: mux_445 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_446;
  wire [0:0] vin0_consume_en_447;
  wire [0:0] vout_canPeek_447;
  wire [7:0] vout_peek_447;
  wire [0:0] v_448;
  wire [0:0] v_449;
  function [0:0] mux_449(input [0:0] sel);
    case (sel) 0: mux_449 = 1'h0; 1: mux_449 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_450;
  function [0:0] mux_450(input [0:0] sel);
    case (sel) 0: mux_450 = 1'h0; 1: mux_450 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_451;
  wire [0:0] v_452;
  wire [0:0] v_453;
  wire [0:0] v_454;
  wire [0:0] v_455;
  wire [0:0] v_456;
  wire [0:0] v_457;
  function [0:0] mux_457(input [0:0] sel);
    case (sel) 0: mux_457 = 1'h0; 1: mux_457 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_458;
  wire [0:0] v_459;
  wire [0:0] v_460;
  wire [0:0] v_461;
  wire [0:0] v_462;
  function [0:0] mux_462(input [0:0] sel);
    case (sel) 0: mux_462 = 1'h0; 1: mux_462 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_463;
  wire [0:0] v_464;
  wire [0:0] v_465;
  wire [0:0] v_466;
  function [0:0] mux_466(input [0:0] sel);
    case (sel) 0: mux_466 = 1'h0; 1: mux_466 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_467;
  function [0:0] mux_467(input [0:0] sel);
    case (sel) 0: mux_467 = 1'h0; 1: mux_467 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_468 = 1'h0;
  wire [0:0] v_469;
  wire [0:0] v_470;
  wire [0:0] act_471;
  wire [0:0] v_472;
  wire [0:0] v_473;
  wire [0:0] v_474;
  wire [0:0] vin0_consume_en_475;
  wire [0:0] vout_canPeek_475;
  wire [7:0] vout_peek_475;
  wire [0:0] v_476;
  wire [0:0] v_477;
  function [0:0] mux_477(input [0:0] sel);
    case (sel) 0: mux_477 = 1'h0; 1: mux_477 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_478;
  wire [0:0] v_479;
  wire [0:0] v_480;
  wire [0:0] v_481;
  wire [0:0] v_482;
  function [0:0] mux_482(input [0:0] sel);
    case (sel) 0: mux_482 = 1'h0; 1: mux_482 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_483;
  wire [0:0] vin0_consume_en_484;
  wire [0:0] vout_canPeek_484;
  wire [7:0] vout_peek_484;
  wire [0:0] v_485;
  wire [0:0] v_486;
  function [0:0] mux_486(input [0:0] sel);
    case (sel) 0: mux_486 = 1'h0; 1: mux_486 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_487;
  function [0:0] mux_487(input [0:0] sel);
    case (sel) 0: mux_487 = 1'h0; 1: mux_487 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_488;
  wire [0:0] v_489;
  wire [0:0] v_490;
  wire [0:0] v_491;
  wire [0:0] v_492;
  wire [0:0] v_493;
  wire [0:0] v_494;
  function [0:0] mux_494(input [0:0] sel);
    case (sel) 0: mux_494 = 1'h0; 1: mux_494 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_495;
  function [0:0] mux_495(input [0:0] sel);
    case (sel) 0: mux_495 = 1'h0; 1: mux_495 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_496;
  wire [0:0] v_497;
  wire [0:0] v_498;
  wire [0:0] v_499;
  function [0:0] mux_499(input [0:0] sel);
    case (sel) 0: mux_499 = 1'h0; 1: mux_499 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_500;
  function [0:0] mux_500(input [0:0] sel);
    case (sel) 0: mux_500 = 1'h0; 1: mux_500 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_501;
  wire [0:0] v_502;
  wire [0:0] v_503;
  wire [0:0] v_504;
  wire [0:0] v_505;
  wire [0:0] v_506;
  function [0:0] mux_506(input [0:0] sel);
    case (sel) 0: mux_506 = 1'h0; 1: mux_506 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_507;
  wire [0:0] v_508;
  wire [0:0] v_509;
  wire [0:0] v_510;
  wire [0:0] v_511;
  function [0:0] mux_511(input [0:0] sel);
    case (sel) 0: mux_511 = 1'h0; 1: mux_511 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_512;
  wire [0:0] v_513;
  wire [0:0] v_514;
  wire [0:0] v_515;
  function [0:0] mux_515(input [0:0] sel);
    case (sel) 0: mux_515 = 1'h0; 1: mux_515 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_516;
  function [0:0] mux_516(input [0:0] sel);
    case (sel) 0: mux_516 = 1'h0; 1: mux_516 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_517 = 1'h0;
  wire [0:0] v_518;
  wire [0:0] v_519;
  wire [0:0] act_520;
  wire [0:0] v_521;
  wire [0:0] v_522;
  wire [0:0] v_523;
  reg [0:0] v_524 = 1'h0;
  wire [0:0] v_525;
  wire [0:0] v_526;
  wire [0:0] act_527;
  wire [0:0] v_528;
  wire [0:0] v_529;
  wire [0:0] v_530;
  wire [0:0] vin0_consume_en_531;
  wire [0:0] vout_canPeek_531;
  wire [7:0] vout_peek_531;
  wire [0:0] v_532;
  wire [0:0] v_533;
  function [0:0] mux_533(input [0:0] sel);
    case (sel) 0: mux_533 = 1'h0; 1: mux_533 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_534;
  wire [0:0] v_535;
  wire [0:0] v_536;
  wire [0:0] v_537;
  wire [0:0] v_538;
  function [0:0] mux_538(input [0:0] sel);
    case (sel) 0: mux_538 = 1'h0; 1: mux_538 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_539;
  wire [0:0] vin0_consume_en_540;
  wire [0:0] vout_canPeek_540;
  wire [7:0] vout_peek_540;
  wire [0:0] v_541;
  wire [0:0] v_542;
  function [0:0] mux_542(input [0:0] sel);
    case (sel) 0: mux_542 = 1'h0; 1: mux_542 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_543;
  function [0:0] mux_543(input [0:0] sel);
    case (sel) 0: mux_543 = 1'h0; 1: mux_543 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_544;
  wire [0:0] v_545;
  wire [0:0] v_546;
  wire [0:0] v_547;
  wire [0:0] v_548;
  wire [0:0] v_549;
  wire [0:0] v_550;
  function [0:0] mux_550(input [0:0] sel);
    case (sel) 0: mux_550 = 1'h0; 1: mux_550 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_551;
  wire [0:0] v_552;
  wire [0:0] v_553;
  wire [0:0] v_554;
  wire [0:0] v_555;
  function [0:0] mux_555(input [0:0] sel);
    case (sel) 0: mux_555 = 1'h0; 1: mux_555 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_556;
  wire [0:0] v_557;
  wire [0:0] v_558;
  wire [0:0] v_559;
  function [0:0] mux_559(input [0:0] sel);
    case (sel) 0: mux_559 = 1'h0; 1: mux_559 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_560;
  function [0:0] mux_560(input [0:0] sel);
    case (sel) 0: mux_560 = 1'h0; 1: mux_560 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_561 = 1'h0;
  wire [0:0] v_562;
  wire [0:0] v_563;
  wire [0:0] act_564;
  wire [0:0] v_565;
  wire [0:0] v_566;
  wire [0:0] v_567;
  wire [0:0] vin0_consume_en_568;
  wire [0:0] vout_canPeek_568;
  wire [7:0] vout_peek_568;
  wire [0:0] v_569;
  wire [0:0] v_570;
  function [0:0] mux_570(input [0:0] sel);
    case (sel) 0: mux_570 = 1'h0; 1: mux_570 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_571;
  wire [0:0] v_572;
  wire [0:0] v_573;
  wire [0:0] v_574;
  wire [0:0] v_575;
  function [0:0] mux_575(input [0:0] sel);
    case (sel) 0: mux_575 = 1'h0; 1: mux_575 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_576;
  wire [0:0] vin0_consume_en_577;
  wire [0:0] vout_canPeek_577;
  wire [7:0] vout_peek_577;
  wire [0:0] v_578;
  wire [0:0] v_579;
  function [0:0] mux_579(input [0:0] sel);
    case (sel) 0: mux_579 = 1'h0; 1: mux_579 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_580;
  function [0:0] mux_580(input [0:0] sel);
    case (sel) 0: mux_580 = 1'h0; 1: mux_580 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_581;
  wire [0:0] v_582;
  wire [0:0] v_583;
  wire [0:0] v_584;
  wire [0:0] v_585;
  wire [0:0] v_586;
  wire [0:0] v_587;
  function [0:0] mux_587(input [0:0] sel);
    case (sel) 0: mux_587 = 1'h0; 1: mux_587 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_588;
  function [0:0] mux_588(input [0:0] sel);
    case (sel) 0: mux_588 = 1'h0; 1: mux_588 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_589;
  wire [0:0] v_590;
  wire [0:0] v_591;
  wire [0:0] v_592;
  function [0:0] mux_592(input [0:0] sel);
    case (sel) 0: mux_592 = 1'h0; 1: mux_592 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_593;
  function [0:0] mux_593(input [0:0] sel);
    case (sel) 0: mux_593 = 1'h0; 1: mux_593 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_594;
  wire [0:0] v_595;
  wire [0:0] v_596;
  wire [0:0] v_597;
  wire [0:0] v_598;
  wire [0:0] v_599;
  function [0:0] mux_599(input [0:0] sel);
    case (sel) 0: mux_599 = 1'h0; 1: mux_599 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_600;
  function [0:0] mux_600(input [0:0] sel);
    case (sel) 0: mux_600 = 1'h0; 1: mux_600 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_601;
  wire [0:0] v_602;
  wire [0:0] v_603;
  wire [0:0] v_604;
  function [0:0] mux_604(input [0:0] sel);
    case (sel) 0: mux_604 = 1'h0; 1: mux_604 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_605;
  function [0:0] mux_605(input [0:0] sel);
    case (sel) 0: mux_605 = 1'h0; 1: mux_605 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_606;
  wire [0:0] v_607;
  wire [0:0] v_608;
  wire [0:0] v_609;
  wire [0:0] v_610;
  wire [0:0] v_611;
  function [0:0] mux_611(input [0:0] sel);
    case (sel) 0: mux_611 = 1'h0; 1: mux_611 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_612;
  wire [0:0] v_613;
  wire [0:0] v_614;
  wire [0:0] v_615;
  wire [0:0] v_616;
  function [0:0] mux_616(input [0:0] sel);
    case (sel) 0: mux_616 = 1'h0; 1: mux_616 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_617;
  wire [0:0] v_618;
  wire [0:0] v_619;
  wire [0:0] v_620;
  function [0:0] mux_620(input [0:0] sel);
    case (sel) 0: mux_620 = 1'h0; 1: mux_620 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_621;
  function [0:0] mux_621(input [0:0] sel);
    case (sel) 0: mux_621 = 1'h0; 1: mux_621 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_622 = 1'h0;
  wire [0:0] v_623;
  wire [0:0] v_624;
  wire [0:0] act_625;
  wire [0:0] v_626;
  wire [0:0] v_627;
  wire [0:0] v_628;
  reg [0:0] v_629 = 1'h0;
  wire [0:0] v_630;
  wire [0:0] v_631;
  wire [0:0] act_632;
  wire [0:0] v_633;
  wire [0:0] v_634;
  wire [0:0] v_635;
  reg [0:0] v_636 = 1'h0;
  wire [0:0] v_637;
  wire [0:0] v_638;
  wire [0:0] act_639;
  wire [0:0] v_640;
  wire [0:0] v_641;
  wire [0:0] v_642;
  wire [0:0] vin0_consume_en_643;
  wire [0:0] vout_canPeek_643;
  wire [7:0] vout_peek_643;
  wire [0:0] v_644;
  wire [0:0] v_645;
  function [0:0] mux_645(input [0:0] sel);
    case (sel) 0: mux_645 = 1'h0; 1: mux_645 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_646;
  wire [0:0] v_647;
  wire [0:0] v_648;
  wire [0:0] v_649;
  wire [0:0] v_650;
  function [0:0] mux_650(input [0:0] sel);
    case (sel) 0: mux_650 = 1'h0; 1: mux_650 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_651;
  wire [0:0] vin0_consume_en_652;
  wire [0:0] vout_canPeek_652;
  wire [7:0] vout_peek_652;
  wire [0:0] v_653;
  wire [0:0] v_654;
  function [0:0] mux_654(input [0:0] sel);
    case (sel) 0: mux_654 = 1'h0; 1: mux_654 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_655;
  function [0:0] mux_655(input [0:0] sel);
    case (sel) 0: mux_655 = 1'h0; 1: mux_655 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_656;
  wire [0:0] v_657;
  wire [0:0] v_658;
  wire [0:0] v_659;
  wire [0:0] v_660;
  wire [0:0] v_661;
  wire [0:0] v_662;
  function [0:0] mux_662(input [0:0] sel);
    case (sel) 0: mux_662 = 1'h0; 1: mux_662 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_663;
  wire [0:0] v_664;
  wire [0:0] v_665;
  wire [0:0] v_666;
  wire [0:0] v_667;
  function [0:0] mux_667(input [0:0] sel);
    case (sel) 0: mux_667 = 1'h0; 1: mux_667 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_668;
  wire [0:0] v_669;
  wire [0:0] v_670;
  wire [0:0] v_671;
  function [0:0] mux_671(input [0:0] sel);
    case (sel) 0: mux_671 = 1'h0; 1: mux_671 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_672;
  function [0:0] mux_672(input [0:0] sel);
    case (sel) 0: mux_672 = 1'h0; 1: mux_672 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_673 = 1'h0;
  wire [0:0] v_674;
  wire [0:0] v_675;
  wire [0:0] act_676;
  wire [0:0] v_677;
  wire [0:0] v_678;
  wire [0:0] v_679;
  wire [0:0] vin0_consume_en_680;
  wire [0:0] vout_canPeek_680;
  wire [7:0] vout_peek_680;
  wire [0:0] v_681;
  wire [0:0] v_682;
  function [0:0] mux_682(input [0:0] sel);
    case (sel) 0: mux_682 = 1'h0; 1: mux_682 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_683;
  wire [0:0] v_684;
  wire [0:0] v_685;
  wire [0:0] v_686;
  wire [0:0] v_687;
  function [0:0] mux_687(input [0:0] sel);
    case (sel) 0: mux_687 = 1'h0; 1: mux_687 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_688;
  wire [0:0] vin0_consume_en_689;
  wire [0:0] vout_canPeek_689;
  wire [7:0] vout_peek_689;
  wire [0:0] v_690;
  wire [0:0] v_691;
  function [0:0] mux_691(input [0:0] sel);
    case (sel) 0: mux_691 = 1'h0; 1: mux_691 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_692;
  function [0:0] mux_692(input [0:0] sel);
    case (sel) 0: mux_692 = 1'h0; 1: mux_692 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_693;
  wire [0:0] v_694;
  wire [0:0] v_695;
  wire [0:0] v_696;
  wire [0:0] v_697;
  wire [0:0] v_698;
  wire [0:0] v_699;
  function [0:0] mux_699(input [0:0] sel);
    case (sel) 0: mux_699 = 1'h0; 1: mux_699 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_700;
  function [0:0] mux_700(input [0:0] sel);
    case (sel) 0: mux_700 = 1'h0; 1: mux_700 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_701;
  wire [0:0] v_702;
  wire [0:0] v_703;
  wire [0:0] v_704;
  function [0:0] mux_704(input [0:0] sel);
    case (sel) 0: mux_704 = 1'h0; 1: mux_704 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_705;
  function [0:0] mux_705(input [0:0] sel);
    case (sel) 0: mux_705 = 1'h0; 1: mux_705 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_706;
  wire [0:0] v_707;
  wire [0:0] v_708;
  wire [0:0] v_709;
  wire [0:0] v_710;
  wire [0:0] v_711;
  function [0:0] mux_711(input [0:0] sel);
    case (sel) 0: mux_711 = 1'h0; 1: mux_711 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_712;
  wire [0:0] v_713;
  wire [0:0] v_714;
  wire [0:0] v_715;
  wire [0:0] v_716;
  function [0:0] mux_716(input [0:0] sel);
    case (sel) 0: mux_716 = 1'h0; 1: mux_716 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_717;
  wire [0:0] v_718;
  wire [0:0] v_719;
  wire [0:0] v_720;
  function [0:0] mux_720(input [0:0] sel);
    case (sel) 0: mux_720 = 1'h0; 1: mux_720 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_721;
  function [0:0] mux_721(input [0:0] sel);
    case (sel) 0: mux_721 = 1'h0; 1: mux_721 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_722 = 1'h0;
  wire [0:0] v_723;
  wire [0:0] v_724;
  wire [0:0] act_725;
  wire [0:0] v_726;
  wire [0:0] v_727;
  wire [0:0] v_728;
  reg [0:0] v_729 = 1'h0;
  wire [0:0] v_730;
  wire [0:0] v_731;
  wire [0:0] act_732;
  wire [0:0] v_733;
  wire [0:0] v_734;
  wire [0:0] v_735;
  wire [0:0] vin0_consume_en_736;
  wire [0:0] vout_canPeek_736;
  wire [7:0] vout_peek_736;
  wire [0:0] v_737;
  wire [0:0] v_738;
  function [0:0] mux_738(input [0:0] sel);
    case (sel) 0: mux_738 = 1'h0; 1: mux_738 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_739;
  wire [0:0] v_740;
  wire [0:0] v_741;
  wire [0:0] v_742;
  wire [0:0] v_743;
  function [0:0] mux_743(input [0:0] sel);
    case (sel) 0: mux_743 = 1'h0; 1: mux_743 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_744;
  wire [0:0] vin0_consume_en_745;
  wire [0:0] vout_canPeek_745;
  wire [7:0] vout_peek_745;
  wire [0:0] v_746;
  wire [0:0] v_747;
  function [0:0] mux_747(input [0:0] sel);
    case (sel) 0: mux_747 = 1'h0; 1: mux_747 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_748;
  function [0:0] mux_748(input [0:0] sel);
    case (sel) 0: mux_748 = 1'h0; 1: mux_748 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_749;
  wire [0:0] v_750;
  wire [0:0] v_751;
  wire [0:0] v_752;
  wire [0:0] v_753;
  wire [0:0] v_754;
  wire [0:0] v_755;
  function [0:0] mux_755(input [0:0] sel);
    case (sel) 0: mux_755 = 1'h0; 1: mux_755 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_756;
  wire [0:0] v_757;
  wire [0:0] v_758;
  wire [0:0] v_759;
  wire [0:0] v_760;
  function [0:0] mux_760(input [0:0] sel);
    case (sel) 0: mux_760 = 1'h0; 1: mux_760 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_761;
  wire [0:0] v_762;
  wire [0:0] v_763;
  wire [0:0] v_764;
  function [0:0] mux_764(input [0:0] sel);
    case (sel) 0: mux_764 = 1'h0; 1: mux_764 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_765;
  function [0:0] mux_765(input [0:0] sel);
    case (sel) 0: mux_765 = 1'h0; 1: mux_765 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_766 = 1'h0;
  wire [0:0] v_767;
  wire [0:0] v_768;
  wire [0:0] act_769;
  wire [0:0] v_770;
  wire [0:0] v_771;
  wire [0:0] v_772;
  wire [0:0] vin0_consume_en_773;
  wire [0:0] vout_canPeek_773;
  wire [7:0] vout_peek_773;
  wire [0:0] v_774;
  wire [0:0] v_775;
  function [0:0] mux_775(input [0:0] sel);
    case (sel) 0: mux_775 = 1'h0; 1: mux_775 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_776;
  wire [0:0] v_777;
  wire [0:0] v_778;
  wire [0:0] v_779;
  wire [0:0] v_780;
  function [0:0] mux_780(input [0:0] sel);
    case (sel) 0: mux_780 = 1'h0; 1: mux_780 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_781;
  wire [0:0] vin0_consume_en_782;
  wire [0:0] vout_canPeek_782;
  wire [7:0] vout_peek_782;
  wire [0:0] v_783;
  wire [0:0] v_784;
  function [0:0] mux_784(input [0:0] sel);
    case (sel) 0: mux_784 = 1'h0; 1: mux_784 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_785;
  function [0:0] mux_785(input [0:0] sel);
    case (sel) 0: mux_785 = 1'h0; 1: mux_785 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_786;
  wire [0:0] v_787;
  wire [0:0] v_788;
  wire [0:0] v_789;
  wire [0:0] v_790;
  wire [0:0] v_791;
  wire [0:0] v_792;
  function [0:0] mux_792(input [0:0] sel);
    case (sel) 0: mux_792 = 1'h0; 1: mux_792 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_793;
  function [0:0] mux_793(input [0:0] sel);
    case (sel) 0: mux_793 = 1'h0; 1: mux_793 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_794;
  wire [0:0] v_795;
  wire [0:0] v_796;
  wire [0:0] v_797;
  function [0:0] mux_797(input [0:0] sel);
    case (sel) 0: mux_797 = 1'h0; 1: mux_797 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_798;
  function [0:0] mux_798(input [0:0] sel);
    case (sel) 0: mux_798 = 1'h0; 1: mux_798 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_799;
  wire [0:0] v_800;
  wire [0:0] v_801;
  wire [0:0] v_802;
  wire [0:0] v_803;
  wire [0:0] v_804;
  function [0:0] mux_804(input [0:0] sel);
    case (sel) 0: mux_804 = 1'h0; 1: mux_804 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_805;
  function [0:0] mux_805(input [0:0] sel);
    case (sel) 0: mux_805 = 1'h0; 1: mux_805 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_806;
  wire [0:0] v_807;
  wire [0:0] v_808;
  wire [0:0] v_809;
  function [0:0] mux_809(input [0:0] sel);
    case (sel) 0: mux_809 = 1'h0; 1: mux_809 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_810;
  function [0:0] mux_810(input [0:0] sel);
    case (sel) 0: mux_810 = 1'h0; 1: mux_810 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_811;
  wire [0:0] v_812;
  wire [0:0] v_813;
  wire [0:0] v_814;
  wire [0:0] v_815;
  wire [0:0] v_816;
  function [0:0] mux_816(input [0:0] sel);
    case (sel) 0: mux_816 = 1'h0; 1: mux_816 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_817;
  function [0:0] mux_817(input [0:0] sel);
    case (sel) 0: mux_817 = 1'h0; 1: mux_817 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_818;
  wire [0:0] v_819;
  wire [0:0] v_820;
  wire [0:0] v_821;
  function [0:0] mux_821(input [0:0] sel);
    case (sel) 0: mux_821 = 1'h0; 1: mux_821 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_822;
  function [0:0] mux_822(input [0:0] sel);
    case (sel) 0: mux_822 = 1'h0; 1: mux_822 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_823;
  wire [0:0] v_824;
  wire [0:0] v_825;
  wire [0:0] v_826;
  wire [0:0] v_827;
  wire [0:0] v_828;
  function [0:0] mux_828(input [0:0] sel);
    case (sel) 0: mux_828 = 1'h0; 1: mux_828 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_829;
  function [0:0] mux_829(input [0:0] sel);
    case (sel) 0: mux_829 = 1'h0; 1: mux_829 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_830;
  wire [0:0] v_831;
  wire [0:0] v_832;
  wire [0:0] v_833;
  function [0:0] mux_833(input [0:0] sel);
    case (sel) 0: mux_833 = 1'h0; 1: mux_833 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_834;
  function [0:0] mux_834(input [0:0] sel);
    case (sel) 0: mux_834 = 1'h0; 1: mux_834 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_835;
  wire [0:0] v_836;
  wire [0:0] v_837;
  wire [0:0] v_838;
  wire [0:0] v_839;
  wire [0:0] v_840;
  function [0:0] mux_840(input [0:0] sel);
    case (sel) 0: mux_840 = 1'h0; 1: mux_840 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_841;
  wire [0:0] v_842;
  wire [0:0] v_843;
  wire [0:0] v_844;
  reg [0:0] v_845 = 1'h0;
  wire [0:0] v_846;
  wire [0:0] v_847;
  wire [0:0] act_848;
  wire [0:0] v_849;
  wire [0:0] v_850;
  wire [0:0] v_851;
  reg [0:0] v_852 = 1'h0;
  wire [0:0] v_853;
  wire [0:0] v_854;
  wire [0:0] act_855;
  wire [0:0] v_856;
  wire [0:0] v_857;
  wire [0:0] v_858;
  reg [0:0] v_859 = 1'h0;
  wire [0:0] v_860;
  wire [0:0] v_861;
  wire [0:0] act_862;
  wire [0:0] v_863;
  wire [0:0] v_864;
  wire [0:0] v_865;
  reg [0:0] v_866 = 1'h0;
  wire [0:0] v_867;
  wire [0:0] v_868;
  wire [0:0] act_869;
  wire [0:0] v_870;
  wire [0:0] v_871;
  wire [0:0] v_872;
  reg [0:0] v_873 = 1'h0;
  wire [0:0] v_874;
  wire [0:0] v_875;
  wire [0:0] act_876;
  wire [0:0] v_877;
  wire [0:0] v_878;
  wire [0:0] v_879;
  reg [0:0] v_880 = 1'h0;
  wire [0:0] v_881;
  wire [0:0] v_882;
  wire [0:0] act_883;
  wire [0:0] v_884;
  wire [0:0] v_885;
  wire [0:0] v_886;
  wire [0:0] vin0_consume_en_887;
  wire [0:0] vout_canPeek_887;
  wire [7:0] vout_peek_887;
  wire [0:0] v_888;
  wire [0:0] v_889;
  function [0:0] mux_889(input [0:0] sel);
    case (sel) 0: mux_889 = 1'h0; 1: mux_889 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_890;
  wire [0:0] v_891;
  wire [0:0] v_892;
  wire [0:0] v_893;
  wire [0:0] v_894;
  function [0:0] mux_894(input [0:0] sel);
    case (sel) 0: mux_894 = 1'h0; 1: mux_894 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_895;
  wire [0:0] vin0_consume_en_896;
  wire [0:0] vout_canPeek_896;
  wire [7:0] vout_peek_896;
  wire [0:0] v_897;
  wire [0:0] v_898;
  function [0:0] mux_898(input [0:0] sel);
    case (sel) 0: mux_898 = 1'h0; 1: mux_898 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_899;
  function [0:0] mux_899(input [0:0] sel);
    case (sel) 0: mux_899 = 1'h0; 1: mux_899 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_900;
  wire [0:0] v_901;
  wire [0:0] v_902;
  wire [0:0] v_903;
  wire [0:0] v_904;
  wire [0:0] v_905;
  wire [0:0] v_906;
  function [0:0] mux_906(input [0:0] sel);
    case (sel) 0: mux_906 = 1'h0; 1: mux_906 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_907;
  wire [0:0] v_908;
  wire [0:0] v_909;
  wire [0:0] v_910;
  wire [0:0] v_911;
  function [0:0] mux_911(input [0:0] sel);
    case (sel) 0: mux_911 = 1'h0; 1: mux_911 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_912;
  wire [0:0] v_913;
  wire [0:0] v_914;
  wire [0:0] v_915;
  function [0:0] mux_915(input [0:0] sel);
    case (sel) 0: mux_915 = 1'h0; 1: mux_915 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_916;
  function [0:0] mux_916(input [0:0] sel);
    case (sel) 0: mux_916 = 1'h0; 1: mux_916 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_917 = 1'h0;
  wire [0:0] v_918;
  wire [0:0] v_919;
  wire [0:0] act_920;
  wire [0:0] v_921;
  wire [0:0] v_922;
  wire [0:0] v_923;
  wire [0:0] vin0_consume_en_924;
  wire [0:0] vout_canPeek_924;
  wire [7:0] vout_peek_924;
  wire [0:0] v_925;
  wire [0:0] v_926;
  function [0:0] mux_926(input [0:0] sel);
    case (sel) 0: mux_926 = 1'h0; 1: mux_926 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_927;
  wire [0:0] v_928;
  wire [0:0] v_929;
  wire [0:0] v_930;
  wire [0:0] v_931;
  function [0:0] mux_931(input [0:0] sel);
    case (sel) 0: mux_931 = 1'h0; 1: mux_931 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_932;
  wire [0:0] vin0_consume_en_933;
  wire [0:0] vout_canPeek_933;
  wire [7:0] vout_peek_933;
  wire [0:0] v_934;
  wire [0:0] v_935;
  function [0:0] mux_935(input [0:0] sel);
    case (sel) 0: mux_935 = 1'h0; 1: mux_935 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_936;
  function [0:0] mux_936(input [0:0] sel);
    case (sel) 0: mux_936 = 1'h0; 1: mux_936 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_937;
  wire [0:0] v_938;
  wire [0:0] v_939;
  wire [0:0] v_940;
  wire [0:0] v_941;
  wire [0:0] v_942;
  wire [0:0] v_943;
  function [0:0] mux_943(input [0:0] sel);
    case (sel) 0: mux_943 = 1'h0; 1: mux_943 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_944;
  function [0:0] mux_944(input [0:0] sel);
    case (sel) 0: mux_944 = 1'h0; 1: mux_944 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_945;
  wire [0:0] v_946;
  wire [0:0] v_947;
  wire [0:0] v_948;
  function [0:0] mux_948(input [0:0] sel);
    case (sel) 0: mux_948 = 1'h0; 1: mux_948 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_949;
  function [0:0] mux_949(input [0:0] sel);
    case (sel) 0: mux_949 = 1'h0; 1: mux_949 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_950;
  wire [0:0] v_951;
  wire [0:0] v_952;
  wire [0:0] v_953;
  wire [0:0] v_954;
  wire [0:0] v_955;
  function [0:0] mux_955(input [0:0] sel);
    case (sel) 0: mux_955 = 1'h0; 1: mux_955 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_956;
  wire [0:0] v_957;
  wire [0:0] v_958;
  wire [0:0] v_959;
  wire [0:0] v_960;
  function [0:0] mux_960(input [0:0] sel);
    case (sel) 0: mux_960 = 1'h0; 1: mux_960 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_961;
  wire [0:0] v_962;
  wire [0:0] v_963;
  wire [0:0] v_964;
  function [0:0] mux_964(input [0:0] sel);
    case (sel) 0: mux_964 = 1'h0; 1: mux_964 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_965;
  function [0:0] mux_965(input [0:0] sel);
    case (sel) 0: mux_965 = 1'h0; 1: mux_965 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_966 = 1'h0;
  wire [0:0] v_967;
  wire [0:0] v_968;
  wire [0:0] act_969;
  wire [0:0] v_970;
  wire [0:0] v_971;
  wire [0:0] v_972;
  reg [0:0] v_973 = 1'h0;
  wire [0:0] v_974;
  wire [0:0] v_975;
  wire [0:0] act_976;
  wire [0:0] v_977;
  wire [0:0] v_978;
  wire [0:0] v_979;
  wire [0:0] vin0_consume_en_980;
  wire [0:0] vout_canPeek_980;
  wire [7:0] vout_peek_980;
  wire [0:0] v_981;
  wire [0:0] v_982;
  function [0:0] mux_982(input [0:0] sel);
    case (sel) 0: mux_982 = 1'h0; 1: mux_982 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_983;
  wire [0:0] v_984;
  wire [0:0] v_985;
  wire [0:0] v_986;
  wire [0:0] v_987;
  function [0:0] mux_987(input [0:0] sel);
    case (sel) 0: mux_987 = 1'h0; 1: mux_987 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_988;
  wire [0:0] vin0_consume_en_989;
  wire [0:0] vout_canPeek_989;
  wire [7:0] vout_peek_989;
  wire [0:0] v_990;
  wire [0:0] v_991;
  function [0:0] mux_991(input [0:0] sel);
    case (sel) 0: mux_991 = 1'h0; 1: mux_991 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_992;
  function [0:0] mux_992(input [0:0] sel);
    case (sel) 0: mux_992 = 1'h0; 1: mux_992 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_993;
  wire [0:0] v_994;
  wire [0:0] v_995;
  wire [0:0] v_996;
  wire [0:0] v_997;
  wire [0:0] v_998;
  wire [0:0] v_999;
  function [0:0] mux_999(input [0:0] sel);
    case (sel) 0: mux_999 = 1'h0; 1: mux_999 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1000;
  wire [0:0] v_1001;
  wire [0:0] v_1002;
  wire [0:0] v_1003;
  wire [0:0] v_1004;
  function [0:0] mux_1004(input [0:0] sel);
    case (sel) 0: mux_1004 = 1'h0; 1: mux_1004 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1005;
  wire [0:0] v_1006;
  wire [0:0] v_1007;
  wire [0:0] v_1008;
  function [0:0] mux_1008(input [0:0] sel);
    case (sel) 0: mux_1008 = 1'h0; 1: mux_1008 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1009;
  function [0:0] mux_1009(input [0:0] sel);
    case (sel) 0: mux_1009 = 1'h0; 1: mux_1009 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_1010 = 1'h0;
  wire [0:0] v_1011;
  wire [0:0] v_1012;
  wire [0:0] act_1013;
  wire [0:0] v_1014;
  wire [0:0] v_1015;
  wire [0:0] v_1016;
  wire [0:0] vin0_consume_en_1017;
  wire [0:0] vout_canPeek_1017;
  wire [7:0] vout_peek_1017;
  wire [0:0] v_1018;
  wire [0:0] v_1019;
  function [0:0] mux_1019(input [0:0] sel);
    case (sel) 0: mux_1019 = 1'h0; 1: mux_1019 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1020;
  wire [0:0] v_1021;
  wire [0:0] v_1022;
  wire [0:0] v_1023;
  wire [0:0] v_1024;
  function [0:0] mux_1024(input [0:0] sel);
    case (sel) 0: mux_1024 = 1'h0; 1: mux_1024 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1025;
  wire [0:0] vin0_consume_en_1026;
  wire [0:0] vout_canPeek_1026;
  wire [7:0] vout_peek_1026;
  wire [0:0] v_1027;
  wire [0:0] v_1028;
  function [0:0] mux_1028(input [0:0] sel);
    case (sel) 0: mux_1028 = 1'h0; 1: mux_1028 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1029;
  function [0:0] mux_1029(input [0:0] sel);
    case (sel) 0: mux_1029 = 1'h0; 1: mux_1029 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1030;
  wire [0:0] v_1031;
  wire [0:0] v_1032;
  wire [0:0] v_1033;
  wire [0:0] v_1034;
  wire [0:0] v_1035;
  wire [0:0] v_1036;
  function [0:0] mux_1036(input [0:0] sel);
    case (sel) 0: mux_1036 = 1'h0; 1: mux_1036 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1037;
  function [0:0] mux_1037(input [0:0] sel);
    case (sel) 0: mux_1037 = 1'h0; 1: mux_1037 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1038;
  wire [0:0] v_1039;
  wire [0:0] v_1040;
  wire [0:0] v_1041;
  function [0:0] mux_1041(input [0:0] sel);
    case (sel) 0: mux_1041 = 1'h0; 1: mux_1041 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1042;
  function [0:0] mux_1042(input [0:0] sel);
    case (sel) 0: mux_1042 = 1'h0; 1: mux_1042 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1043;
  wire [0:0] v_1044;
  wire [0:0] v_1045;
  wire [0:0] v_1046;
  wire [0:0] v_1047;
  wire [0:0] v_1048;
  function [0:0] mux_1048(input [0:0] sel);
    case (sel) 0: mux_1048 = 1'h0; 1: mux_1048 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1049;
  function [0:0] mux_1049(input [0:0] sel);
    case (sel) 0: mux_1049 = 1'h0; 1: mux_1049 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1050;
  wire [0:0] v_1051;
  wire [0:0] v_1052;
  wire [0:0] v_1053;
  function [0:0] mux_1053(input [0:0] sel);
    case (sel) 0: mux_1053 = 1'h0; 1: mux_1053 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1054;
  function [0:0] mux_1054(input [0:0] sel);
    case (sel) 0: mux_1054 = 1'h0; 1: mux_1054 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1055;
  wire [0:0] v_1056;
  wire [0:0] v_1057;
  wire [0:0] v_1058;
  wire [0:0] v_1059;
  wire [0:0] v_1060;
  function [0:0] mux_1060(input [0:0] sel);
    case (sel) 0: mux_1060 = 1'h0; 1: mux_1060 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1061;
  wire [0:0] v_1062;
  wire [0:0] v_1063;
  wire [0:0] v_1064;
  wire [0:0] v_1065;
  function [0:0] mux_1065(input [0:0] sel);
    case (sel) 0: mux_1065 = 1'h0; 1: mux_1065 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1066;
  wire [0:0] v_1067;
  wire [0:0] v_1068;
  wire [0:0] v_1069;
  function [0:0] mux_1069(input [0:0] sel);
    case (sel) 0: mux_1069 = 1'h0; 1: mux_1069 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1070;
  function [0:0] mux_1070(input [0:0] sel);
    case (sel) 0: mux_1070 = 1'h0; 1: mux_1070 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_1071 = 1'h0;
  wire [0:0] v_1072;
  wire [0:0] v_1073;
  wire [0:0] act_1074;
  wire [0:0] v_1075;
  wire [0:0] v_1076;
  wire [0:0] v_1077;
  reg [0:0] v_1078 = 1'h0;
  wire [0:0] v_1079;
  wire [0:0] v_1080;
  wire [0:0] act_1081;
  wire [0:0] v_1082;
  wire [0:0] v_1083;
  wire [0:0] v_1084;
  reg [0:0] v_1085 = 1'h0;
  wire [0:0] v_1086;
  wire [0:0] v_1087;
  wire [0:0] act_1088;
  wire [0:0] v_1089;
  wire [0:0] v_1090;
  wire [0:0] v_1091;
  wire [0:0] vin0_consume_en_1092;
  wire [0:0] vout_canPeek_1092;
  wire [7:0] vout_peek_1092;
  wire [0:0] v_1093;
  wire [0:0] v_1094;
  function [0:0] mux_1094(input [0:0] sel);
    case (sel) 0: mux_1094 = 1'h0; 1: mux_1094 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1095;
  wire [0:0] v_1096;
  wire [0:0] v_1097;
  wire [0:0] v_1098;
  wire [0:0] v_1099;
  function [0:0] mux_1099(input [0:0] sel);
    case (sel) 0: mux_1099 = 1'h0; 1: mux_1099 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1100;
  wire [0:0] vin0_consume_en_1101;
  wire [0:0] vout_canPeek_1101;
  wire [7:0] vout_peek_1101;
  wire [0:0] v_1102;
  wire [0:0] v_1103;
  function [0:0] mux_1103(input [0:0] sel);
    case (sel) 0: mux_1103 = 1'h0; 1: mux_1103 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1104;
  function [0:0] mux_1104(input [0:0] sel);
    case (sel) 0: mux_1104 = 1'h0; 1: mux_1104 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1105;
  wire [0:0] v_1106;
  wire [0:0] v_1107;
  wire [0:0] v_1108;
  wire [0:0] v_1109;
  wire [0:0] v_1110;
  wire [0:0] v_1111;
  function [0:0] mux_1111(input [0:0] sel);
    case (sel) 0: mux_1111 = 1'h0; 1: mux_1111 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1112;
  wire [0:0] v_1113;
  wire [0:0] v_1114;
  wire [0:0] v_1115;
  wire [0:0] v_1116;
  function [0:0] mux_1116(input [0:0] sel);
    case (sel) 0: mux_1116 = 1'h0; 1: mux_1116 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1117;
  wire [0:0] v_1118;
  wire [0:0] v_1119;
  wire [0:0] v_1120;
  function [0:0] mux_1120(input [0:0] sel);
    case (sel) 0: mux_1120 = 1'h0; 1: mux_1120 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1121;
  function [0:0] mux_1121(input [0:0] sel);
    case (sel) 0: mux_1121 = 1'h0; 1: mux_1121 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_1122 = 1'h0;
  wire [0:0] v_1123;
  wire [0:0] v_1124;
  wire [0:0] act_1125;
  wire [0:0] v_1126;
  wire [0:0] v_1127;
  wire [0:0] v_1128;
  wire [0:0] vin0_consume_en_1129;
  wire [0:0] vout_canPeek_1129;
  wire [7:0] vout_peek_1129;
  wire [0:0] v_1130;
  wire [0:0] v_1131;
  function [0:0] mux_1131(input [0:0] sel);
    case (sel) 0: mux_1131 = 1'h0; 1: mux_1131 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1132;
  wire [0:0] v_1133;
  wire [0:0] v_1134;
  wire [0:0] v_1135;
  wire [0:0] v_1136;
  function [0:0] mux_1136(input [0:0] sel);
    case (sel) 0: mux_1136 = 1'h0; 1: mux_1136 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1137;
  wire [0:0] vin0_consume_en_1138;
  wire [0:0] vout_canPeek_1138;
  wire [7:0] vout_peek_1138;
  wire [0:0] v_1139;
  wire [0:0] v_1140;
  function [0:0] mux_1140(input [0:0] sel);
    case (sel) 0: mux_1140 = 1'h0; 1: mux_1140 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1141;
  function [0:0] mux_1141(input [0:0] sel);
    case (sel) 0: mux_1141 = 1'h0; 1: mux_1141 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1142;
  wire [0:0] v_1143;
  wire [0:0] v_1144;
  wire [0:0] v_1145;
  wire [0:0] v_1146;
  wire [0:0] v_1147;
  wire [0:0] v_1148;
  function [0:0] mux_1148(input [0:0] sel);
    case (sel) 0: mux_1148 = 1'h0; 1: mux_1148 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1149;
  function [0:0] mux_1149(input [0:0] sel);
    case (sel) 0: mux_1149 = 1'h0; 1: mux_1149 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1150;
  wire [0:0] v_1151;
  wire [0:0] v_1152;
  wire [0:0] v_1153;
  function [0:0] mux_1153(input [0:0] sel);
    case (sel) 0: mux_1153 = 1'h0; 1: mux_1153 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1154;
  function [0:0] mux_1154(input [0:0] sel);
    case (sel) 0: mux_1154 = 1'h0; 1: mux_1154 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1155;
  wire [0:0] v_1156;
  wire [0:0] v_1157;
  wire [0:0] v_1158;
  wire [0:0] v_1159;
  wire [0:0] v_1160;
  function [0:0] mux_1160(input [0:0] sel);
    case (sel) 0: mux_1160 = 1'h0; 1: mux_1160 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1161;
  wire [0:0] v_1162;
  wire [0:0] v_1163;
  wire [0:0] v_1164;
  wire [0:0] v_1165;
  function [0:0] mux_1165(input [0:0] sel);
    case (sel) 0: mux_1165 = 1'h0; 1: mux_1165 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1166;
  wire [0:0] v_1167;
  wire [0:0] v_1168;
  wire [0:0] v_1169;
  function [0:0] mux_1169(input [0:0] sel);
    case (sel) 0: mux_1169 = 1'h0; 1: mux_1169 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1170;
  function [0:0] mux_1170(input [0:0] sel);
    case (sel) 0: mux_1170 = 1'h0; 1: mux_1170 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_1171 = 1'h0;
  wire [0:0] v_1172;
  wire [0:0] v_1173;
  wire [0:0] act_1174;
  wire [0:0] v_1175;
  wire [0:0] v_1176;
  wire [0:0] v_1177;
  reg [0:0] v_1178 = 1'h0;
  wire [0:0] v_1179;
  wire [0:0] v_1180;
  wire [0:0] act_1181;
  wire [0:0] v_1182;
  wire [0:0] v_1183;
  wire [0:0] v_1184;
  wire [0:0] vin0_consume_en_1185;
  wire [0:0] vout_canPeek_1185;
  wire [7:0] vout_peek_1185;
  wire [0:0] v_1186;
  wire [0:0] v_1187;
  function [0:0] mux_1187(input [0:0] sel);
    case (sel) 0: mux_1187 = 1'h0; 1: mux_1187 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1188;
  wire [0:0] v_1189;
  wire [0:0] v_1190;
  wire [0:0] v_1191;
  wire [0:0] v_1192;
  function [0:0] mux_1192(input [0:0] sel);
    case (sel) 0: mux_1192 = 1'h0; 1: mux_1192 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1193;
  wire [0:0] vin0_consume_en_1194;
  wire [0:0] vout_canPeek_1194;
  wire [7:0] vout_peek_1194;
  wire [0:0] v_1195;
  wire [0:0] v_1196;
  function [0:0] mux_1196(input [0:0] sel);
    case (sel) 0: mux_1196 = 1'h0; 1: mux_1196 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1197;
  function [0:0] mux_1197(input [0:0] sel);
    case (sel) 0: mux_1197 = 1'h0; 1: mux_1197 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1198;
  wire [0:0] v_1199;
  wire [0:0] v_1200;
  wire [0:0] v_1201;
  wire [0:0] v_1202;
  wire [0:0] v_1203;
  wire [0:0] v_1204;
  function [0:0] mux_1204(input [0:0] sel);
    case (sel) 0: mux_1204 = 1'h0; 1: mux_1204 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1205;
  wire [0:0] v_1206;
  wire [0:0] v_1207;
  wire [0:0] v_1208;
  wire [0:0] v_1209;
  function [0:0] mux_1209(input [0:0] sel);
    case (sel) 0: mux_1209 = 1'h0; 1: mux_1209 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1210;
  wire [0:0] v_1211;
  wire [0:0] v_1212;
  wire [0:0] v_1213;
  function [0:0] mux_1213(input [0:0] sel);
    case (sel) 0: mux_1213 = 1'h0; 1: mux_1213 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1214;
  function [0:0] mux_1214(input [0:0] sel);
    case (sel) 0: mux_1214 = 1'h0; 1: mux_1214 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_1215 = 1'h0;
  wire [0:0] v_1216;
  wire [0:0] v_1217;
  wire [0:0] act_1218;
  wire [0:0] v_1219;
  wire [0:0] v_1220;
  wire [0:0] v_1221;
  wire [0:0] vin0_consume_en_1222;
  wire [0:0] vout_canPeek_1222;
  wire [7:0] vout_peek_1222;
  wire [0:0] v_1223;
  wire [0:0] v_1224;
  function [0:0] mux_1224(input [0:0] sel);
    case (sel) 0: mux_1224 = 1'h0; 1: mux_1224 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1225;
  wire [0:0] v_1226;
  wire [0:0] v_1227;
  wire [0:0] v_1228;
  wire [0:0] v_1229;
  function [0:0] mux_1229(input [0:0] sel);
    case (sel) 0: mux_1229 = 1'h0; 1: mux_1229 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1230;
  wire [0:0] vin0_consume_en_1231;
  wire [0:0] vout_canPeek_1231;
  wire [7:0] vout_peek_1231;
  wire [0:0] v_1232;
  wire [0:0] v_1233;
  function [0:0] mux_1233(input [0:0] sel);
    case (sel) 0: mux_1233 = 1'h0; 1: mux_1233 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1234;
  function [0:0] mux_1234(input [0:0] sel);
    case (sel) 0: mux_1234 = 1'h0; 1: mux_1234 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1235;
  wire [0:0] v_1236;
  wire [0:0] v_1237;
  wire [0:0] v_1238;
  wire [0:0] v_1239;
  wire [0:0] v_1240;
  wire [0:0] v_1241;
  function [0:0] mux_1241(input [0:0] sel);
    case (sel) 0: mux_1241 = 1'h0; 1: mux_1241 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1242;
  function [0:0] mux_1242(input [0:0] sel);
    case (sel) 0: mux_1242 = 1'h0; 1: mux_1242 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1243;
  wire [0:0] v_1244;
  wire [0:0] v_1245;
  wire [0:0] v_1246;
  function [0:0] mux_1246(input [0:0] sel);
    case (sel) 0: mux_1246 = 1'h0; 1: mux_1246 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1247;
  function [0:0] mux_1247(input [0:0] sel);
    case (sel) 0: mux_1247 = 1'h0; 1: mux_1247 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1248;
  wire [0:0] v_1249;
  wire [0:0] v_1250;
  wire [0:0] v_1251;
  wire [0:0] v_1252;
  wire [0:0] v_1253;
  function [0:0] mux_1253(input [0:0] sel);
    case (sel) 0: mux_1253 = 1'h0; 1: mux_1253 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1254;
  function [0:0] mux_1254(input [0:0] sel);
    case (sel) 0: mux_1254 = 1'h0; 1: mux_1254 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1255;
  wire [0:0] v_1256;
  wire [0:0] v_1257;
  wire [0:0] v_1258;
  function [0:0] mux_1258(input [0:0] sel);
    case (sel) 0: mux_1258 = 1'h0; 1: mux_1258 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1259;
  function [0:0] mux_1259(input [0:0] sel);
    case (sel) 0: mux_1259 = 1'h0; 1: mux_1259 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1260;
  wire [0:0] v_1261;
  wire [0:0] v_1262;
  wire [0:0] v_1263;
  wire [0:0] v_1264;
  wire [0:0] v_1265;
  function [0:0] mux_1265(input [0:0] sel);
    case (sel) 0: mux_1265 = 1'h0; 1: mux_1265 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1266;
  function [0:0] mux_1266(input [0:0] sel);
    case (sel) 0: mux_1266 = 1'h0; 1: mux_1266 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1267;
  wire [0:0] v_1268;
  wire [0:0] v_1269;
  wire [0:0] v_1270;
  function [0:0] mux_1270(input [0:0] sel);
    case (sel) 0: mux_1270 = 1'h0; 1: mux_1270 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1271;
  function [0:0] mux_1271(input [0:0] sel);
    case (sel) 0: mux_1271 = 1'h0; 1: mux_1271 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1272;
  wire [0:0] v_1273;
  wire [0:0] v_1274;
  wire [0:0] v_1275;
  wire [0:0] v_1276;
  wire [0:0] v_1277;
  function [0:0] mux_1277(input [0:0] sel);
    case (sel) 0: mux_1277 = 1'h0; 1: mux_1277 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1278;
  wire [0:0] v_1279;
  wire [0:0] v_1280;
  wire [0:0] v_1281;
  wire [0:0] v_1282;
  function [0:0] mux_1282(input [0:0] sel);
    case (sel) 0: mux_1282 = 1'h0; 1: mux_1282 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1283;
  wire [0:0] v_1284;
  wire [0:0] v_1285;
  wire [0:0] v_1286;
  function [0:0] mux_1286(input [0:0] sel);
    case (sel) 0: mux_1286 = 1'h0; 1: mux_1286 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1287;
  function [0:0] mux_1287(input [0:0] sel);
    case (sel) 0: mux_1287 = 1'h0; 1: mux_1287 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_1288 = 1'h0;
  wire [0:0] v_1289;
  wire [0:0] v_1290;
  wire [0:0] act_1291;
  wire [0:0] v_1292;
  wire [0:0] v_1293;
  wire [0:0] v_1294;
  reg [0:0] v_1295 = 1'h0;
  wire [0:0] v_1296;
  wire [0:0] v_1297;
  wire [0:0] act_1298;
  wire [0:0] v_1299;
  wire [0:0] v_1300;
  wire [0:0] v_1301;
  reg [0:0] v_1302 = 1'h0;
  wire [0:0] v_1303;
  wire [0:0] v_1304;
  wire [0:0] act_1305;
  wire [0:0] v_1306;
  wire [0:0] v_1307;
  wire [0:0] v_1308;
  reg [0:0] v_1309 = 1'h0;
  wire [0:0] v_1310;
  wire [0:0] v_1311;
  wire [0:0] act_1312;
  wire [0:0] v_1313;
  wire [0:0] v_1314;
  wire [0:0] v_1315;
  wire [0:0] vin0_consume_en_1316;
  wire [0:0] vout_canPeek_1316;
  wire [7:0] vout_peek_1316;
  wire [0:0] v_1317;
  wire [0:0] v_1318;
  function [0:0] mux_1318(input [0:0] sel);
    case (sel) 0: mux_1318 = 1'h0; 1: mux_1318 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1319;
  wire [0:0] v_1320;
  wire [0:0] v_1321;
  wire [0:0] v_1322;
  wire [0:0] v_1323;
  function [0:0] mux_1323(input [0:0] sel);
    case (sel) 0: mux_1323 = 1'h0; 1: mux_1323 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1324;
  wire [0:0] vin0_consume_en_1325;
  wire [0:0] vout_canPeek_1325;
  wire [7:0] vout_peek_1325;
  wire [0:0] v_1326;
  wire [0:0] v_1327;
  function [0:0] mux_1327(input [0:0] sel);
    case (sel) 0: mux_1327 = 1'h0; 1: mux_1327 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1328;
  function [0:0] mux_1328(input [0:0] sel);
    case (sel) 0: mux_1328 = 1'h0; 1: mux_1328 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1329;
  wire [0:0] v_1330;
  wire [0:0] v_1331;
  wire [0:0] v_1332;
  wire [0:0] v_1333;
  wire [0:0] v_1334;
  wire [0:0] v_1335;
  function [0:0] mux_1335(input [0:0] sel);
    case (sel) 0: mux_1335 = 1'h0; 1: mux_1335 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1336;
  wire [0:0] v_1337;
  wire [0:0] v_1338;
  wire [0:0] v_1339;
  wire [0:0] v_1340;
  function [0:0] mux_1340(input [0:0] sel);
    case (sel) 0: mux_1340 = 1'h0; 1: mux_1340 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1341;
  wire [0:0] v_1342;
  wire [0:0] v_1343;
  wire [0:0] v_1344;
  function [0:0] mux_1344(input [0:0] sel);
    case (sel) 0: mux_1344 = 1'h0; 1: mux_1344 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1345;
  function [0:0] mux_1345(input [0:0] sel);
    case (sel) 0: mux_1345 = 1'h0; 1: mux_1345 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_1346 = 1'h0;
  wire [0:0] v_1347;
  wire [0:0] v_1348;
  wire [0:0] act_1349;
  wire [0:0] v_1350;
  wire [0:0] v_1351;
  wire [0:0] v_1352;
  wire [0:0] vin0_consume_en_1353;
  wire [0:0] vout_canPeek_1353;
  wire [7:0] vout_peek_1353;
  wire [0:0] v_1354;
  wire [0:0] v_1355;
  function [0:0] mux_1355(input [0:0] sel);
    case (sel) 0: mux_1355 = 1'h0; 1: mux_1355 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1356;
  wire [0:0] v_1357;
  wire [0:0] v_1358;
  wire [0:0] v_1359;
  wire [0:0] v_1360;
  function [0:0] mux_1360(input [0:0] sel);
    case (sel) 0: mux_1360 = 1'h0; 1: mux_1360 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1361;
  wire [0:0] vin0_consume_en_1362;
  wire [0:0] vout_canPeek_1362;
  wire [7:0] vout_peek_1362;
  wire [0:0] v_1363;
  wire [0:0] v_1364;
  function [0:0] mux_1364(input [0:0] sel);
    case (sel) 0: mux_1364 = 1'h0; 1: mux_1364 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1365;
  function [0:0] mux_1365(input [0:0] sel);
    case (sel) 0: mux_1365 = 1'h0; 1: mux_1365 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1366;
  wire [0:0] v_1367;
  wire [0:0] v_1368;
  wire [0:0] v_1369;
  wire [0:0] v_1370;
  wire [0:0] v_1371;
  wire [0:0] v_1372;
  function [0:0] mux_1372(input [0:0] sel);
    case (sel) 0: mux_1372 = 1'h0; 1: mux_1372 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1373;
  function [0:0] mux_1373(input [0:0] sel);
    case (sel) 0: mux_1373 = 1'h0; 1: mux_1373 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1374;
  wire [0:0] v_1375;
  wire [0:0] v_1376;
  wire [0:0] v_1377;
  function [0:0] mux_1377(input [0:0] sel);
    case (sel) 0: mux_1377 = 1'h0; 1: mux_1377 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1378;
  function [0:0] mux_1378(input [0:0] sel);
    case (sel) 0: mux_1378 = 1'h0; 1: mux_1378 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1379;
  wire [0:0] v_1380;
  wire [0:0] v_1381;
  wire [0:0] v_1382;
  wire [0:0] v_1383;
  wire [0:0] v_1384;
  function [0:0] mux_1384(input [0:0] sel);
    case (sel) 0: mux_1384 = 1'h0; 1: mux_1384 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1385;
  wire [0:0] v_1386;
  wire [0:0] v_1387;
  wire [0:0] v_1388;
  wire [0:0] v_1389;
  function [0:0] mux_1389(input [0:0] sel);
    case (sel) 0: mux_1389 = 1'h0; 1: mux_1389 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1390;
  wire [0:0] v_1391;
  wire [0:0] v_1392;
  wire [0:0] v_1393;
  function [0:0] mux_1393(input [0:0] sel);
    case (sel) 0: mux_1393 = 1'h0; 1: mux_1393 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1394;
  function [0:0] mux_1394(input [0:0] sel);
    case (sel) 0: mux_1394 = 1'h0; 1: mux_1394 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_1395 = 1'h0;
  wire [0:0] v_1396;
  wire [0:0] v_1397;
  wire [0:0] act_1398;
  wire [0:0] v_1399;
  wire [0:0] v_1400;
  wire [0:0] v_1401;
  reg [0:0] v_1402 = 1'h0;
  wire [0:0] v_1403;
  wire [0:0] v_1404;
  wire [0:0] act_1405;
  wire [0:0] v_1406;
  wire [0:0] v_1407;
  wire [0:0] v_1408;
  wire [0:0] vin0_consume_en_1409;
  wire [0:0] vout_canPeek_1409;
  wire [7:0] vout_peek_1409;
  wire [0:0] v_1410;
  wire [0:0] v_1411;
  function [0:0] mux_1411(input [0:0] sel);
    case (sel) 0: mux_1411 = 1'h0; 1: mux_1411 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1412;
  wire [0:0] v_1413;
  wire [0:0] v_1414;
  wire [0:0] v_1415;
  wire [0:0] v_1416;
  function [0:0] mux_1416(input [0:0] sel);
    case (sel) 0: mux_1416 = 1'h0; 1: mux_1416 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1417;
  wire [0:0] vin0_consume_en_1418;
  wire [0:0] vout_canPeek_1418;
  wire [7:0] vout_peek_1418;
  wire [0:0] v_1419;
  wire [0:0] v_1420;
  function [0:0] mux_1420(input [0:0] sel);
    case (sel) 0: mux_1420 = 1'h0; 1: mux_1420 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1421;
  function [0:0] mux_1421(input [0:0] sel);
    case (sel) 0: mux_1421 = 1'h0; 1: mux_1421 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1422;
  wire [0:0] v_1423;
  wire [0:0] v_1424;
  wire [0:0] v_1425;
  wire [0:0] v_1426;
  wire [0:0] v_1427;
  wire [0:0] v_1428;
  function [0:0] mux_1428(input [0:0] sel);
    case (sel) 0: mux_1428 = 1'h0; 1: mux_1428 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1429;
  wire [0:0] v_1430;
  wire [0:0] v_1431;
  wire [0:0] v_1432;
  wire [0:0] v_1433;
  function [0:0] mux_1433(input [0:0] sel);
    case (sel) 0: mux_1433 = 1'h0; 1: mux_1433 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1434;
  wire [0:0] v_1435;
  wire [0:0] v_1436;
  wire [0:0] v_1437;
  function [0:0] mux_1437(input [0:0] sel);
    case (sel) 0: mux_1437 = 1'h0; 1: mux_1437 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1438;
  function [0:0] mux_1438(input [0:0] sel);
    case (sel) 0: mux_1438 = 1'h0; 1: mux_1438 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_1439 = 1'h0;
  wire [0:0] v_1440;
  wire [0:0] v_1441;
  wire [0:0] act_1442;
  wire [0:0] v_1443;
  wire [0:0] v_1444;
  wire [0:0] v_1445;
  wire [0:0] vin0_consume_en_1446;
  wire [0:0] vout_canPeek_1446;
  wire [7:0] vout_peek_1446;
  wire [0:0] v_1447;
  wire [0:0] v_1448;
  function [0:0] mux_1448(input [0:0] sel);
    case (sel) 0: mux_1448 = 1'h0; 1: mux_1448 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1449;
  wire [0:0] v_1450;
  wire [0:0] v_1451;
  wire [0:0] v_1452;
  wire [0:0] v_1453;
  function [0:0] mux_1453(input [0:0] sel);
    case (sel) 0: mux_1453 = 1'h0; 1: mux_1453 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1454;
  wire [0:0] vin0_consume_en_1455;
  wire [0:0] vout_canPeek_1455;
  wire [7:0] vout_peek_1455;
  wire [0:0] v_1456;
  wire [0:0] v_1457;
  function [0:0] mux_1457(input [0:0] sel);
    case (sel) 0: mux_1457 = 1'h0; 1: mux_1457 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1458;
  function [0:0] mux_1458(input [0:0] sel);
    case (sel) 0: mux_1458 = 1'h0; 1: mux_1458 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1459;
  wire [0:0] v_1460;
  wire [0:0] v_1461;
  wire [0:0] v_1462;
  wire [0:0] v_1463;
  wire [0:0] v_1464;
  wire [0:0] v_1465;
  function [0:0] mux_1465(input [0:0] sel);
    case (sel) 0: mux_1465 = 1'h0; 1: mux_1465 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1466;
  function [0:0] mux_1466(input [0:0] sel);
    case (sel) 0: mux_1466 = 1'h0; 1: mux_1466 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1467;
  wire [0:0] v_1468;
  wire [0:0] v_1469;
  wire [0:0] v_1470;
  function [0:0] mux_1470(input [0:0] sel);
    case (sel) 0: mux_1470 = 1'h0; 1: mux_1470 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1471;
  function [0:0] mux_1471(input [0:0] sel);
    case (sel) 0: mux_1471 = 1'h0; 1: mux_1471 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1472;
  wire [0:0] v_1473;
  wire [0:0] v_1474;
  wire [0:0] v_1475;
  wire [0:0] v_1476;
  wire [0:0] v_1477;
  function [0:0] mux_1477(input [0:0] sel);
    case (sel) 0: mux_1477 = 1'h0; 1: mux_1477 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1478;
  function [0:0] mux_1478(input [0:0] sel);
    case (sel) 0: mux_1478 = 1'h0; 1: mux_1478 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1479;
  wire [0:0] v_1480;
  wire [0:0] v_1481;
  wire [0:0] v_1482;
  function [0:0] mux_1482(input [0:0] sel);
    case (sel) 0: mux_1482 = 1'h0; 1: mux_1482 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1483;
  function [0:0] mux_1483(input [0:0] sel);
    case (sel) 0: mux_1483 = 1'h0; 1: mux_1483 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1484;
  wire [0:0] v_1485;
  wire [0:0] v_1486;
  wire [0:0] v_1487;
  wire [0:0] v_1488;
  wire [0:0] v_1489;
  function [0:0] mux_1489(input [0:0] sel);
    case (sel) 0: mux_1489 = 1'h0; 1: mux_1489 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1490;
  wire [0:0] v_1491;
  wire [0:0] v_1492;
  wire [0:0] v_1493;
  wire [0:0] v_1494;
  function [0:0] mux_1494(input [0:0] sel);
    case (sel) 0: mux_1494 = 1'h0; 1: mux_1494 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1495;
  wire [0:0] v_1496;
  wire [0:0] v_1497;
  wire [0:0] v_1498;
  function [0:0] mux_1498(input [0:0] sel);
    case (sel) 0: mux_1498 = 1'h0; 1: mux_1498 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1499;
  function [0:0] mux_1499(input [0:0] sel);
    case (sel) 0: mux_1499 = 1'h0; 1: mux_1499 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_1500 = 1'h0;
  wire [0:0] v_1501;
  wire [0:0] v_1502;
  wire [0:0] act_1503;
  wire [0:0] v_1504;
  wire [0:0] v_1505;
  wire [0:0] v_1506;
  reg [0:0] v_1507 = 1'h0;
  wire [0:0] v_1508;
  wire [0:0] v_1509;
  wire [0:0] act_1510;
  wire [0:0] v_1511;
  wire [0:0] v_1512;
  wire [0:0] v_1513;
  reg [0:0] v_1514 = 1'h0;
  wire [0:0] v_1515;
  wire [0:0] v_1516;
  wire [0:0] act_1517;
  wire [0:0] v_1518;
  wire [0:0] v_1519;
  wire [0:0] v_1520;
  wire [0:0] vin0_consume_en_1521;
  wire [0:0] vout_canPeek_1521;
  wire [7:0] vout_peek_1521;
  wire [0:0] v_1522;
  wire [0:0] v_1523;
  function [0:0] mux_1523(input [0:0] sel);
    case (sel) 0: mux_1523 = 1'h0; 1: mux_1523 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1524;
  wire [0:0] v_1525;
  wire [0:0] v_1526;
  wire [0:0] v_1527;
  wire [0:0] v_1528;
  function [0:0] mux_1528(input [0:0] sel);
    case (sel) 0: mux_1528 = 1'h0; 1: mux_1528 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1529;
  wire [0:0] vin0_consume_en_1530;
  wire [0:0] vout_canPeek_1530;
  wire [7:0] vout_peek_1530;
  wire [0:0] v_1531;
  wire [0:0] v_1532;
  function [0:0] mux_1532(input [0:0] sel);
    case (sel) 0: mux_1532 = 1'h0; 1: mux_1532 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1533;
  function [0:0] mux_1533(input [0:0] sel);
    case (sel) 0: mux_1533 = 1'h0; 1: mux_1533 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1534;
  wire [0:0] v_1535;
  wire [0:0] v_1536;
  wire [0:0] v_1537;
  wire [0:0] v_1538;
  wire [0:0] v_1539;
  wire [0:0] v_1540;
  function [0:0] mux_1540(input [0:0] sel);
    case (sel) 0: mux_1540 = 1'h0; 1: mux_1540 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1541;
  wire [0:0] v_1542;
  wire [0:0] v_1543;
  wire [0:0] v_1544;
  wire [0:0] v_1545;
  function [0:0] mux_1545(input [0:0] sel);
    case (sel) 0: mux_1545 = 1'h0; 1: mux_1545 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1546;
  wire [0:0] v_1547;
  wire [0:0] v_1548;
  wire [0:0] v_1549;
  function [0:0] mux_1549(input [0:0] sel);
    case (sel) 0: mux_1549 = 1'h0; 1: mux_1549 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1550;
  function [0:0] mux_1550(input [0:0] sel);
    case (sel) 0: mux_1550 = 1'h0; 1: mux_1550 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_1551 = 1'h0;
  wire [0:0] v_1552;
  wire [0:0] v_1553;
  wire [0:0] act_1554;
  wire [0:0] v_1555;
  wire [0:0] v_1556;
  wire [0:0] v_1557;
  wire [0:0] vin0_consume_en_1558;
  wire [0:0] vout_canPeek_1558;
  wire [7:0] vout_peek_1558;
  wire [0:0] v_1559;
  wire [0:0] v_1560;
  function [0:0] mux_1560(input [0:0] sel);
    case (sel) 0: mux_1560 = 1'h0; 1: mux_1560 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1561;
  wire [0:0] v_1562;
  wire [0:0] v_1563;
  wire [0:0] v_1564;
  wire [0:0] v_1565;
  function [0:0] mux_1565(input [0:0] sel);
    case (sel) 0: mux_1565 = 1'h0; 1: mux_1565 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1566;
  wire [0:0] vin0_consume_en_1567;
  wire [0:0] vout_canPeek_1567;
  wire [7:0] vout_peek_1567;
  wire [0:0] v_1568;
  wire [0:0] v_1569;
  function [0:0] mux_1569(input [0:0] sel);
    case (sel) 0: mux_1569 = 1'h0; 1: mux_1569 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1570;
  function [0:0] mux_1570(input [0:0] sel);
    case (sel) 0: mux_1570 = 1'h0; 1: mux_1570 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1571;
  wire [0:0] v_1572;
  wire [0:0] v_1573;
  wire [0:0] v_1574;
  wire [0:0] v_1575;
  wire [0:0] v_1576;
  wire [0:0] v_1577;
  function [0:0] mux_1577(input [0:0] sel);
    case (sel) 0: mux_1577 = 1'h0; 1: mux_1577 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1578;
  function [0:0] mux_1578(input [0:0] sel);
    case (sel) 0: mux_1578 = 1'h0; 1: mux_1578 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1579;
  wire [0:0] v_1580;
  wire [0:0] v_1581;
  wire [0:0] v_1582;
  function [0:0] mux_1582(input [0:0] sel);
    case (sel) 0: mux_1582 = 1'h0; 1: mux_1582 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1583;
  function [0:0] mux_1583(input [0:0] sel);
    case (sel) 0: mux_1583 = 1'h0; 1: mux_1583 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1584;
  wire [0:0] v_1585;
  wire [0:0] v_1586;
  wire [0:0] v_1587;
  wire [0:0] v_1588;
  wire [0:0] v_1589;
  function [0:0] mux_1589(input [0:0] sel);
    case (sel) 0: mux_1589 = 1'h0; 1: mux_1589 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1590;
  wire [0:0] v_1591;
  wire [0:0] v_1592;
  wire [0:0] v_1593;
  wire [0:0] v_1594;
  function [0:0] mux_1594(input [0:0] sel);
    case (sel) 0: mux_1594 = 1'h0; 1: mux_1594 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1595;
  wire [0:0] v_1596;
  wire [0:0] v_1597;
  wire [0:0] v_1598;
  function [0:0] mux_1598(input [0:0] sel);
    case (sel) 0: mux_1598 = 1'h0; 1: mux_1598 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1599;
  function [0:0] mux_1599(input [0:0] sel);
    case (sel) 0: mux_1599 = 1'h0; 1: mux_1599 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_1600 = 1'h0;
  wire [0:0] v_1601;
  wire [0:0] v_1602;
  wire [0:0] act_1603;
  wire [0:0] v_1604;
  wire [0:0] v_1605;
  wire [0:0] v_1606;
  reg [0:0] v_1607 = 1'h0;
  wire [0:0] v_1608;
  wire [0:0] v_1609;
  wire [0:0] act_1610;
  wire [0:0] v_1611;
  wire [0:0] v_1612;
  wire [0:0] v_1613;
  wire [0:0] vin0_consume_en_1614;
  wire [0:0] vout_canPeek_1614;
  wire [7:0] vout_peek_1614;
  wire [0:0] v_1615;
  wire [0:0] v_1616;
  function [0:0] mux_1616(input [0:0] sel);
    case (sel) 0: mux_1616 = 1'h0; 1: mux_1616 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1617;
  wire [0:0] v_1618;
  wire [0:0] v_1619;
  wire [0:0] v_1620;
  wire [0:0] v_1621;
  function [0:0] mux_1621(input [0:0] sel);
    case (sel) 0: mux_1621 = 1'h0; 1: mux_1621 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1622;
  wire [0:0] vin0_consume_en_1623;
  wire [0:0] vout_canPeek_1623;
  wire [7:0] vout_peek_1623;
  wire [0:0] v_1624;
  wire [0:0] v_1625;
  function [0:0] mux_1625(input [0:0] sel);
    case (sel) 0: mux_1625 = 1'h0; 1: mux_1625 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1626;
  function [0:0] mux_1626(input [0:0] sel);
    case (sel) 0: mux_1626 = 1'h0; 1: mux_1626 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1627;
  wire [0:0] v_1628;
  wire [0:0] v_1629;
  wire [0:0] v_1630;
  wire [0:0] v_1631;
  wire [0:0] v_1632;
  wire [0:0] v_1633;
  function [0:0] mux_1633(input [0:0] sel);
    case (sel) 0: mux_1633 = 1'h0; 1: mux_1633 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1634;
  wire [0:0] v_1635;
  wire [0:0] v_1636;
  wire [0:0] v_1637;
  wire [0:0] v_1638;
  function [0:0] mux_1638(input [0:0] sel);
    case (sel) 0: mux_1638 = 1'h0; 1: mux_1638 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1639;
  wire [0:0] v_1640;
  wire [0:0] v_1641;
  wire [0:0] v_1642;
  function [0:0] mux_1642(input [0:0] sel);
    case (sel) 0: mux_1642 = 1'h0; 1: mux_1642 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1643;
  function [0:0] mux_1643(input [0:0] sel);
    case (sel) 0: mux_1643 = 1'h0; 1: mux_1643 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_1644 = 1'h0;
  wire [0:0] v_1645;
  wire [0:0] v_1646;
  wire [0:0] act_1647;
  wire [0:0] v_1648;
  wire [0:0] v_1649;
  wire [0:0] v_1650;
  wire [0:0] vin0_consume_en_1651;
  wire [0:0] vout_canPeek_1651;
  wire [7:0] vout_peek_1651;
  wire [0:0] v_1652;
  wire [0:0] v_1653;
  function [0:0] mux_1653(input [0:0] sel);
    case (sel) 0: mux_1653 = 1'h0; 1: mux_1653 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1654;
  wire [0:0] v_1655;
  wire [0:0] v_1656;
  wire [0:0] v_1657;
  wire [0:0] v_1658;
  function [0:0] mux_1658(input [0:0] sel);
    case (sel) 0: mux_1658 = 1'h0; 1: mux_1658 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1659;
  wire [0:0] vin0_consume_en_1660;
  wire [0:0] vout_canPeek_1660;
  wire [7:0] vout_peek_1660;
  wire [0:0] v_1661;
  wire [0:0] v_1662;
  function [0:0] mux_1662(input [0:0] sel);
    case (sel) 0: mux_1662 = 1'h0; 1: mux_1662 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1663;
  function [0:0] mux_1663(input [0:0] sel);
    case (sel) 0: mux_1663 = 1'h0; 1: mux_1663 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1664;
  wire [0:0] v_1665;
  wire [0:0] v_1666;
  wire [0:0] v_1667;
  wire [0:0] v_1668;
  wire [0:0] v_1669;
  wire [0:0] v_1670;
  function [0:0] mux_1670(input [0:0] sel);
    case (sel) 0: mux_1670 = 1'h0; 1: mux_1670 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1671;
  function [0:0] mux_1671(input [0:0] sel);
    case (sel) 0: mux_1671 = 1'h0; 1: mux_1671 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1672;
  wire [0:0] v_1673;
  wire [0:0] v_1674;
  wire [0:0] v_1675;
  function [0:0] mux_1675(input [0:0] sel);
    case (sel) 0: mux_1675 = 1'h0; 1: mux_1675 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1676;
  function [0:0] mux_1676(input [0:0] sel);
    case (sel) 0: mux_1676 = 1'h0; 1: mux_1676 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1677;
  wire [0:0] v_1678;
  wire [0:0] v_1679;
  wire [0:0] v_1680;
  wire [0:0] v_1681;
  wire [0:0] v_1682;
  function [0:0] mux_1682(input [0:0] sel);
    case (sel) 0: mux_1682 = 1'h0; 1: mux_1682 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1683;
  function [0:0] mux_1683(input [0:0] sel);
    case (sel) 0: mux_1683 = 1'h0; 1: mux_1683 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1684;
  wire [0:0] v_1685;
  wire [0:0] v_1686;
  wire [0:0] v_1687;
  function [0:0] mux_1687(input [0:0] sel);
    case (sel) 0: mux_1687 = 1'h0; 1: mux_1687 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1688;
  function [0:0] mux_1688(input [0:0] sel);
    case (sel) 0: mux_1688 = 1'h0; 1: mux_1688 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1689;
  wire [0:0] v_1690;
  wire [0:0] v_1691;
  wire [0:0] v_1692;
  wire [0:0] v_1693;
  wire [0:0] v_1694;
  function [0:0] mux_1694(input [0:0] sel);
    case (sel) 0: mux_1694 = 1'h0; 1: mux_1694 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1695;
  function [0:0] mux_1695(input [0:0] sel);
    case (sel) 0: mux_1695 = 1'h0; 1: mux_1695 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1696;
  wire [0:0] v_1697;
  wire [0:0] v_1698;
  wire [0:0] v_1699;
  function [0:0] mux_1699(input [0:0] sel);
    case (sel) 0: mux_1699 = 1'h0; 1: mux_1699 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1700;
  function [0:0] mux_1700(input [0:0] sel);
    case (sel) 0: mux_1700 = 1'h0; 1: mux_1700 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1701;
  wire [0:0] v_1702;
  wire [0:0] v_1703;
  wire [0:0] v_1704;
  wire [0:0] v_1705;
  wire [0:0] v_1706;
  function [0:0] mux_1706(input [0:0] sel);
    case (sel) 0: mux_1706 = 1'h0; 1: mux_1706 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1707;
  function [0:0] mux_1707(input [0:0] sel);
    case (sel) 0: mux_1707 = 1'h0; 1: mux_1707 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1708;
  wire [0:0] v_1709;
  wire [0:0] v_1710;
  wire [0:0] v_1711;
  function [0:0] mux_1711(input [0:0] sel);
    case (sel) 0: mux_1711 = 1'h0; 1: mux_1711 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1712;
  function [0:0] mux_1712(input [0:0] sel);
    case (sel) 0: mux_1712 = 1'h0; 1: mux_1712 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1713;
  wire [0:0] v_1714;
  wire [0:0] v_1715;
  wire [0:0] v_1716;
  wire [0:0] v_1717;
  wire [0:0] v_1718;
  function [0:0] mux_1718(input [0:0] sel);
    case (sel) 0: mux_1718 = 1'h0; 1: mux_1718 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1719;
  function [0:0] mux_1719(input [0:0] sel);
    case (sel) 0: mux_1719 = 1'h0; 1: mux_1719 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1720;
  wire [0:0] v_1721;
  wire [0:0] v_1722;
  wire [0:0] v_1723;
  function [0:0] mux_1723(input [0:0] sel);
    case (sel) 0: mux_1723 = 1'h0; 1: mux_1723 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1724;
  function [0:0] mux_1724(input [0:0] sel);
    case (sel) 0: mux_1724 = 1'h0; 1: mux_1724 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1725;
  wire [0:0] v_1726;
  wire [0:0] v_1727;
  wire [0:0] v_1728;
  wire [0:0] v_1729;
  wire [0:0] v_1730;
  function [0:0] mux_1730(input [0:0] sel);
    case (sel) 0: mux_1730 = 1'h0; 1: mux_1730 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1731;
  wire [0:0] v_1732;
  wire [0:0] v_1733;
  reg [0:0] v_1734 = 1'h0;
  wire [0:0] v_1735;
  wire [0:0] v_1736;
  wire [0:0] act_1737;
  wire [0:0] v_1738;
  wire [0:0] v_1739;
  wire [0:0] v_1740;
  reg [0:0] v_1741 = 1'h0;
  wire [0:0] v_1742;
  wire [0:0] v_1743;
  wire [0:0] act_1744;
  wire [0:0] v_1745;
  wire [0:0] v_1746;
  wire [0:0] v_1747;
  reg [0:0] v_1748 = 1'h0;
  wire [0:0] v_1749;
  wire [0:0] v_1750;
  wire [0:0] act_1751;
  wire [0:0] v_1752;
  wire [0:0] v_1753;
  wire [0:0] v_1754;
  reg [0:0] v_1755 = 1'h0;
  wire [0:0] v_1756;
  wire [0:0] v_1757;
  wire [0:0] act_1758;
  wire [0:0] v_1759;
  wire [0:0] v_1760;
  wire [0:0] v_1761;
  reg [0:0] v_1762 = 1'h0;
  wire [0:0] v_1763;
  wire [0:0] v_1764;
  wire [0:0] act_1765;
  wire [0:0] v_1766;
  wire [0:0] v_1767;
  wire [0:0] v_1768;
  wire [0:0] vin0_consume_en_1769;
  wire [0:0] vout_canPeek_1769;
  wire [7:0] vout_peek_1769;
  wire [0:0] v_1770;
  wire [0:0] v_1771;
  function [0:0] mux_1771(input [0:0] sel);
    case (sel) 0: mux_1771 = 1'h0; 1: mux_1771 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1772;
  wire [0:0] v_1773;
  wire [0:0] v_1774;
  wire [0:0] v_1775;
  wire [0:0] v_1776;
  function [0:0] mux_1776(input [0:0] sel);
    case (sel) 0: mux_1776 = 1'h0; 1: mux_1776 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1777;
  wire [0:0] vin0_consume_en_1778;
  wire [0:0] vout_canPeek_1778;
  wire [7:0] vout_peek_1778;
  wire [0:0] v_1779;
  wire [0:0] v_1780;
  function [0:0] mux_1780(input [0:0] sel);
    case (sel) 0: mux_1780 = 1'h0; 1: mux_1780 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1781;
  function [0:0] mux_1781(input [0:0] sel);
    case (sel) 0: mux_1781 = 1'h0; 1: mux_1781 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1782;
  wire [0:0] v_1783;
  wire [0:0] v_1784;
  wire [0:0] v_1785;
  wire [0:0] v_1786;
  wire [0:0] v_1787;
  wire [0:0] v_1788;
  function [0:0] mux_1788(input [0:0] sel);
    case (sel) 0: mux_1788 = 1'h0; 1: mux_1788 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1789;
  wire [0:0] v_1790;
  wire [0:0] v_1791;
  wire [0:0] v_1792;
  wire [0:0] v_1793;
  function [0:0] mux_1793(input [0:0] sel);
    case (sel) 0: mux_1793 = 1'h0; 1: mux_1793 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1794;
  wire [0:0] v_1795;
  wire [0:0] v_1796;
  wire [0:0] v_1797;
  function [0:0] mux_1797(input [0:0] sel);
    case (sel) 0: mux_1797 = 1'h0; 1: mux_1797 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1798;
  function [0:0] mux_1798(input [0:0] sel);
    case (sel) 0: mux_1798 = 1'h0; 1: mux_1798 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_1799 = 1'h0;
  wire [0:0] v_1800;
  wire [0:0] v_1801;
  wire [0:0] act_1802;
  wire [0:0] v_1803;
  wire [0:0] v_1804;
  wire [0:0] v_1805;
  wire [0:0] vin0_consume_en_1806;
  wire [0:0] vout_canPeek_1806;
  wire [7:0] vout_peek_1806;
  wire [0:0] v_1807;
  wire [0:0] v_1808;
  function [0:0] mux_1808(input [0:0] sel);
    case (sel) 0: mux_1808 = 1'h0; 1: mux_1808 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1809;
  wire [0:0] v_1810;
  wire [0:0] v_1811;
  wire [0:0] v_1812;
  wire [0:0] v_1813;
  function [0:0] mux_1813(input [0:0] sel);
    case (sel) 0: mux_1813 = 1'h0; 1: mux_1813 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1814;
  wire [0:0] vin0_consume_en_1815;
  wire [0:0] vout_canPeek_1815;
  wire [7:0] vout_peek_1815;
  wire [0:0] v_1816;
  wire [0:0] v_1817;
  function [0:0] mux_1817(input [0:0] sel);
    case (sel) 0: mux_1817 = 1'h0; 1: mux_1817 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1818;
  function [0:0] mux_1818(input [0:0] sel);
    case (sel) 0: mux_1818 = 1'h0; 1: mux_1818 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1819;
  wire [0:0] v_1820;
  wire [0:0] v_1821;
  wire [0:0] v_1822;
  wire [0:0] v_1823;
  wire [0:0] v_1824;
  wire [0:0] v_1825;
  function [0:0] mux_1825(input [0:0] sel);
    case (sel) 0: mux_1825 = 1'h0; 1: mux_1825 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1826;
  function [0:0] mux_1826(input [0:0] sel);
    case (sel) 0: mux_1826 = 1'h0; 1: mux_1826 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1827;
  wire [0:0] v_1828;
  wire [0:0] v_1829;
  wire [0:0] v_1830;
  function [0:0] mux_1830(input [0:0] sel);
    case (sel) 0: mux_1830 = 1'h0; 1: mux_1830 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1831;
  function [0:0] mux_1831(input [0:0] sel);
    case (sel) 0: mux_1831 = 1'h0; 1: mux_1831 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1832;
  wire [0:0] v_1833;
  wire [0:0] v_1834;
  wire [0:0] v_1835;
  wire [0:0] v_1836;
  wire [0:0] v_1837;
  function [0:0] mux_1837(input [0:0] sel);
    case (sel) 0: mux_1837 = 1'h0; 1: mux_1837 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1838;
  wire [0:0] v_1839;
  wire [0:0] v_1840;
  wire [0:0] v_1841;
  wire [0:0] v_1842;
  function [0:0] mux_1842(input [0:0] sel);
    case (sel) 0: mux_1842 = 1'h0; 1: mux_1842 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1843;
  wire [0:0] v_1844;
  wire [0:0] v_1845;
  wire [0:0] v_1846;
  function [0:0] mux_1846(input [0:0] sel);
    case (sel) 0: mux_1846 = 1'h0; 1: mux_1846 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1847;
  function [0:0] mux_1847(input [0:0] sel);
    case (sel) 0: mux_1847 = 1'h0; 1: mux_1847 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_1848 = 1'h0;
  wire [0:0] v_1849;
  wire [0:0] v_1850;
  wire [0:0] act_1851;
  wire [0:0] v_1852;
  wire [0:0] v_1853;
  wire [0:0] v_1854;
  reg [0:0] v_1855 = 1'h0;
  wire [0:0] v_1856;
  wire [0:0] v_1857;
  wire [0:0] act_1858;
  wire [0:0] v_1859;
  wire [0:0] v_1860;
  wire [0:0] v_1861;
  wire [0:0] vin0_consume_en_1862;
  wire [0:0] vout_canPeek_1862;
  wire [7:0] vout_peek_1862;
  wire [0:0] v_1863;
  wire [0:0] v_1864;
  function [0:0] mux_1864(input [0:0] sel);
    case (sel) 0: mux_1864 = 1'h0; 1: mux_1864 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1865;
  wire [0:0] v_1866;
  wire [0:0] v_1867;
  wire [0:0] v_1868;
  wire [0:0] v_1869;
  function [0:0] mux_1869(input [0:0] sel);
    case (sel) 0: mux_1869 = 1'h0; 1: mux_1869 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1870;
  wire [0:0] vin0_consume_en_1871;
  wire [0:0] vout_canPeek_1871;
  wire [7:0] vout_peek_1871;
  wire [0:0] v_1872;
  wire [0:0] v_1873;
  function [0:0] mux_1873(input [0:0] sel);
    case (sel) 0: mux_1873 = 1'h0; 1: mux_1873 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1874;
  function [0:0] mux_1874(input [0:0] sel);
    case (sel) 0: mux_1874 = 1'h0; 1: mux_1874 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1875;
  wire [0:0] v_1876;
  wire [0:0] v_1877;
  wire [0:0] v_1878;
  wire [0:0] v_1879;
  wire [0:0] v_1880;
  wire [0:0] v_1881;
  function [0:0] mux_1881(input [0:0] sel);
    case (sel) 0: mux_1881 = 1'h0; 1: mux_1881 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1882;
  wire [0:0] v_1883;
  wire [0:0] v_1884;
  wire [0:0] v_1885;
  wire [0:0] v_1886;
  function [0:0] mux_1886(input [0:0] sel);
    case (sel) 0: mux_1886 = 1'h0; 1: mux_1886 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1887;
  wire [0:0] v_1888;
  wire [0:0] v_1889;
  wire [0:0] v_1890;
  function [0:0] mux_1890(input [0:0] sel);
    case (sel) 0: mux_1890 = 1'h0; 1: mux_1890 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1891;
  function [0:0] mux_1891(input [0:0] sel);
    case (sel) 0: mux_1891 = 1'h0; 1: mux_1891 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_1892 = 1'h0;
  wire [0:0] v_1893;
  wire [0:0] v_1894;
  wire [0:0] act_1895;
  wire [0:0] v_1896;
  wire [0:0] v_1897;
  wire [0:0] v_1898;
  wire [0:0] vin0_consume_en_1899;
  wire [0:0] vout_canPeek_1899;
  wire [7:0] vout_peek_1899;
  wire [0:0] v_1900;
  wire [0:0] v_1901;
  function [0:0] mux_1901(input [0:0] sel);
    case (sel) 0: mux_1901 = 1'h0; 1: mux_1901 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1902;
  wire [0:0] v_1903;
  wire [0:0] v_1904;
  wire [0:0] v_1905;
  wire [0:0] v_1906;
  function [0:0] mux_1906(input [0:0] sel);
    case (sel) 0: mux_1906 = 1'h0; 1: mux_1906 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1907;
  wire [0:0] vin0_consume_en_1908;
  wire [0:0] vout_canPeek_1908;
  wire [7:0] vout_peek_1908;
  wire [0:0] v_1909;
  wire [0:0] v_1910;
  function [0:0] mux_1910(input [0:0] sel);
    case (sel) 0: mux_1910 = 1'h0; 1: mux_1910 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1911;
  function [0:0] mux_1911(input [0:0] sel);
    case (sel) 0: mux_1911 = 1'h0; 1: mux_1911 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1912;
  wire [0:0] v_1913;
  wire [0:0] v_1914;
  wire [0:0] v_1915;
  wire [0:0] v_1916;
  wire [0:0] v_1917;
  wire [0:0] v_1918;
  function [0:0] mux_1918(input [0:0] sel);
    case (sel) 0: mux_1918 = 1'h0; 1: mux_1918 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1919;
  function [0:0] mux_1919(input [0:0] sel);
    case (sel) 0: mux_1919 = 1'h0; 1: mux_1919 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1920;
  wire [0:0] v_1921;
  wire [0:0] v_1922;
  wire [0:0] v_1923;
  function [0:0] mux_1923(input [0:0] sel);
    case (sel) 0: mux_1923 = 1'h0; 1: mux_1923 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1924;
  function [0:0] mux_1924(input [0:0] sel);
    case (sel) 0: mux_1924 = 1'h0; 1: mux_1924 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1925;
  wire [0:0] v_1926;
  wire [0:0] v_1927;
  wire [0:0] v_1928;
  wire [0:0] v_1929;
  wire [0:0] v_1930;
  function [0:0] mux_1930(input [0:0] sel);
    case (sel) 0: mux_1930 = 1'h0; 1: mux_1930 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1931;
  function [0:0] mux_1931(input [0:0] sel);
    case (sel) 0: mux_1931 = 1'h0; 1: mux_1931 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1932;
  wire [0:0] v_1933;
  wire [0:0] v_1934;
  wire [0:0] v_1935;
  function [0:0] mux_1935(input [0:0] sel);
    case (sel) 0: mux_1935 = 1'h0; 1: mux_1935 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1936;
  function [0:0] mux_1936(input [0:0] sel);
    case (sel) 0: mux_1936 = 1'h0; 1: mux_1936 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1937;
  wire [0:0] v_1938;
  wire [0:0] v_1939;
  wire [0:0] v_1940;
  wire [0:0] v_1941;
  wire [0:0] v_1942;
  function [0:0] mux_1942(input [0:0] sel);
    case (sel) 0: mux_1942 = 1'h0; 1: mux_1942 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1943;
  wire [0:0] v_1944;
  wire [0:0] v_1945;
  wire [0:0] v_1946;
  wire [0:0] v_1947;
  function [0:0] mux_1947(input [0:0] sel);
    case (sel) 0: mux_1947 = 1'h0; 1: mux_1947 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1948;
  wire [0:0] v_1949;
  wire [0:0] v_1950;
  wire [0:0] v_1951;
  function [0:0] mux_1951(input [0:0] sel);
    case (sel) 0: mux_1951 = 1'h0; 1: mux_1951 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1952;
  function [0:0] mux_1952(input [0:0] sel);
    case (sel) 0: mux_1952 = 1'h0; 1: mux_1952 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_1953 = 1'h0;
  wire [0:0] v_1954;
  wire [0:0] v_1955;
  wire [0:0] act_1956;
  wire [0:0] v_1957;
  wire [0:0] v_1958;
  wire [0:0] v_1959;
  reg [0:0] v_1960 = 1'h0;
  wire [0:0] v_1961;
  wire [0:0] v_1962;
  wire [0:0] act_1963;
  wire [0:0] v_1964;
  wire [0:0] v_1965;
  wire [0:0] v_1966;
  reg [0:0] v_1967 = 1'h0;
  wire [0:0] v_1968;
  wire [0:0] v_1969;
  wire [0:0] act_1970;
  wire [0:0] v_1971;
  wire [0:0] v_1972;
  wire [0:0] v_1973;
  wire [0:0] vin0_consume_en_1974;
  wire [0:0] vout_canPeek_1974;
  wire [7:0] vout_peek_1974;
  wire [0:0] v_1975;
  wire [0:0] v_1976;
  function [0:0] mux_1976(input [0:0] sel);
    case (sel) 0: mux_1976 = 1'h0; 1: mux_1976 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1977;
  wire [0:0] v_1978;
  wire [0:0] v_1979;
  wire [0:0] v_1980;
  wire [0:0] v_1981;
  function [0:0] mux_1981(input [0:0] sel);
    case (sel) 0: mux_1981 = 1'h0; 1: mux_1981 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1982;
  wire [0:0] vin0_consume_en_1983;
  wire [0:0] vout_canPeek_1983;
  wire [7:0] vout_peek_1983;
  wire [0:0] v_1984;
  wire [0:0] v_1985;
  function [0:0] mux_1985(input [0:0] sel);
    case (sel) 0: mux_1985 = 1'h0; 1: mux_1985 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1986;
  function [0:0] mux_1986(input [0:0] sel);
    case (sel) 0: mux_1986 = 1'h0; 1: mux_1986 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1987;
  wire [0:0] v_1988;
  wire [0:0] v_1989;
  wire [0:0] v_1990;
  wire [0:0] v_1991;
  wire [0:0] v_1992;
  wire [0:0] v_1993;
  function [0:0] mux_1993(input [0:0] sel);
    case (sel) 0: mux_1993 = 1'h0; 1: mux_1993 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1994;
  wire [0:0] v_1995;
  wire [0:0] v_1996;
  wire [0:0] v_1997;
  wire [0:0] v_1998;
  function [0:0] mux_1998(input [0:0] sel);
    case (sel) 0: mux_1998 = 1'h0; 1: mux_1998 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1999;
  wire [0:0] v_2000;
  wire [0:0] v_2001;
  wire [0:0] v_2002;
  function [0:0] mux_2002(input [0:0] sel);
    case (sel) 0: mux_2002 = 1'h0; 1: mux_2002 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2003;
  function [0:0] mux_2003(input [0:0] sel);
    case (sel) 0: mux_2003 = 1'h0; 1: mux_2003 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2004 = 1'h0;
  wire [0:0] v_2005;
  wire [0:0] v_2006;
  wire [0:0] act_2007;
  wire [0:0] v_2008;
  wire [0:0] v_2009;
  wire [0:0] v_2010;
  wire [0:0] vin0_consume_en_2011;
  wire [0:0] vout_canPeek_2011;
  wire [7:0] vout_peek_2011;
  wire [0:0] v_2012;
  wire [0:0] v_2013;
  function [0:0] mux_2013(input [0:0] sel);
    case (sel) 0: mux_2013 = 1'h0; 1: mux_2013 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2014;
  wire [0:0] v_2015;
  wire [0:0] v_2016;
  wire [0:0] v_2017;
  wire [0:0] v_2018;
  function [0:0] mux_2018(input [0:0] sel);
    case (sel) 0: mux_2018 = 1'h0; 1: mux_2018 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2019;
  wire [0:0] vin0_consume_en_2020;
  wire [0:0] vout_canPeek_2020;
  wire [7:0] vout_peek_2020;
  wire [0:0] v_2021;
  wire [0:0] v_2022;
  function [0:0] mux_2022(input [0:0] sel);
    case (sel) 0: mux_2022 = 1'h0; 1: mux_2022 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2023;
  function [0:0] mux_2023(input [0:0] sel);
    case (sel) 0: mux_2023 = 1'h0; 1: mux_2023 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2024;
  wire [0:0] v_2025;
  wire [0:0] v_2026;
  wire [0:0] v_2027;
  wire [0:0] v_2028;
  wire [0:0] v_2029;
  wire [0:0] v_2030;
  function [0:0] mux_2030(input [0:0] sel);
    case (sel) 0: mux_2030 = 1'h0; 1: mux_2030 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2031;
  function [0:0] mux_2031(input [0:0] sel);
    case (sel) 0: mux_2031 = 1'h0; 1: mux_2031 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2032;
  wire [0:0] v_2033;
  wire [0:0] v_2034;
  wire [0:0] v_2035;
  function [0:0] mux_2035(input [0:0] sel);
    case (sel) 0: mux_2035 = 1'h0; 1: mux_2035 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2036;
  function [0:0] mux_2036(input [0:0] sel);
    case (sel) 0: mux_2036 = 1'h0; 1: mux_2036 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2037;
  wire [0:0] v_2038;
  wire [0:0] v_2039;
  wire [0:0] v_2040;
  wire [0:0] v_2041;
  wire [0:0] v_2042;
  function [0:0] mux_2042(input [0:0] sel);
    case (sel) 0: mux_2042 = 1'h0; 1: mux_2042 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2043;
  wire [0:0] v_2044;
  wire [0:0] v_2045;
  wire [0:0] v_2046;
  wire [0:0] v_2047;
  function [0:0] mux_2047(input [0:0] sel);
    case (sel) 0: mux_2047 = 1'h0; 1: mux_2047 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2048;
  wire [0:0] v_2049;
  wire [0:0] v_2050;
  wire [0:0] v_2051;
  function [0:0] mux_2051(input [0:0] sel);
    case (sel) 0: mux_2051 = 1'h0; 1: mux_2051 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2052;
  function [0:0] mux_2052(input [0:0] sel);
    case (sel) 0: mux_2052 = 1'h0; 1: mux_2052 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2053 = 1'h0;
  wire [0:0] v_2054;
  wire [0:0] v_2055;
  wire [0:0] act_2056;
  wire [0:0] v_2057;
  wire [0:0] v_2058;
  wire [0:0] v_2059;
  reg [0:0] v_2060 = 1'h0;
  wire [0:0] v_2061;
  wire [0:0] v_2062;
  wire [0:0] act_2063;
  wire [0:0] v_2064;
  wire [0:0] v_2065;
  wire [0:0] v_2066;
  wire [0:0] vin0_consume_en_2067;
  wire [0:0] vout_canPeek_2067;
  wire [7:0] vout_peek_2067;
  wire [0:0] v_2068;
  wire [0:0] v_2069;
  function [0:0] mux_2069(input [0:0] sel);
    case (sel) 0: mux_2069 = 1'h0; 1: mux_2069 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2070;
  wire [0:0] v_2071;
  wire [0:0] v_2072;
  wire [0:0] v_2073;
  wire [0:0] v_2074;
  function [0:0] mux_2074(input [0:0] sel);
    case (sel) 0: mux_2074 = 1'h0; 1: mux_2074 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2075;
  wire [0:0] vin0_consume_en_2076;
  wire [0:0] vout_canPeek_2076;
  wire [7:0] vout_peek_2076;
  wire [0:0] v_2077;
  wire [0:0] v_2078;
  function [0:0] mux_2078(input [0:0] sel);
    case (sel) 0: mux_2078 = 1'h0; 1: mux_2078 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2079;
  function [0:0] mux_2079(input [0:0] sel);
    case (sel) 0: mux_2079 = 1'h0; 1: mux_2079 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2080;
  wire [0:0] v_2081;
  wire [0:0] v_2082;
  wire [0:0] v_2083;
  wire [0:0] v_2084;
  wire [0:0] v_2085;
  wire [0:0] v_2086;
  function [0:0] mux_2086(input [0:0] sel);
    case (sel) 0: mux_2086 = 1'h0; 1: mux_2086 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2087;
  wire [0:0] v_2088;
  wire [0:0] v_2089;
  wire [0:0] v_2090;
  wire [0:0] v_2091;
  function [0:0] mux_2091(input [0:0] sel);
    case (sel) 0: mux_2091 = 1'h0; 1: mux_2091 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2092;
  wire [0:0] v_2093;
  wire [0:0] v_2094;
  wire [0:0] v_2095;
  function [0:0] mux_2095(input [0:0] sel);
    case (sel) 0: mux_2095 = 1'h0; 1: mux_2095 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2096;
  function [0:0] mux_2096(input [0:0] sel);
    case (sel) 0: mux_2096 = 1'h0; 1: mux_2096 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2097 = 1'h0;
  wire [0:0] v_2098;
  wire [0:0] v_2099;
  wire [0:0] act_2100;
  wire [0:0] v_2101;
  wire [0:0] v_2102;
  wire [0:0] v_2103;
  wire [0:0] vin0_consume_en_2104;
  wire [0:0] vout_canPeek_2104;
  wire [7:0] vout_peek_2104;
  wire [0:0] v_2105;
  wire [0:0] v_2106;
  function [0:0] mux_2106(input [0:0] sel);
    case (sel) 0: mux_2106 = 1'h0; 1: mux_2106 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2107;
  wire [0:0] v_2108;
  wire [0:0] v_2109;
  wire [0:0] v_2110;
  wire [0:0] v_2111;
  function [0:0] mux_2111(input [0:0] sel);
    case (sel) 0: mux_2111 = 1'h0; 1: mux_2111 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2112;
  wire [0:0] vin0_consume_en_2113;
  wire [0:0] vout_canPeek_2113;
  wire [7:0] vout_peek_2113;
  wire [0:0] v_2114;
  wire [0:0] v_2115;
  function [0:0] mux_2115(input [0:0] sel);
    case (sel) 0: mux_2115 = 1'h0; 1: mux_2115 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2116;
  function [0:0] mux_2116(input [0:0] sel);
    case (sel) 0: mux_2116 = 1'h0; 1: mux_2116 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2117;
  wire [0:0] v_2118;
  wire [0:0] v_2119;
  wire [0:0] v_2120;
  wire [0:0] v_2121;
  wire [0:0] v_2122;
  wire [0:0] v_2123;
  function [0:0] mux_2123(input [0:0] sel);
    case (sel) 0: mux_2123 = 1'h0; 1: mux_2123 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2124;
  function [0:0] mux_2124(input [0:0] sel);
    case (sel) 0: mux_2124 = 1'h0; 1: mux_2124 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2125;
  wire [0:0] v_2126;
  wire [0:0] v_2127;
  wire [0:0] v_2128;
  function [0:0] mux_2128(input [0:0] sel);
    case (sel) 0: mux_2128 = 1'h0; 1: mux_2128 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2129;
  function [0:0] mux_2129(input [0:0] sel);
    case (sel) 0: mux_2129 = 1'h0; 1: mux_2129 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2130;
  wire [0:0] v_2131;
  wire [0:0] v_2132;
  wire [0:0] v_2133;
  wire [0:0] v_2134;
  wire [0:0] v_2135;
  function [0:0] mux_2135(input [0:0] sel);
    case (sel) 0: mux_2135 = 1'h0; 1: mux_2135 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2136;
  function [0:0] mux_2136(input [0:0] sel);
    case (sel) 0: mux_2136 = 1'h0; 1: mux_2136 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2137;
  wire [0:0] v_2138;
  wire [0:0] v_2139;
  wire [0:0] v_2140;
  function [0:0] mux_2140(input [0:0] sel);
    case (sel) 0: mux_2140 = 1'h0; 1: mux_2140 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2141;
  function [0:0] mux_2141(input [0:0] sel);
    case (sel) 0: mux_2141 = 1'h0; 1: mux_2141 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2142;
  wire [0:0] v_2143;
  wire [0:0] v_2144;
  wire [0:0] v_2145;
  wire [0:0] v_2146;
  wire [0:0] v_2147;
  function [0:0] mux_2147(input [0:0] sel);
    case (sel) 0: mux_2147 = 1'h0; 1: mux_2147 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2148;
  function [0:0] mux_2148(input [0:0] sel);
    case (sel) 0: mux_2148 = 1'h0; 1: mux_2148 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2149;
  wire [0:0] v_2150;
  wire [0:0] v_2151;
  wire [0:0] v_2152;
  function [0:0] mux_2152(input [0:0] sel);
    case (sel) 0: mux_2152 = 1'h0; 1: mux_2152 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2153;
  function [0:0] mux_2153(input [0:0] sel);
    case (sel) 0: mux_2153 = 1'h0; 1: mux_2153 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2154;
  wire [0:0] v_2155;
  wire [0:0] v_2156;
  wire [0:0] v_2157;
  wire [0:0] v_2158;
  wire [0:0] v_2159;
  function [0:0] mux_2159(input [0:0] sel);
    case (sel) 0: mux_2159 = 1'h0; 1: mux_2159 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2160;
  wire [0:0] v_2161;
  wire [0:0] v_2162;
  wire [0:0] v_2163;
  wire [0:0] v_2164;
  function [0:0] mux_2164(input [0:0] sel);
    case (sel) 0: mux_2164 = 1'h0; 1: mux_2164 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2165;
  wire [0:0] v_2166;
  wire [0:0] v_2167;
  wire [0:0] v_2168;
  function [0:0] mux_2168(input [0:0] sel);
    case (sel) 0: mux_2168 = 1'h0; 1: mux_2168 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2169;
  function [0:0] mux_2169(input [0:0] sel);
    case (sel) 0: mux_2169 = 1'h0; 1: mux_2169 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2170 = 1'h0;
  wire [0:0] v_2171;
  wire [0:0] v_2172;
  wire [0:0] act_2173;
  wire [0:0] v_2174;
  wire [0:0] v_2175;
  wire [0:0] v_2176;
  reg [0:0] v_2177 = 1'h0;
  wire [0:0] v_2178;
  wire [0:0] v_2179;
  wire [0:0] act_2180;
  wire [0:0] v_2181;
  wire [0:0] v_2182;
  wire [0:0] v_2183;
  reg [0:0] v_2184 = 1'h0;
  wire [0:0] v_2185;
  wire [0:0] v_2186;
  wire [0:0] act_2187;
  wire [0:0] v_2188;
  wire [0:0] v_2189;
  wire [0:0] v_2190;
  reg [0:0] v_2191 = 1'h0;
  wire [0:0] v_2192;
  wire [0:0] v_2193;
  wire [0:0] act_2194;
  wire [0:0] v_2195;
  wire [0:0] v_2196;
  wire [0:0] v_2197;
  wire [0:0] vin0_consume_en_2198;
  wire [0:0] vout_canPeek_2198;
  wire [7:0] vout_peek_2198;
  wire [0:0] v_2199;
  wire [0:0] v_2200;
  function [0:0] mux_2200(input [0:0] sel);
    case (sel) 0: mux_2200 = 1'h0; 1: mux_2200 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2201;
  wire [0:0] v_2202;
  wire [0:0] v_2203;
  wire [0:0] v_2204;
  wire [0:0] v_2205;
  function [0:0] mux_2205(input [0:0] sel);
    case (sel) 0: mux_2205 = 1'h0; 1: mux_2205 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2206;
  wire [0:0] vin0_consume_en_2207;
  wire [0:0] vout_canPeek_2207;
  wire [7:0] vout_peek_2207;
  wire [0:0] v_2208;
  wire [0:0] v_2209;
  function [0:0] mux_2209(input [0:0] sel);
    case (sel) 0: mux_2209 = 1'h0; 1: mux_2209 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2210;
  function [0:0] mux_2210(input [0:0] sel);
    case (sel) 0: mux_2210 = 1'h0; 1: mux_2210 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2211;
  wire [0:0] v_2212;
  wire [0:0] v_2213;
  wire [0:0] v_2214;
  wire [0:0] v_2215;
  wire [0:0] v_2216;
  wire [0:0] v_2217;
  function [0:0] mux_2217(input [0:0] sel);
    case (sel) 0: mux_2217 = 1'h0; 1: mux_2217 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2218;
  wire [0:0] v_2219;
  wire [0:0] v_2220;
  wire [0:0] v_2221;
  wire [0:0] v_2222;
  function [0:0] mux_2222(input [0:0] sel);
    case (sel) 0: mux_2222 = 1'h0; 1: mux_2222 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2223;
  wire [0:0] v_2224;
  wire [0:0] v_2225;
  wire [0:0] v_2226;
  function [0:0] mux_2226(input [0:0] sel);
    case (sel) 0: mux_2226 = 1'h0; 1: mux_2226 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2227;
  function [0:0] mux_2227(input [0:0] sel);
    case (sel) 0: mux_2227 = 1'h0; 1: mux_2227 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2228 = 1'h0;
  wire [0:0] v_2229;
  wire [0:0] v_2230;
  wire [0:0] act_2231;
  wire [0:0] v_2232;
  wire [0:0] v_2233;
  wire [0:0] v_2234;
  wire [0:0] vin0_consume_en_2235;
  wire [0:0] vout_canPeek_2235;
  wire [7:0] vout_peek_2235;
  wire [0:0] v_2236;
  wire [0:0] v_2237;
  function [0:0] mux_2237(input [0:0] sel);
    case (sel) 0: mux_2237 = 1'h0; 1: mux_2237 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2238;
  wire [0:0] v_2239;
  wire [0:0] v_2240;
  wire [0:0] v_2241;
  wire [0:0] v_2242;
  function [0:0] mux_2242(input [0:0] sel);
    case (sel) 0: mux_2242 = 1'h0; 1: mux_2242 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2243;
  wire [0:0] vin0_consume_en_2244;
  wire [0:0] vout_canPeek_2244;
  wire [7:0] vout_peek_2244;
  wire [0:0] v_2245;
  wire [0:0] v_2246;
  function [0:0] mux_2246(input [0:0] sel);
    case (sel) 0: mux_2246 = 1'h0; 1: mux_2246 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2247;
  function [0:0] mux_2247(input [0:0] sel);
    case (sel) 0: mux_2247 = 1'h0; 1: mux_2247 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2248;
  wire [0:0] v_2249;
  wire [0:0] v_2250;
  wire [0:0] v_2251;
  wire [0:0] v_2252;
  wire [0:0] v_2253;
  wire [0:0] v_2254;
  function [0:0] mux_2254(input [0:0] sel);
    case (sel) 0: mux_2254 = 1'h0; 1: mux_2254 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2255;
  function [0:0] mux_2255(input [0:0] sel);
    case (sel) 0: mux_2255 = 1'h0; 1: mux_2255 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2256;
  wire [0:0] v_2257;
  wire [0:0] v_2258;
  wire [0:0] v_2259;
  function [0:0] mux_2259(input [0:0] sel);
    case (sel) 0: mux_2259 = 1'h0; 1: mux_2259 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2260;
  function [0:0] mux_2260(input [0:0] sel);
    case (sel) 0: mux_2260 = 1'h0; 1: mux_2260 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2261;
  wire [0:0] v_2262;
  wire [0:0] v_2263;
  wire [0:0] v_2264;
  wire [0:0] v_2265;
  wire [0:0] v_2266;
  function [0:0] mux_2266(input [0:0] sel);
    case (sel) 0: mux_2266 = 1'h0; 1: mux_2266 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2267;
  wire [0:0] v_2268;
  wire [0:0] v_2269;
  wire [0:0] v_2270;
  wire [0:0] v_2271;
  function [0:0] mux_2271(input [0:0] sel);
    case (sel) 0: mux_2271 = 1'h0; 1: mux_2271 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2272;
  wire [0:0] v_2273;
  wire [0:0] v_2274;
  wire [0:0] v_2275;
  function [0:0] mux_2275(input [0:0] sel);
    case (sel) 0: mux_2275 = 1'h0; 1: mux_2275 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2276;
  function [0:0] mux_2276(input [0:0] sel);
    case (sel) 0: mux_2276 = 1'h0; 1: mux_2276 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2277 = 1'h0;
  wire [0:0] v_2278;
  wire [0:0] v_2279;
  wire [0:0] act_2280;
  wire [0:0] v_2281;
  wire [0:0] v_2282;
  wire [0:0] v_2283;
  reg [0:0] v_2284 = 1'h0;
  wire [0:0] v_2285;
  wire [0:0] v_2286;
  wire [0:0] act_2287;
  wire [0:0] v_2288;
  wire [0:0] v_2289;
  wire [0:0] v_2290;
  wire [0:0] vin0_consume_en_2291;
  wire [0:0] vout_canPeek_2291;
  wire [7:0] vout_peek_2291;
  wire [0:0] v_2292;
  wire [0:0] v_2293;
  function [0:0] mux_2293(input [0:0] sel);
    case (sel) 0: mux_2293 = 1'h0; 1: mux_2293 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2294;
  wire [0:0] v_2295;
  wire [0:0] v_2296;
  wire [0:0] v_2297;
  wire [0:0] v_2298;
  function [0:0] mux_2298(input [0:0] sel);
    case (sel) 0: mux_2298 = 1'h0; 1: mux_2298 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2299;
  wire [0:0] vin0_consume_en_2300;
  wire [0:0] vout_canPeek_2300;
  wire [7:0] vout_peek_2300;
  wire [0:0] v_2301;
  wire [0:0] v_2302;
  function [0:0] mux_2302(input [0:0] sel);
    case (sel) 0: mux_2302 = 1'h0; 1: mux_2302 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2303;
  function [0:0] mux_2303(input [0:0] sel);
    case (sel) 0: mux_2303 = 1'h0; 1: mux_2303 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2304;
  wire [0:0] v_2305;
  wire [0:0] v_2306;
  wire [0:0] v_2307;
  wire [0:0] v_2308;
  wire [0:0] v_2309;
  wire [0:0] v_2310;
  function [0:0] mux_2310(input [0:0] sel);
    case (sel) 0: mux_2310 = 1'h0; 1: mux_2310 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2311;
  wire [0:0] v_2312;
  wire [0:0] v_2313;
  wire [0:0] v_2314;
  wire [0:0] v_2315;
  function [0:0] mux_2315(input [0:0] sel);
    case (sel) 0: mux_2315 = 1'h0; 1: mux_2315 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2316;
  wire [0:0] v_2317;
  wire [0:0] v_2318;
  wire [0:0] v_2319;
  function [0:0] mux_2319(input [0:0] sel);
    case (sel) 0: mux_2319 = 1'h0; 1: mux_2319 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2320;
  function [0:0] mux_2320(input [0:0] sel);
    case (sel) 0: mux_2320 = 1'h0; 1: mux_2320 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2321 = 1'h0;
  wire [0:0] v_2322;
  wire [0:0] v_2323;
  wire [0:0] act_2324;
  wire [0:0] v_2325;
  wire [0:0] v_2326;
  wire [0:0] v_2327;
  wire [0:0] vin0_consume_en_2328;
  wire [0:0] vout_canPeek_2328;
  wire [7:0] vout_peek_2328;
  wire [0:0] v_2329;
  wire [0:0] v_2330;
  function [0:0] mux_2330(input [0:0] sel);
    case (sel) 0: mux_2330 = 1'h0; 1: mux_2330 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2331;
  wire [0:0] v_2332;
  wire [0:0] v_2333;
  wire [0:0] v_2334;
  wire [0:0] v_2335;
  function [0:0] mux_2335(input [0:0] sel);
    case (sel) 0: mux_2335 = 1'h0; 1: mux_2335 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2336;
  wire [0:0] vin0_consume_en_2337;
  wire [0:0] vout_canPeek_2337;
  wire [7:0] vout_peek_2337;
  wire [0:0] v_2338;
  wire [0:0] v_2339;
  function [0:0] mux_2339(input [0:0] sel);
    case (sel) 0: mux_2339 = 1'h0; 1: mux_2339 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2340;
  function [0:0] mux_2340(input [0:0] sel);
    case (sel) 0: mux_2340 = 1'h0; 1: mux_2340 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2341;
  wire [0:0] v_2342;
  wire [0:0] v_2343;
  wire [0:0] v_2344;
  wire [0:0] v_2345;
  wire [0:0] v_2346;
  wire [0:0] v_2347;
  function [0:0] mux_2347(input [0:0] sel);
    case (sel) 0: mux_2347 = 1'h0; 1: mux_2347 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2348;
  function [0:0] mux_2348(input [0:0] sel);
    case (sel) 0: mux_2348 = 1'h0; 1: mux_2348 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2349;
  wire [0:0] v_2350;
  wire [0:0] v_2351;
  wire [0:0] v_2352;
  function [0:0] mux_2352(input [0:0] sel);
    case (sel) 0: mux_2352 = 1'h0; 1: mux_2352 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2353;
  function [0:0] mux_2353(input [0:0] sel);
    case (sel) 0: mux_2353 = 1'h0; 1: mux_2353 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2354;
  wire [0:0] v_2355;
  wire [0:0] v_2356;
  wire [0:0] v_2357;
  wire [0:0] v_2358;
  wire [0:0] v_2359;
  function [0:0] mux_2359(input [0:0] sel);
    case (sel) 0: mux_2359 = 1'h0; 1: mux_2359 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2360;
  function [0:0] mux_2360(input [0:0] sel);
    case (sel) 0: mux_2360 = 1'h0; 1: mux_2360 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2361;
  wire [0:0] v_2362;
  wire [0:0] v_2363;
  wire [0:0] v_2364;
  function [0:0] mux_2364(input [0:0] sel);
    case (sel) 0: mux_2364 = 1'h0; 1: mux_2364 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2365;
  function [0:0] mux_2365(input [0:0] sel);
    case (sel) 0: mux_2365 = 1'h0; 1: mux_2365 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2366;
  wire [0:0] v_2367;
  wire [0:0] v_2368;
  wire [0:0] v_2369;
  wire [0:0] v_2370;
  wire [0:0] v_2371;
  function [0:0] mux_2371(input [0:0] sel);
    case (sel) 0: mux_2371 = 1'h0; 1: mux_2371 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2372;
  wire [0:0] v_2373;
  wire [0:0] v_2374;
  wire [0:0] v_2375;
  wire [0:0] v_2376;
  function [0:0] mux_2376(input [0:0] sel);
    case (sel) 0: mux_2376 = 1'h0; 1: mux_2376 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2377;
  wire [0:0] v_2378;
  wire [0:0] v_2379;
  wire [0:0] v_2380;
  function [0:0] mux_2380(input [0:0] sel);
    case (sel) 0: mux_2380 = 1'h0; 1: mux_2380 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2381;
  function [0:0] mux_2381(input [0:0] sel);
    case (sel) 0: mux_2381 = 1'h0; 1: mux_2381 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2382 = 1'h0;
  wire [0:0] v_2383;
  wire [0:0] v_2384;
  wire [0:0] act_2385;
  wire [0:0] v_2386;
  wire [0:0] v_2387;
  wire [0:0] v_2388;
  reg [0:0] v_2389 = 1'h0;
  wire [0:0] v_2390;
  wire [0:0] v_2391;
  wire [0:0] act_2392;
  wire [0:0] v_2393;
  wire [0:0] v_2394;
  wire [0:0] v_2395;
  reg [0:0] v_2396 = 1'h0;
  wire [0:0] v_2397;
  wire [0:0] v_2398;
  wire [0:0] act_2399;
  wire [0:0] v_2400;
  wire [0:0] v_2401;
  wire [0:0] v_2402;
  wire [0:0] vin0_consume_en_2403;
  wire [0:0] vout_canPeek_2403;
  wire [7:0] vout_peek_2403;
  wire [0:0] v_2404;
  wire [0:0] v_2405;
  function [0:0] mux_2405(input [0:0] sel);
    case (sel) 0: mux_2405 = 1'h0; 1: mux_2405 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2406;
  wire [0:0] v_2407;
  wire [0:0] v_2408;
  wire [0:0] v_2409;
  wire [0:0] v_2410;
  function [0:0] mux_2410(input [0:0] sel);
    case (sel) 0: mux_2410 = 1'h0; 1: mux_2410 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2411;
  wire [0:0] vin0_consume_en_2412;
  wire [0:0] vout_canPeek_2412;
  wire [7:0] vout_peek_2412;
  wire [0:0] v_2413;
  wire [0:0] v_2414;
  function [0:0] mux_2414(input [0:0] sel);
    case (sel) 0: mux_2414 = 1'h0; 1: mux_2414 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2415;
  function [0:0] mux_2415(input [0:0] sel);
    case (sel) 0: mux_2415 = 1'h0; 1: mux_2415 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2416;
  wire [0:0] v_2417;
  wire [0:0] v_2418;
  wire [0:0] v_2419;
  wire [0:0] v_2420;
  wire [0:0] v_2421;
  wire [0:0] v_2422;
  function [0:0] mux_2422(input [0:0] sel);
    case (sel) 0: mux_2422 = 1'h0; 1: mux_2422 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2423;
  wire [0:0] v_2424;
  wire [0:0] v_2425;
  wire [0:0] v_2426;
  wire [0:0] v_2427;
  function [0:0] mux_2427(input [0:0] sel);
    case (sel) 0: mux_2427 = 1'h0; 1: mux_2427 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2428;
  wire [0:0] v_2429;
  wire [0:0] v_2430;
  wire [0:0] v_2431;
  function [0:0] mux_2431(input [0:0] sel);
    case (sel) 0: mux_2431 = 1'h0; 1: mux_2431 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2432;
  function [0:0] mux_2432(input [0:0] sel);
    case (sel) 0: mux_2432 = 1'h0; 1: mux_2432 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2433 = 1'h0;
  wire [0:0] v_2434;
  wire [0:0] v_2435;
  wire [0:0] act_2436;
  wire [0:0] v_2437;
  wire [0:0] v_2438;
  wire [0:0] v_2439;
  wire [0:0] vin0_consume_en_2440;
  wire [0:0] vout_canPeek_2440;
  wire [7:0] vout_peek_2440;
  wire [0:0] v_2441;
  wire [0:0] v_2442;
  function [0:0] mux_2442(input [0:0] sel);
    case (sel) 0: mux_2442 = 1'h0; 1: mux_2442 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2443;
  wire [0:0] v_2444;
  wire [0:0] v_2445;
  wire [0:0] v_2446;
  wire [0:0] v_2447;
  function [0:0] mux_2447(input [0:0] sel);
    case (sel) 0: mux_2447 = 1'h0; 1: mux_2447 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2448;
  wire [0:0] vin0_consume_en_2449;
  wire [0:0] vout_canPeek_2449;
  wire [7:0] vout_peek_2449;
  wire [0:0] v_2450;
  wire [0:0] v_2451;
  function [0:0] mux_2451(input [0:0] sel);
    case (sel) 0: mux_2451 = 1'h0; 1: mux_2451 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2452;
  function [0:0] mux_2452(input [0:0] sel);
    case (sel) 0: mux_2452 = 1'h0; 1: mux_2452 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2453;
  wire [0:0] v_2454;
  wire [0:0] v_2455;
  wire [0:0] v_2456;
  wire [0:0] v_2457;
  wire [0:0] v_2458;
  wire [0:0] v_2459;
  function [0:0] mux_2459(input [0:0] sel);
    case (sel) 0: mux_2459 = 1'h0; 1: mux_2459 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2460;
  function [0:0] mux_2460(input [0:0] sel);
    case (sel) 0: mux_2460 = 1'h0; 1: mux_2460 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2461;
  wire [0:0] v_2462;
  wire [0:0] v_2463;
  wire [0:0] v_2464;
  function [0:0] mux_2464(input [0:0] sel);
    case (sel) 0: mux_2464 = 1'h0; 1: mux_2464 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2465;
  function [0:0] mux_2465(input [0:0] sel);
    case (sel) 0: mux_2465 = 1'h0; 1: mux_2465 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2466;
  wire [0:0] v_2467;
  wire [0:0] v_2468;
  wire [0:0] v_2469;
  wire [0:0] v_2470;
  wire [0:0] v_2471;
  function [0:0] mux_2471(input [0:0] sel);
    case (sel) 0: mux_2471 = 1'h0; 1: mux_2471 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2472;
  wire [0:0] v_2473;
  wire [0:0] v_2474;
  wire [0:0] v_2475;
  wire [0:0] v_2476;
  function [0:0] mux_2476(input [0:0] sel);
    case (sel) 0: mux_2476 = 1'h0; 1: mux_2476 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2477;
  wire [0:0] v_2478;
  wire [0:0] v_2479;
  wire [0:0] v_2480;
  function [0:0] mux_2480(input [0:0] sel);
    case (sel) 0: mux_2480 = 1'h0; 1: mux_2480 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2481;
  function [0:0] mux_2481(input [0:0] sel);
    case (sel) 0: mux_2481 = 1'h0; 1: mux_2481 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2482 = 1'h0;
  wire [0:0] v_2483;
  wire [0:0] v_2484;
  wire [0:0] act_2485;
  wire [0:0] v_2486;
  wire [0:0] v_2487;
  wire [0:0] v_2488;
  reg [0:0] v_2489 = 1'h0;
  wire [0:0] v_2490;
  wire [0:0] v_2491;
  wire [0:0] act_2492;
  wire [0:0] v_2493;
  wire [0:0] v_2494;
  wire [0:0] v_2495;
  wire [0:0] vin0_consume_en_2496;
  wire [0:0] vout_canPeek_2496;
  wire [7:0] vout_peek_2496;
  wire [0:0] v_2497;
  wire [0:0] v_2498;
  function [0:0] mux_2498(input [0:0] sel);
    case (sel) 0: mux_2498 = 1'h0; 1: mux_2498 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2499;
  wire [0:0] v_2500;
  wire [0:0] v_2501;
  wire [0:0] v_2502;
  wire [0:0] v_2503;
  function [0:0] mux_2503(input [0:0] sel);
    case (sel) 0: mux_2503 = 1'h0; 1: mux_2503 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2504;
  wire [0:0] vin0_consume_en_2505;
  wire [0:0] vout_canPeek_2505;
  wire [7:0] vout_peek_2505;
  wire [0:0] v_2506;
  wire [0:0] v_2507;
  function [0:0] mux_2507(input [0:0] sel);
    case (sel) 0: mux_2507 = 1'h0; 1: mux_2507 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2508;
  function [0:0] mux_2508(input [0:0] sel);
    case (sel) 0: mux_2508 = 1'h0; 1: mux_2508 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2509;
  wire [0:0] v_2510;
  wire [0:0] v_2511;
  wire [0:0] v_2512;
  wire [0:0] v_2513;
  wire [0:0] v_2514;
  wire [0:0] v_2515;
  function [0:0] mux_2515(input [0:0] sel);
    case (sel) 0: mux_2515 = 1'h0; 1: mux_2515 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2516;
  wire [0:0] v_2517;
  wire [0:0] v_2518;
  wire [0:0] v_2519;
  wire [0:0] v_2520;
  function [0:0] mux_2520(input [0:0] sel);
    case (sel) 0: mux_2520 = 1'h0; 1: mux_2520 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2521;
  wire [0:0] v_2522;
  wire [0:0] v_2523;
  wire [0:0] v_2524;
  function [0:0] mux_2524(input [0:0] sel);
    case (sel) 0: mux_2524 = 1'h0; 1: mux_2524 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2525;
  function [0:0] mux_2525(input [0:0] sel);
    case (sel) 0: mux_2525 = 1'h0; 1: mux_2525 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2526 = 1'h0;
  wire [0:0] v_2527;
  wire [0:0] v_2528;
  wire [0:0] act_2529;
  wire [0:0] v_2530;
  wire [0:0] v_2531;
  wire [0:0] v_2532;
  wire [0:0] vin0_consume_en_2533;
  wire [0:0] vout_canPeek_2533;
  wire [7:0] vout_peek_2533;
  wire [0:0] v_2534;
  wire [0:0] v_2535;
  function [0:0] mux_2535(input [0:0] sel);
    case (sel) 0: mux_2535 = 1'h0; 1: mux_2535 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2536;
  wire [0:0] v_2537;
  wire [0:0] v_2538;
  wire [0:0] v_2539;
  wire [0:0] v_2540;
  function [0:0] mux_2540(input [0:0] sel);
    case (sel) 0: mux_2540 = 1'h0; 1: mux_2540 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2541;
  wire [0:0] vin0_consume_en_2542;
  wire [0:0] vout_canPeek_2542;
  wire [7:0] vout_peek_2542;
  wire [0:0] v_2543;
  wire [0:0] v_2544;
  function [0:0] mux_2544(input [0:0] sel);
    case (sel) 0: mux_2544 = 1'h0; 1: mux_2544 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2545;
  function [0:0] mux_2545(input [0:0] sel);
    case (sel) 0: mux_2545 = 1'h0; 1: mux_2545 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2546;
  wire [0:0] v_2547;
  wire [0:0] v_2548;
  wire [0:0] v_2549;
  wire [0:0] v_2550;
  wire [0:0] v_2551;
  wire [0:0] v_2552;
  function [0:0] mux_2552(input [0:0] sel);
    case (sel) 0: mux_2552 = 1'h0; 1: mux_2552 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2553;
  function [0:0] mux_2553(input [0:0] sel);
    case (sel) 0: mux_2553 = 1'h0; 1: mux_2553 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2554;
  wire [0:0] v_2555;
  wire [0:0] v_2556;
  wire [0:0] v_2557;
  function [0:0] mux_2557(input [0:0] sel);
    case (sel) 0: mux_2557 = 1'h0; 1: mux_2557 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2558;
  function [0:0] mux_2558(input [0:0] sel);
    case (sel) 0: mux_2558 = 1'h0; 1: mux_2558 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2559;
  wire [0:0] v_2560;
  wire [0:0] v_2561;
  wire [0:0] v_2562;
  wire [0:0] v_2563;
  wire [0:0] v_2564;
  function [0:0] mux_2564(input [0:0] sel);
    case (sel) 0: mux_2564 = 1'h0; 1: mux_2564 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2565;
  function [0:0] mux_2565(input [0:0] sel);
    case (sel) 0: mux_2565 = 1'h0; 1: mux_2565 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2566;
  wire [0:0] v_2567;
  wire [0:0] v_2568;
  wire [0:0] v_2569;
  function [0:0] mux_2569(input [0:0] sel);
    case (sel) 0: mux_2569 = 1'h0; 1: mux_2569 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2570;
  function [0:0] mux_2570(input [0:0] sel);
    case (sel) 0: mux_2570 = 1'h0; 1: mux_2570 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2571;
  wire [0:0] v_2572;
  wire [0:0] v_2573;
  wire [0:0] v_2574;
  wire [0:0] v_2575;
  wire [0:0] v_2576;
  function [0:0] mux_2576(input [0:0] sel);
    case (sel) 0: mux_2576 = 1'h0; 1: mux_2576 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2577;
  function [0:0] mux_2577(input [0:0] sel);
    case (sel) 0: mux_2577 = 1'h0; 1: mux_2577 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2578;
  wire [0:0] v_2579;
  wire [0:0] v_2580;
  wire [0:0] v_2581;
  function [0:0] mux_2581(input [0:0] sel);
    case (sel) 0: mux_2581 = 1'h0; 1: mux_2581 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2582;
  function [0:0] mux_2582(input [0:0] sel);
    case (sel) 0: mux_2582 = 1'h0; 1: mux_2582 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2583;
  wire [0:0] v_2584;
  wire [0:0] v_2585;
  wire [0:0] v_2586;
  wire [0:0] v_2587;
  wire [0:0] v_2588;
  function [0:0] mux_2588(input [0:0] sel);
    case (sel) 0: mux_2588 = 1'h0; 1: mux_2588 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2589;
  function [0:0] mux_2589(input [0:0] sel);
    case (sel) 0: mux_2589 = 1'h0; 1: mux_2589 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2590;
  wire [0:0] v_2591;
  wire [0:0] v_2592;
  wire [0:0] v_2593;
  function [0:0] mux_2593(input [0:0] sel);
    case (sel) 0: mux_2593 = 1'h0; 1: mux_2593 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2594;
  function [0:0] mux_2594(input [0:0] sel);
    case (sel) 0: mux_2594 = 1'h0; 1: mux_2594 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2595;
  wire [0:0] v_2596;
  wire [0:0] v_2597;
  wire [0:0] v_2598;
  wire [0:0] v_2599;
  wire [0:0] v_2600;
  function [0:0] mux_2600(input [0:0] sel);
    case (sel) 0: mux_2600 = 1'h0; 1: mux_2600 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2601;
  wire [0:0] v_2602;
  wire [0:0] v_2603;
  wire [0:0] v_2604;
  reg [0:0] v_2605 = 1'h0;
  wire [0:0] v_2606;
  wire [0:0] v_2607;
  wire [0:0] act_2608;
  wire [0:0] v_2609;
  wire [0:0] v_2610;
  wire [0:0] v_2611;
  wire [0:0] v_2612;
  wire [0:0] v_2613;
  wire [0:0] v_2614;
  function [0:0] mux_2614(input [0:0] sel);
    case (sel) 0: mux_2614 = 1'h0; 1: mux_2614 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2615;
  wire [0:0] v_2616;
  wire [0:0] v_2617;
  reg [0:0] v_2618 = 1'h0;
  wire [0:0] v_2619;
  wire [0:0] v_2620;
  wire [0:0] act_2621;
  wire [0:0] v_2622;
  wire [0:0] v_2623;
  wire [0:0] v_2624;
  reg [0:0] v_2625 = 1'h0;
  wire [0:0] v_2626;
  wire [0:0] v_2627;
  wire [0:0] act_2628;
  wire [0:0] v_2629;
  wire [0:0] v_2630;
  wire [0:0] v_2631;
  reg [0:0] v_2632 = 1'h0;
  wire [0:0] v_2633;
  wire [0:0] v_2634;
  wire [0:0] act_2635;
  wire [0:0] v_2636;
  wire [0:0] v_2637;
  wire [0:0] v_2638;
  reg [0:0] v_2639 = 1'h0;
  wire [0:0] v_2640;
  wire [0:0] v_2641;
  wire [0:0] act_2642;
  wire [0:0] v_2643;
  wire [0:0] v_2644;
  wire [0:0] v_2645;
  reg [0:0] v_2646 = 1'h0;
  wire [0:0] v_2647;
  wire [0:0] v_2648;
  wire [0:0] act_2649;
  wire [0:0] v_2650;
  wire [0:0] v_2651;
  wire [0:0] v_2652;
  reg [0:0] v_2653 = 1'h0;
  wire [0:0] v_2654;
  wire [0:0] v_2655;
  wire [0:0] act_2656;
  wire [0:0] v_2657;
  wire [0:0] v_2658;
  wire [0:0] v_2659;
  wire [0:0] vin0_consume_en_2660;
  wire [0:0] vout_canPeek_2660;
  wire [7:0] vout_peek_2660;
  wire [0:0] v_2661;
  wire [0:0] v_2662;
  function [0:0] mux_2662(input [0:0] sel);
    case (sel) 0: mux_2662 = 1'h0; 1: mux_2662 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2663;
  wire [0:0] v_2664;
  wire [0:0] v_2665;
  wire [0:0] v_2666;
  wire [0:0] v_2667;
  function [0:0] mux_2667(input [0:0] sel);
    case (sel) 0: mux_2667 = 1'h0; 1: mux_2667 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2668;
  wire [0:0] vin0_consume_en_2669;
  wire [0:0] vout_canPeek_2669;
  wire [7:0] vout_peek_2669;
  wire [0:0] v_2670;
  wire [0:0] v_2671;
  function [0:0] mux_2671(input [0:0] sel);
    case (sel) 0: mux_2671 = 1'h0; 1: mux_2671 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2672;
  function [0:0] mux_2672(input [0:0] sel);
    case (sel) 0: mux_2672 = 1'h0; 1: mux_2672 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2673;
  wire [0:0] v_2674;
  wire [0:0] v_2675;
  wire [0:0] v_2676;
  wire [0:0] v_2677;
  wire [0:0] v_2678;
  wire [0:0] v_2679;
  function [0:0] mux_2679(input [0:0] sel);
    case (sel) 0: mux_2679 = 1'h0; 1: mux_2679 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2680;
  wire [0:0] v_2681;
  wire [0:0] v_2682;
  wire [0:0] v_2683;
  wire [0:0] v_2684;
  function [0:0] mux_2684(input [0:0] sel);
    case (sel) 0: mux_2684 = 1'h0; 1: mux_2684 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2685;
  wire [0:0] v_2686;
  wire [0:0] v_2687;
  wire [0:0] v_2688;
  function [0:0] mux_2688(input [0:0] sel);
    case (sel) 0: mux_2688 = 1'h0; 1: mux_2688 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2689;
  function [0:0] mux_2689(input [0:0] sel);
    case (sel) 0: mux_2689 = 1'h0; 1: mux_2689 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2690 = 1'h0;
  wire [0:0] v_2691;
  wire [0:0] v_2692;
  wire [0:0] act_2693;
  wire [0:0] v_2694;
  wire [0:0] v_2695;
  wire [0:0] v_2696;
  wire [0:0] vin0_consume_en_2697;
  wire [0:0] vout_canPeek_2697;
  wire [7:0] vout_peek_2697;
  wire [0:0] v_2698;
  wire [0:0] v_2699;
  function [0:0] mux_2699(input [0:0] sel);
    case (sel) 0: mux_2699 = 1'h0; 1: mux_2699 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2700;
  wire [0:0] v_2701;
  wire [0:0] v_2702;
  wire [0:0] v_2703;
  wire [0:0] v_2704;
  function [0:0] mux_2704(input [0:0] sel);
    case (sel) 0: mux_2704 = 1'h0; 1: mux_2704 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2705;
  wire [0:0] vin0_consume_en_2706;
  wire [0:0] vout_canPeek_2706;
  wire [7:0] vout_peek_2706;
  wire [0:0] v_2707;
  wire [0:0] v_2708;
  function [0:0] mux_2708(input [0:0] sel);
    case (sel) 0: mux_2708 = 1'h0; 1: mux_2708 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2709;
  function [0:0] mux_2709(input [0:0] sel);
    case (sel) 0: mux_2709 = 1'h0; 1: mux_2709 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2710;
  wire [0:0] v_2711;
  wire [0:0] v_2712;
  wire [0:0] v_2713;
  wire [0:0] v_2714;
  wire [0:0] v_2715;
  wire [0:0] v_2716;
  function [0:0] mux_2716(input [0:0] sel);
    case (sel) 0: mux_2716 = 1'h0; 1: mux_2716 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2717;
  function [0:0] mux_2717(input [0:0] sel);
    case (sel) 0: mux_2717 = 1'h0; 1: mux_2717 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2718;
  wire [0:0] v_2719;
  wire [0:0] v_2720;
  wire [0:0] v_2721;
  function [0:0] mux_2721(input [0:0] sel);
    case (sel) 0: mux_2721 = 1'h0; 1: mux_2721 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2722;
  function [0:0] mux_2722(input [0:0] sel);
    case (sel) 0: mux_2722 = 1'h0; 1: mux_2722 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2723;
  wire [0:0] v_2724;
  wire [0:0] v_2725;
  wire [0:0] v_2726;
  wire [0:0] v_2727;
  wire [0:0] v_2728;
  function [0:0] mux_2728(input [0:0] sel);
    case (sel) 0: mux_2728 = 1'h0; 1: mux_2728 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2729;
  wire [0:0] v_2730;
  wire [0:0] v_2731;
  wire [0:0] v_2732;
  wire [0:0] v_2733;
  function [0:0] mux_2733(input [0:0] sel);
    case (sel) 0: mux_2733 = 1'h0; 1: mux_2733 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2734;
  wire [0:0] v_2735;
  wire [0:0] v_2736;
  wire [0:0] v_2737;
  function [0:0] mux_2737(input [0:0] sel);
    case (sel) 0: mux_2737 = 1'h0; 1: mux_2737 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2738;
  function [0:0] mux_2738(input [0:0] sel);
    case (sel) 0: mux_2738 = 1'h0; 1: mux_2738 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2739 = 1'h0;
  wire [0:0] v_2740;
  wire [0:0] v_2741;
  wire [0:0] act_2742;
  wire [0:0] v_2743;
  wire [0:0] v_2744;
  wire [0:0] v_2745;
  reg [0:0] v_2746 = 1'h0;
  wire [0:0] v_2747;
  wire [0:0] v_2748;
  wire [0:0] act_2749;
  wire [0:0] v_2750;
  wire [0:0] v_2751;
  wire [0:0] v_2752;
  wire [0:0] vin0_consume_en_2753;
  wire [0:0] vout_canPeek_2753;
  wire [7:0] vout_peek_2753;
  wire [0:0] v_2754;
  wire [0:0] v_2755;
  function [0:0] mux_2755(input [0:0] sel);
    case (sel) 0: mux_2755 = 1'h0; 1: mux_2755 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2756;
  wire [0:0] v_2757;
  wire [0:0] v_2758;
  wire [0:0] v_2759;
  wire [0:0] v_2760;
  function [0:0] mux_2760(input [0:0] sel);
    case (sel) 0: mux_2760 = 1'h0; 1: mux_2760 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2761;
  wire [0:0] vin0_consume_en_2762;
  wire [0:0] vout_canPeek_2762;
  wire [7:0] vout_peek_2762;
  wire [0:0] v_2763;
  wire [0:0] v_2764;
  function [0:0] mux_2764(input [0:0] sel);
    case (sel) 0: mux_2764 = 1'h0; 1: mux_2764 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2765;
  function [0:0] mux_2765(input [0:0] sel);
    case (sel) 0: mux_2765 = 1'h0; 1: mux_2765 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2766;
  wire [0:0] v_2767;
  wire [0:0] v_2768;
  wire [0:0] v_2769;
  wire [0:0] v_2770;
  wire [0:0] v_2771;
  wire [0:0] v_2772;
  function [0:0] mux_2772(input [0:0] sel);
    case (sel) 0: mux_2772 = 1'h0; 1: mux_2772 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2773;
  wire [0:0] v_2774;
  wire [0:0] v_2775;
  wire [0:0] v_2776;
  wire [0:0] v_2777;
  function [0:0] mux_2777(input [0:0] sel);
    case (sel) 0: mux_2777 = 1'h0; 1: mux_2777 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2778;
  wire [0:0] v_2779;
  wire [0:0] v_2780;
  wire [0:0] v_2781;
  function [0:0] mux_2781(input [0:0] sel);
    case (sel) 0: mux_2781 = 1'h0; 1: mux_2781 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2782;
  function [0:0] mux_2782(input [0:0] sel);
    case (sel) 0: mux_2782 = 1'h0; 1: mux_2782 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2783 = 1'h0;
  wire [0:0] v_2784;
  wire [0:0] v_2785;
  wire [0:0] act_2786;
  wire [0:0] v_2787;
  wire [0:0] v_2788;
  wire [0:0] v_2789;
  wire [0:0] vin0_consume_en_2790;
  wire [0:0] vout_canPeek_2790;
  wire [7:0] vout_peek_2790;
  wire [0:0] v_2791;
  wire [0:0] v_2792;
  function [0:0] mux_2792(input [0:0] sel);
    case (sel) 0: mux_2792 = 1'h0; 1: mux_2792 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2793;
  wire [0:0] v_2794;
  wire [0:0] v_2795;
  wire [0:0] v_2796;
  wire [0:0] v_2797;
  function [0:0] mux_2797(input [0:0] sel);
    case (sel) 0: mux_2797 = 1'h0; 1: mux_2797 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2798;
  wire [0:0] vin0_consume_en_2799;
  wire [0:0] vout_canPeek_2799;
  wire [7:0] vout_peek_2799;
  wire [0:0] v_2800;
  wire [0:0] v_2801;
  function [0:0] mux_2801(input [0:0] sel);
    case (sel) 0: mux_2801 = 1'h0; 1: mux_2801 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2802;
  function [0:0] mux_2802(input [0:0] sel);
    case (sel) 0: mux_2802 = 1'h0; 1: mux_2802 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2803;
  wire [0:0] v_2804;
  wire [0:0] v_2805;
  wire [0:0] v_2806;
  wire [0:0] v_2807;
  wire [0:0] v_2808;
  wire [0:0] v_2809;
  function [0:0] mux_2809(input [0:0] sel);
    case (sel) 0: mux_2809 = 1'h0; 1: mux_2809 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2810;
  function [0:0] mux_2810(input [0:0] sel);
    case (sel) 0: mux_2810 = 1'h0; 1: mux_2810 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2811;
  wire [0:0] v_2812;
  wire [0:0] v_2813;
  wire [0:0] v_2814;
  function [0:0] mux_2814(input [0:0] sel);
    case (sel) 0: mux_2814 = 1'h0; 1: mux_2814 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2815;
  function [0:0] mux_2815(input [0:0] sel);
    case (sel) 0: mux_2815 = 1'h0; 1: mux_2815 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2816;
  wire [0:0] v_2817;
  wire [0:0] v_2818;
  wire [0:0] v_2819;
  wire [0:0] v_2820;
  wire [0:0] v_2821;
  function [0:0] mux_2821(input [0:0] sel);
    case (sel) 0: mux_2821 = 1'h0; 1: mux_2821 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2822;
  function [0:0] mux_2822(input [0:0] sel);
    case (sel) 0: mux_2822 = 1'h0; 1: mux_2822 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2823;
  wire [0:0] v_2824;
  wire [0:0] v_2825;
  wire [0:0] v_2826;
  function [0:0] mux_2826(input [0:0] sel);
    case (sel) 0: mux_2826 = 1'h0; 1: mux_2826 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2827;
  function [0:0] mux_2827(input [0:0] sel);
    case (sel) 0: mux_2827 = 1'h0; 1: mux_2827 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2828;
  wire [0:0] v_2829;
  wire [0:0] v_2830;
  wire [0:0] v_2831;
  wire [0:0] v_2832;
  wire [0:0] v_2833;
  function [0:0] mux_2833(input [0:0] sel);
    case (sel) 0: mux_2833 = 1'h0; 1: mux_2833 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2834;
  wire [0:0] v_2835;
  wire [0:0] v_2836;
  wire [0:0] v_2837;
  wire [0:0] v_2838;
  function [0:0] mux_2838(input [0:0] sel);
    case (sel) 0: mux_2838 = 1'h0; 1: mux_2838 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2839;
  wire [0:0] v_2840;
  wire [0:0] v_2841;
  wire [0:0] v_2842;
  function [0:0] mux_2842(input [0:0] sel);
    case (sel) 0: mux_2842 = 1'h0; 1: mux_2842 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2843;
  function [0:0] mux_2843(input [0:0] sel);
    case (sel) 0: mux_2843 = 1'h0; 1: mux_2843 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2844 = 1'h0;
  wire [0:0] v_2845;
  wire [0:0] v_2846;
  wire [0:0] act_2847;
  wire [0:0] v_2848;
  wire [0:0] v_2849;
  wire [0:0] v_2850;
  reg [0:0] v_2851 = 1'h0;
  wire [0:0] v_2852;
  wire [0:0] v_2853;
  wire [0:0] act_2854;
  wire [0:0] v_2855;
  wire [0:0] v_2856;
  wire [0:0] v_2857;
  reg [0:0] v_2858 = 1'h0;
  wire [0:0] v_2859;
  wire [0:0] v_2860;
  wire [0:0] act_2861;
  wire [0:0] v_2862;
  wire [0:0] v_2863;
  wire [0:0] v_2864;
  wire [0:0] vin0_consume_en_2865;
  wire [0:0] vout_canPeek_2865;
  wire [7:0] vout_peek_2865;
  wire [0:0] v_2866;
  wire [0:0] v_2867;
  function [0:0] mux_2867(input [0:0] sel);
    case (sel) 0: mux_2867 = 1'h0; 1: mux_2867 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2868;
  wire [0:0] v_2869;
  wire [0:0] v_2870;
  wire [0:0] v_2871;
  wire [0:0] v_2872;
  function [0:0] mux_2872(input [0:0] sel);
    case (sel) 0: mux_2872 = 1'h0; 1: mux_2872 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2873;
  wire [0:0] vin0_consume_en_2874;
  wire [0:0] vout_canPeek_2874;
  wire [7:0] vout_peek_2874;
  wire [0:0] v_2875;
  wire [0:0] v_2876;
  function [0:0] mux_2876(input [0:0] sel);
    case (sel) 0: mux_2876 = 1'h0; 1: mux_2876 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2877;
  function [0:0] mux_2877(input [0:0] sel);
    case (sel) 0: mux_2877 = 1'h0; 1: mux_2877 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2878;
  wire [0:0] v_2879;
  wire [0:0] v_2880;
  wire [0:0] v_2881;
  wire [0:0] v_2882;
  wire [0:0] v_2883;
  wire [0:0] v_2884;
  function [0:0] mux_2884(input [0:0] sel);
    case (sel) 0: mux_2884 = 1'h0; 1: mux_2884 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2885;
  wire [0:0] v_2886;
  wire [0:0] v_2887;
  wire [0:0] v_2888;
  wire [0:0] v_2889;
  function [0:0] mux_2889(input [0:0] sel);
    case (sel) 0: mux_2889 = 1'h0; 1: mux_2889 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2890;
  wire [0:0] v_2891;
  wire [0:0] v_2892;
  wire [0:0] v_2893;
  function [0:0] mux_2893(input [0:0] sel);
    case (sel) 0: mux_2893 = 1'h0; 1: mux_2893 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2894;
  function [0:0] mux_2894(input [0:0] sel);
    case (sel) 0: mux_2894 = 1'h0; 1: mux_2894 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2895 = 1'h0;
  wire [0:0] v_2896;
  wire [0:0] v_2897;
  wire [0:0] act_2898;
  wire [0:0] v_2899;
  wire [0:0] v_2900;
  wire [0:0] v_2901;
  wire [0:0] vin0_consume_en_2902;
  wire [0:0] vout_canPeek_2902;
  wire [7:0] vout_peek_2902;
  wire [0:0] v_2903;
  wire [0:0] v_2904;
  function [0:0] mux_2904(input [0:0] sel);
    case (sel) 0: mux_2904 = 1'h0; 1: mux_2904 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2905;
  wire [0:0] v_2906;
  wire [0:0] v_2907;
  wire [0:0] v_2908;
  wire [0:0] v_2909;
  function [0:0] mux_2909(input [0:0] sel);
    case (sel) 0: mux_2909 = 1'h0; 1: mux_2909 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2910;
  wire [0:0] vin0_consume_en_2911;
  wire [0:0] vout_canPeek_2911;
  wire [7:0] vout_peek_2911;
  wire [0:0] v_2912;
  wire [0:0] v_2913;
  function [0:0] mux_2913(input [0:0] sel);
    case (sel) 0: mux_2913 = 1'h0; 1: mux_2913 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2914;
  function [0:0] mux_2914(input [0:0] sel);
    case (sel) 0: mux_2914 = 1'h0; 1: mux_2914 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2915;
  wire [0:0] v_2916;
  wire [0:0] v_2917;
  wire [0:0] v_2918;
  wire [0:0] v_2919;
  wire [0:0] v_2920;
  wire [0:0] v_2921;
  function [0:0] mux_2921(input [0:0] sel);
    case (sel) 0: mux_2921 = 1'h0; 1: mux_2921 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2922;
  function [0:0] mux_2922(input [0:0] sel);
    case (sel) 0: mux_2922 = 1'h0; 1: mux_2922 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2923;
  wire [0:0] v_2924;
  wire [0:0] v_2925;
  wire [0:0] v_2926;
  function [0:0] mux_2926(input [0:0] sel);
    case (sel) 0: mux_2926 = 1'h0; 1: mux_2926 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2927;
  function [0:0] mux_2927(input [0:0] sel);
    case (sel) 0: mux_2927 = 1'h0; 1: mux_2927 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2928;
  wire [0:0] v_2929;
  wire [0:0] v_2930;
  wire [0:0] v_2931;
  wire [0:0] v_2932;
  wire [0:0] v_2933;
  function [0:0] mux_2933(input [0:0] sel);
    case (sel) 0: mux_2933 = 1'h0; 1: mux_2933 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2934;
  wire [0:0] v_2935;
  wire [0:0] v_2936;
  wire [0:0] v_2937;
  wire [0:0] v_2938;
  function [0:0] mux_2938(input [0:0] sel);
    case (sel) 0: mux_2938 = 1'h0; 1: mux_2938 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2939;
  wire [0:0] v_2940;
  wire [0:0] v_2941;
  wire [0:0] v_2942;
  function [0:0] mux_2942(input [0:0] sel);
    case (sel) 0: mux_2942 = 1'h0; 1: mux_2942 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2943;
  function [0:0] mux_2943(input [0:0] sel);
    case (sel) 0: mux_2943 = 1'h0; 1: mux_2943 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2944 = 1'h0;
  wire [0:0] v_2945;
  wire [0:0] v_2946;
  wire [0:0] act_2947;
  wire [0:0] v_2948;
  wire [0:0] v_2949;
  wire [0:0] v_2950;
  reg [0:0] v_2951 = 1'h0;
  wire [0:0] v_2952;
  wire [0:0] v_2953;
  wire [0:0] act_2954;
  wire [0:0] v_2955;
  wire [0:0] v_2956;
  wire [0:0] v_2957;
  wire [0:0] vin0_consume_en_2958;
  wire [0:0] vout_canPeek_2958;
  wire [7:0] vout_peek_2958;
  wire [0:0] v_2959;
  wire [0:0] v_2960;
  function [0:0] mux_2960(input [0:0] sel);
    case (sel) 0: mux_2960 = 1'h0; 1: mux_2960 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2961;
  wire [0:0] v_2962;
  wire [0:0] v_2963;
  wire [0:0] v_2964;
  wire [0:0] v_2965;
  function [0:0] mux_2965(input [0:0] sel);
    case (sel) 0: mux_2965 = 1'h0; 1: mux_2965 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2966;
  wire [0:0] vin0_consume_en_2967;
  wire [0:0] vout_canPeek_2967;
  wire [7:0] vout_peek_2967;
  wire [0:0] v_2968;
  wire [0:0] v_2969;
  function [0:0] mux_2969(input [0:0] sel);
    case (sel) 0: mux_2969 = 1'h0; 1: mux_2969 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2970;
  function [0:0] mux_2970(input [0:0] sel);
    case (sel) 0: mux_2970 = 1'h0; 1: mux_2970 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2971;
  wire [0:0] v_2972;
  wire [0:0] v_2973;
  wire [0:0] v_2974;
  wire [0:0] v_2975;
  wire [0:0] v_2976;
  wire [0:0] v_2977;
  function [0:0] mux_2977(input [0:0] sel);
    case (sel) 0: mux_2977 = 1'h0; 1: mux_2977 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2978;
  wire [0:0] v_2979;
  wire [0:0] v_2980;
  wire [0:0] v_2981;
  wire [0:0] v_2982;
  function [0:0] mux_2982(input [0:0] sel);
    case (sel) 0: mux_2982 = 1'h0; 1: mux_2982 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2983;
  wire [0:0] v_2984;
  wire [0:0] v_2985;
  wire [0:0] v_2986;
  function [0:0] mux_2986(input [0:0] sel);
    case (sel) 0: mux_2986 = 1'h0; 1: mux_2986 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2987;
  function [0:0] mux_2987(input [0:0] sel);
    case (sel) 0: mux_2987 = 1'h0; 1: mux_2987 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2988 = 1'h0;
  wire [0:0] v_2989;
  wire [0:0] v_2990;
  wire [0:0] act_2991;
  wire [0:0] v_2992;
  wire [0:0] v_2993;
  wire [0:0] v_2994;
  wire [0:0] vin0_consume_en_2995;
  wire [0:0] vout_canPeek_2995;
  wire [7:0] vout_peek_2995;
  wire [0:0] v_2996;
  wire [0:0] v_2997;
  function [0:0] mux_2997(input [0:0] sel);
    case (sel) 0: mux_2997 = 1'h0; 1: mux_2997 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2998;
  wire [0:0] v_2999;
  wire [0:0] v_3000;
  wire [0:0] v_3001;
  wire [0:0] v_3002;
  function [0:0] mux_3002(input [0:0] sel);
    case (sel) 0: mux_3002 = 1'h0; 1: mux_3002 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3003;
  wire [0:0] vin0_consume_en_3004;
  wire [0:0] vout_canPeek_3004;
  wire [7:0] vout_peek_3004;
  wire [0:0] v_3005;
  wire [0:0] v_3006;
  function [0:0] mux_3006(input [0:0] sel);
    case (sel) 0: mux_3006 = 1'h0; 1: mux_3006 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3007;
  function [0:0] mux_3007(input [0:0] sel);
    case (sel) 0: mux_3007 = 1'h0; 1: mux_3007 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3008;
  wire [0:0] v_3009;
  wire [0:0] v_3010;
  wire [0:0] v_3011;
  wire [0:0] v_3012;
  wire [0:0] v_3013;
  wire [0:0] v_3014;
  function [0:0] mux_3014(input [0:0] sel);
    case (sel) 0: mux_3014 = 1'h0; 1: mux_3014 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3015;
  function [0:0] mux_3015(input [0:0] sel);
    case (sel) 0: mux_3015 = 1'h0; 1: mux_3015 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3016;
  wire [0:0] v_3017;
  wire [0:0] v_3018;
  wire [0:0] v_3019;
  function [0:0] mux_3019(input [0:0] sel);
    case (sel) 0: mux_3019 = 1'h0; 1: mux_3019 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3020;
  function [0:0] mux_3020(input [0:0] sel);
    case (sel) 0: mux_3020 = 1'h0; 1: mux_3020 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3021;
  wire [0:0] v_3022;
  wire [0:0] v_3023;
  wire [0:0] v_3024;
  wire [0:0] v_3025;
  wire [0:0] v_3026;
  function [0:0] mux_3026(input [0:0] sel);
    case (sel) 0: mux_3026 = 1'h0; 1: mux_3026 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3027;
  function [0:0] mux_3027(input [0:0] sel);
    case (sel) 0: mux_3027 = 1'h0; 1: mux_3027 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3028;
  wire [0:0] v_3029;
  wire [0:0] v_3030;
  wire [0:0] v_3031;
  function [0:0] mux_3031(input [0:0] sel);
    case (sel) 0: mux_3031 = 1'h0; 1: mux_3031 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3032;
  function [0:0] mux_3032(input [0:0] sel);
    case (sel) 0: mux_3032 = 1'h0; 1: mux_3032 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3033;
  wire [0:0] v_3034;
  wire [0:0] v_3035;
  wire [0:0] v_3036;
  wire [0:0] v_3037;
  wire [0:0] v_3038;
  function [0:0] mux_3038(input [0:0] sel);
    case (sel) 0: mux_3038 = 1'h0; 1: mux_3038 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3039;
  function [0:0] mux_3039(input [0:0] sel);
    case (sel) 0: mux_3039 = 1'h0; 1: mux_3039 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3040;
  wire [0:0] v_3041;
  wire [0:0] v_3042;
  wire [0:0] v_3043;
  function [0:0] mux_3043(input [0:0] sel);
    case (sel) 0: mux_3043 = 1'h0; 1: mux_3043 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3044;
  function [0:0] mux_3044(input [0:0] sel);
    case (sel) 0: mux_3044 = 1'h0; 1: mux_3044 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3045;
  wire [0:0] v_3046;
  wire [0:0] v_3047;
  wire [0:0] v_3048;
  wire [0:0] v_3049;
  wire [0:0] v_3050;
  function [0:0] mux_3050(input [0:0] sel);
    case (sel) 0: mux_3050 = 1'h0; 1: mux_3050 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3051;
  wire [0:0] v_3052;
  wire [0:0] v_3053;
  wire [0:0] v_3054;
  wire [0:0] v_3055;
  function [0:0] mux_3055(input [0:0] sel);
    case (sel) 0: mux_3055 = 1'h0; 1: mux_3055 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3056;
  wire [0:0] v_3057;
  wire [0:0] v_3058;
  wire [0:0] v_3059;
  function [0:0] mux_3059(input [0:0] sel);
    case (sel) 0: mux_3059 = 1'h0; 1: mux_3059 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3060;
  function [0:0] mux_3060(input [0:0] sel);
    case (sel) 0: mux_3060 = 1'h0; 1: mux_3060 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3061 = 1'h0;
  wire [0:0] v_3062;
  wire [0:0] v_3063;
  wire [0:0] act_3064;
  wire [0:0] v_3065;
  wire [0:0] v_3066;
  wire [0:0] v_3067;
  reg [0:0] v_3068 = 1'h0;
  wire [0:0] v_3069;
  wire [0:0] v_3070;
  wire [0:0] act_3071;
  wire [0:0] v_3072;
  wire [0:0] v_3073;
  wire [0:0] v_3074;
  reg [0:0] v_3075 = 1'h0;
  wire [0:0] v_3076;
  wire [0:0] v_3077;
  wire [0:0] act_3078;
  wire [0:0] v_3079;
  wire [0:0] v_3080;
  wire [0:0] v_3081;
  reg [0:0] v_3082 = 1'h0;
  wire [0:0] v_3083;
  wire [0:0] v_3084;
  wire [0:0] act_3085;
  wire [0:0] v_3086;
  wire [0:0] v_3087;
  wire [0:0] v_3088;
  wire [0:0] vin0_consume_en_3089;
  wire [0:0] vout_canPeek_3089;
  wire [7:0] vout_peek_3089;
  wire [0:0] v_3090;
  wire [0:0] v_3091;
  function [0:0] mux_3091(input [0:0] sel);
    case (sel) 0: mux_3091 = 1'h0; 1: mux_3091 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3092;
  wire [0:0] v_3093;
  wire [0:0] v_3094;
  wire [0:0] v_3095;
  wire [0:0] v_3096;
  function [0:0] mux_3096(input [0:0] sel);
    case (sel) 0: mux_3096 = 1'h0; 1: mux_3096 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3097;
  wire [0:0] vin0_consume_en_3098;
  wire [0:0] vout_canPeek_3098;
  wire [7:0] vout_peek_3098;
  wire [0:0] v_3099;
  wire [0:0] v_3100;
  function [0:0] mux_3100(input [0:0] sel);
    case (sel) 0: mux_3100 = 1'h0; 1: mux_3100 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3101;
  function [0:0] mux_3101(input [0:0] sel);
    case (sel) 0: mux_3101 = 1'h0; 1: mux_3101 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3102;
  wire [0:0] v_3103;
  wire [0:0] v_3104;
  wire [0:0] v_3105;
  wire [0:0] v_3106;
  wire [0:0] v_3107;
  wire [0:0] v_3108;
  function [0:0] mux_3108(input [0:0] sel);
    case (sel) 0: mux_3108 = 1'h0; 1: mux_3108 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3109;
  wire [0:0] v_3110;
  wire [0:0] v_3111;
  wire [0:0] v_3112;
  wire [0:0] v_3113;
  function [0:0] mux_3113(input [0:0] sel);
    case (sel) 0: mux_3113 = 1'h0; 1: mux_3113 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3114;
  wire [0:0] v_3115;
  wire [0:0] v_3116;
  wire [0:0] v_3117;
  function [0:0] mux_3117(input [0:0] sel);
    case (sel) 0: mux_3117 = 1'h0; 1: mux_3117 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3118;
  function [0:0] mux_3118(input [0:0] sel);
    case (sel) 0: mux_3118 = 1'h0; 1: mux_3118 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3119 = 1'h0;
  wire [0:0] v_3120;
  wire [0:0] v_3121;
  wire [0:0] act_3122;
  wire [0:0] v_3123;
  wire [0:0] v_3124;
  wire [0:0] v_3125;
  wire [0:0] vin0_consume_en_3126;
  wire [0:0] vout_canPeek_3126;
  wire [7:0] vout_peek_3126;
  wire [0:0] v_3127;
  wire [0:0] v_3128;
  function [0:0] mux_3128(input [0:0] sel);
    case (sel) 0: mux_3128 = 1'h0; 1: mux_3128 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3129;
  wire [0:0] v_3130;
  wire [0:0] v_3131;
  wire [0:0] v_3132;
  wire [0:0] v_3133;
  function [0:0] mux_3133(input [0:0] sel);
    case (sel) 0: mux_3133 = 1'h0; 1: mux_3133 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3134;
  wire [0:0] vin0_consume_en_3135;
  wire [0:0] vout_canPeek_3135;
  wire [7:0] vout_peek_3135;
  wire [0:0] v_3136;
  wire [0:0] v_3137;
  function [0:0] mux_3137(input [0:0] sel);
    case (sel) 0: mux_3137 = 1'h0; 1: mux_3137 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3138;
  function [0:0] mux_3138(input [0:0] sel);
    case (sel) 0: mux_3138 = 1'h0; 1: mux_3138 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3139;
  wire [0:0] v_3140;
  wire [0:0] v_3141;
  wire [0:0] v_3142;
  wire [0:0] v_3143;
  wire [0:0] v_3144;
  wire [0:0] v_3145;
  function [0:0] mux_3145(input [0:0] sel);
    case (sel) 0: mux_3145 = 1'h0; 1: mux_3145 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3146;
  function [0:0] mux_3146(input [0:0] sel);
    case (sel) 0: mux_3146 = 1'h0; 1: mux_3146 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3147;
  wire [0:0] v_3148;
  wire [0:0] v_3149;
  wire [0:0] v_3150;
  function [0:0] mux_3150(input [0:0] sel);
    case (sel) 0: mux_3150 = 1'h0; 1: mux_3150 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3151;
  function [0:0] mux_3151(input [0:0] sel);
    case (sel) 0: mux_3151 = 1'h0; 1: mux_3151 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3152;
  wire [0:0] v_3153;
  wire [0:0] v_3154;
  wire [0:0] v_3155;
  wire [0:0] v_3156;
  wire [0:0] v_3157;
  function [0:0] mux_3157(input [0:0] sel);
    case (sel) 0: mux_3157 = 1'h0; 1: mux_3157 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3158;
  wire [0:0] v_3159;
  wire [0:0] v_3160;
  wire [0:0] v_3161;
  wire [0:0] v_3162;
  function [0:0] mux_3162(input [0:0] sel);
    case (sel) 0: mux_3162 = 1'h0; 1: mux_3162 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3163;
  wire [0:0] v_3164;
  wire [0:0] v_3165;
  wire [0:0] v_3166;
  function [0:0] mux_3166(input [0:0] sel);
    case (sel) 0: mux_3166 = 1'h0; 1: mux_3166 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3167;
  function [0:0] mux_3167(input [0:0] sel);
    case (sel) 0: mux_3167 = 1'h0; 1: mux_3167 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3168 = 1'h0;
  wire [0:0] v_3169;
  wire [0:0] v_3170;
  wire [0:0] act_3171;
  wire [0:0] v_3172;
  wire [0:0] v_3173;
  wire [0:0] v_3174;
  reg [0:0] v_3175 = 1'h0;
  wire [0:0] v_3176;
  wire [0:0] v_3177;
  wire [0:0] act_3178;
  wire [0:0] v_3179;
  wire [0:0] v_3180;
  wire [0:0] v_3181;
  wire [0:0] vin0_consume_en_3182;
  wire [0:0] vout_canPeek_3182;
  wire [7:0] vout_peek_3182;
  wire [0:0] v_3183;
  wire [0:0] v_3184;
  function [0:0] mux_3184(input [0:0] sel);
    case (sel) 0: mux_3184 = 1'h0; 1: mux_3184 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3185;
  wire [0:0] v_3186;
  wire [0:0] v_3187;
  wire [0:0] v_3188;
  wire [0:0] v_3189;
  function [0:0] mux_3189(input [0:0] sel);
    case (sel) 0: mux_3189 = 1'h0; 1: mux_3189 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3190;
  wire [0:0] vin0_consume_en_3191;
  wire [0:0] vout_canPeek_3191;
  wire [7:0] vout_peek_3191;
  wire [0:0] v_3192;
  wire [0:0] v_3193;
  function [0:0] mux_3193(input [0:0] sel);
    case (sel) 0: mux_3193 = 1'h0; 1: mux_3193 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3194;
  function [0:0] mux_3194(input [0:0] sel);
    case (sel) 0: mux_3194 = 1'h0; 1: mux_3194 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3195;
  wire [0:0] v_3196;
  wire [0:0] v_3197;
  wire [0:0] v_3198;
  wire [0:0] v_3199;
  wire [0:0] v_3200;
  wire [0:0] v_3201;
  function [0:0] mux_3201(input [0:0] sel);
    case (sel) 0: mux_3201 = 1'h0; 1: mux_3201 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3202;
  wire [0:0] v_3203;
  wire [0:0] v_3204;
  wire [0:0] v_3205;
  wire [0:0] v_3206;
  function [0:0] mux_3206(input [0:0] sel);
    case (sel) 0: mux_3206 = 1'h0; 1: mux_3206 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3207;
  wire [0:0] v_3208;
  wire [0:0] v_3209;
  wire [0:0] v_3210;
  function [0:0] mux_3210(input [0:0] sel);
    case (sel) 0: mux_3210 = 1'h0; 1: mux_3210 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3211;
  function [0:0] mux_3211(input [0:0] sel);
    case (sel) 0: mux_3211 = 1'h0; 1: mux_3211 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3212 = 1'h0;
  wire [0:0] v_3213;
  wire [0:0] v_3214;
  wire [0:0] act_3215;
  wire [0:0] v_3216;
  wire [0:0] v_3217;
  wire [0:0] v_3218;
  wire [0:0] vin0_consume_en_3219;
  wire [0:0] vout_canPeek_3219;
  wire [7:0] vout_peek_3219;
  wire [0:0] v_3220;
  wire [0:0] v_3221;
  function [0:0] mux_3221(input [0:0] sel);
    case (sel) 0: mux_3221 = 1'h0; 1: mux_3221 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3222;
  wire [0:0] v_3223;
  wire [0:0] v_3224;
  wire [0:0] v_3225;
  wire [0:0] v_3226;
  function [0:0] mux_3226(input [0:0] sel);
    case (sel) 0: mux_3226 = 1'h0; 1: mux_3226 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3227;
  wire [0:0] vin0_consume_en_3228;
  wire [0:0] vout_canPeek_3228;
  wire [7:0] vout_peek_3228;
  wire [0:0] v_3229;
  wire [0:0] v_3230;
  function [0:0] mux_3230(input [0:0] sel);
    case (sel) 0: mux_3230 = 1'h0; 1: mux_3230 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3231;
  function [0:0] mux_3231(input [0:0] sel);
    case (sel) 0: mux_3231 = 1'h0; 1: mux_3231 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3232;
  wire [0:0] v_3233;
  wire [0:0] v_3234;
  wire [0:0] v_3235;
  wire [0:0] v_3236;
  wire [0:0] v_3237;
  wire [0:0] v_3238;
  function [0:0] mux_3238(input [0:0] sel);
    case (sel) 0: mux_3238 = 1'h0; 1: mux_3238 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3239;
  function [0:0] mux_3239(input [0:0] sel);
    case (sel) 0: mux_3239 = 1'h0; 1: mux_3239 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3240;
  wire [0:0] v_3241;
  wire [0:0] v_3242;
  wire [0:0] v_3243;
  function [0:0] mux_3243(input [0:0] sel);
    case (sel) 0: mux_3243 = 1'h0; 1: mux_3243 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3244;
  function [0:0] mux_3244(input [0:0] sel);
    case (sel) 0: mux_3244 = 1'h0; 1: mux_3244 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3245;
  wire [0:0] v_3246;
  wire [0:0] v_3247;
  wire [0:0] v_3248;
  wire [0:0] v_3249;
  wire [0:0] v_3250;
  function [0:0] mux_3250(input [0:0] sel);
    case (sel) 0: mux_3250 = 1'h0; 1: mux_3250 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3251;
  function [0:0] mux_3251(input [0:0] sel);
    case (sel) 0: mux_3251 = 1'h0; 1: mux_3251 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3252;
  wire [0:0] v_3253;
  wire [0:0] v_3254;
  wire [0:0] v_3255;
  function [0:0] mux_3255(input [0:0] sel);
    case (sel) 0: mux_3255 = 1'h0; 1: mux_3255 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3256;
  function [0:0] mux_3256(input [0:0] sel);
    case (sel) 0: mux_3256 = 1'h0; 1: mux_3256 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3257;
  wire [0:0] v_3258;
  wire [0:0] v_3259;
  wire [0:0] v_3260;
  wire [0:0] v_3261;
  wire [0:0] v_3262;
  function [0:0] mux_3262(input [0:0] sel);
    case (sel) 0: mux_3262 = 1'h0; 1: mux_3262 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3263;
  wire [0:0] v_3264;
  wire [0:0] v_3265;
  wire [0:0] v_3266;
  wire [0:0] v_3267;
  function [0:0] mux_3267(input [0:0] sel);
    case (sel) 0: mux_3267 = 1'h0; 1: mux_3267 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3268;
  wire [0:0] v_3269;
  wire [0:0] v_3270;
  wire [0:0] v_3271;
  function [0:0] mux_3271(input [0:0] sel);
    case (sel) 0: mux_3271 = 1'h0; 1: mux_3271 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3272;
  function [0:0] mux_3272(input [0:0] sel);
    case (sel) 0: mux_3272 = 1'h0; 1: mux_3272 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3273 = 1'h0;
  wire [0:0] v_3274;
  wire [0:0] v_3275;
  wire [0:0] act_3276;
  wire [0:0] v_3277;
  wire [0:0] v_3278;
  wire [0:0] v_3279;
  reg [0:0] v_3280 = 1'h0;
  wire [0:0] v_3281;
  wire [0:0] v_3282;
  wire [0:0] act_3283;
  wire [0:0] v_3284;
  wire [0:0] v_3285;
  wire [0:0] v_3286;
  reg [0:0] v_3287 = 1'h0;
  wire [0:0] v_3288;
  wire [0:0] v_3289;
  wire [0:0] act_3290;
  wire [0:0] v_3291;
  wire [0:0] v_3292;
  wire [0:0] v_3293;
  wire [0:0] vin0_consume_en_3294;
  wire [0:0] vout_canPeek_3294;
  wire [7:0] vout_peek_3294;
  wire [0:0] v_3295;
  wire [0:0] v_3296;
  function [0:0] mux_3296(input [0:0] sel);
    case (sel) 0: mux_3296 = 1'h0; 1: mux_3296 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3297;
  wire [0:0] v_3298;
  wire [0:0] v_3299;
  wire [0:0] v_3300;
  wire [0:0] v_3301;
  function [0:0] mux_3301(input [0:0] sel);
    case (sel) 0: mux_3301 = 1'h0; 1: mux_3301 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3302;
  wire [0:0] vin0_consume_en_3303;
  wire [0:0] vout_canPeek_3303;
  wire [7:0] vout_peek_3303;
  wire [0:0] v_3304;
  wire [0:0] v_3305;
  function [0:0] mux_3305(input [0:0] sel);
    case (sel) 0: mux_3305 = 1'h0; 1: mux_3305 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3306;
  function [0:0] mux_3306(input [0:0] sel);
    case (sel) 0: mux_3306 = 1'h0; 1: mux_3306 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3307;
  wire [0:0] v_3308;
  wire [0:0] v_3309;
  wire [0:0] v_3310;
  wire [0:0] v_3311;
  wire [0:0] v_3312;
  wire [0:0] v_3313;
  function [0:0] mux_3313(input [0:0] sel);
    case (sel) 0: mux_3313 = 1'h0; 1: mux_3313 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3314;
  wire [0:0] v_3315;
  wire [0:0] v_3316;
  wire [0:0] v_3317;
  wire [0:0] v_3318;
  function [0:0] mux_3318(input [0:0] sel);
    case (sel) 0: mux_3318 = 1'h0; 1: mux_3318 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3319;
  wire [0:0] v_3320;
  wire [0:0] v_3321;
  wire [0:0] v_3322;
  function [0:0] mux_3322(input [0:0] sel);
    case (sel) 0: mux_3322 = 1'h0; 1: mux_3322 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3323;
  function [0:0] mux_3323(input [0:0] sel);
    case (sel) 0: mux_3323 = 1'h0; 1: mux_3323 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3324 = 1'h0;
  wire [0:0] v_3325;
  wire [0:0] v_3326;
  wire [0:0] act_3327;
  wire [0:0] v_3328;
  wire [0:0] v_3329;
  wire [0:0] v_3330;
  wire [0:0] vin0_consume_en_3331;
  wire [0:0] vout_canPeek_3331;
  wire [7:0] vout_peek_3331;
  wire [0:0] v_3332;
  wire [0:0] v_3333;
  function [0:0] mux_3333(input [0:0] sel);
    case (sel) 0: mux_3333 = 1'h0; 1: mux_3333 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3334;
  wire [0:0] v_3335;
  wire [0:0] v_3336;
  wire [0:0] v_3337;
  wire [0:0] v_3338;
  function [0:0] mux_3338(input [0:0] sel);
    case (sel) 0: mux_3338 = 1'h0; 1: mux_3338 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3339;
  wire [0:0] vin0_consume_en_3340;
  wire [0:0] vout_canPeek_3340;
  wire [7:0] vout_peek_3340;
  wire [0:0] v_3341;
  wire [0:0] v_3342;
  function [0:0] mux_3342(input [0:0] sel);
    case (sel) 0: mux_3342 = 1'h0; 1: mux_3342 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3343;
  function [0:0] mux_3343(input [0:0] sel);
    case (sel) 0: mux_3343 = 1'h0; 1: mux_3343 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3344;
  wire [0:0] v_3345;
  wire [0:0] v_3346;
  wire [0:0] v_3347;
  wire [0:0] v_3348;
  wire [0:0] v_3349;
  wire [0:0] v_3350;
  function [0:0] mux_3350(input [0:0] sel);
    case (sel) 0: mux_3350 = 1'h0; 1: mux_3350 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3351;
  function [0:0] mux_3351(input [0:0] sel);
    case (sel) 0: mux_3351 = 1'h0; 1: mux_3351 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3352;
  wire [0:0] v_3353;
  wire [0:0] v_3354;
  wire [0:0] v_3355;
  function [0:0] mux_3355(input [0:0] sel);
    case (sel) 0: mux_3355 = 1'h0; 1: mux_3355 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3356;
  function [0:0] mux_3356(input [0:0] sel);
    case (sel) 0: mux_3356 = 1'h0; 1: mux_3356 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3357;
  wire [0:0] v_3358;
  wire [0:0] v_3359;
  wire [0:0] v_3360;
  wire [0:0] v_3361;
  wire [0:0] v_3362;
  function [0:0] mux_3362(input [0:0] sel);
    case (sel) 0: mux_3362 = 1'h0; 1: mux_3362 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3363;
  wire [0:0] v_3364;
  wire [0:0] v_3365;
  wire [0:0] v_3366;
  wire [0:0] v_3367;
  function [0:0] mux_3367(input [0:0] sel);
    case (sel) 0: mux_3367 = 1'h0; 1: mux_3367 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3368;
  wire [0:0] v_3369;
  wire [0:0] v_3370;
  wire [0:0] v_3371;
  function [0:0] mux_3371(input [0:0] sel);
    case (sel) 0: mux_3371 = 1'h0; 1: mux_3371 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3372;
  function [0:0] mux_3372(input [0:0] sel);
    case (sel) 0: mux_3372 = 1'h0; 1: mux_3372 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3373 = 1'h0;
  wire [0:0] v_3374;
  wire [0:0] v_3375;
  wire [0:0] act_3376;
  wire [0:0] v_3377;
  wire [0:0] v_3378;
  wire [0:0] v_3379;
  reg [0:0] v_3380 = 1'h0;
  wire [0:0] v_3381;
  wire [0:0] v_3382;
  wire [0:0] act_3383;
  wire [0:0] v_3384;
  wire [0:0] v_3385;
  wire [0:0] v_3386;
  wire [0:0] vin0_consume_en_3387;
  wire [0:0] vout_canPeek_3387;
  wire [7:0] vout_peek_3387;
  wire [0:0] v_3388;
  wire [0:0] v_3389;
  function [0:0] mux_3389(input [0:0] sel);
    case (sel) 0: mux_3389 = 1'h0; 1: mux_3389 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3390;
  wire [0:0] v_3391;
  wire [0:0] v_3392;
  wire [0:0] v_3393;
  wire [0:0] v_3394;
  function [0:0] mux_3394(input [0:0] sel);
    case (sel) 0: mux_3394 = 1'h0; 1: mux_3394 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3395;
  wire [0:0] vin0_consume_en_3396;
  wire [0:0] vout_canPeek_3396;
  wire [7:0] vout_peek_3396;
  wire [0:0] v_3397;
  wire [0:0] v_3398;
  function [0:0] mux_3398(input [0:0] sel);
    case (sel) 0: mux_3398 = 1'h0; 1: mux_3398 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3399;
  function [0:0] mux_3399(input [0:0] sel);
    case (sel) 0: mux_3399 = 1'h0; 1: mux_3399 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3400;
  wire [0:0] v_3401;
  wire [0:0] v_3402;
  wire [0:0] v_3403;
  wire [0:0] v_3404;
  wire [0:0] v_3405;
  wire [0:0] v_3406;
  function [0:0] mux_3406(input [0:0] sel);
    case (sel) 0: mux_3406 = 1'h0; 1: mux_3406 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3407;
  wire [0:0] v_3408;
  wire [0:0] v_3409;
  wire [0:0] v_3410;
  wire [0:0] v_3411;
  function [0:0] mux_3411(input [0:0] sel);
    case (sel) 0: mux_3411 = 1'h0; 1: mux_3411 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3412;
  wire [0:0] v_3413;
  wire [0:0] v_3414;
  wire [0:0] v_3415;
  function [0:0] mux_3415(input [0:0] sel);
    case (sel) 0: mux_3415 = 1'h0; 1: mux_3415 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3416;
  function [0:0] mux_3416(input [0:0] sel);
    case (sel) 0: mux_3416 = 1'h0; 1: mux_3416 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3417 = 1'h0;
  wire [0:0] v_3418;
  wire [0:0] v_3419;
  wire [0:0] act_3420;
  wire [0:0] v_3421;
  wire [0:0] v_3422;
  wire [0:0] v_3423;
  wire [0:0] vin0_consume_en_3424;
  wire [0:0] vout_canPeek_3424;
  wire [7:0] vout_peek_3424;
  wire [0:0] v_3425;
  wire [0:0] v_3426;
  function [0:0] mux_3426(input [0:0] sel);
    case (sel) 0: mux_3426 = 1'h0; 1: mux_3426 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3427;
  wire [0:0] v_3428;
  wire [0:0] v_3429;
  wire [0:0] v_3430;
  wire [0:0] v_3431;
  function [0:0] mux_3431(input [0:0] sel);
    case (sel) 0: mux_3431 = 1'h0; 1: mux_3431 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3432;
  wire [0:0] vin0_consume_en_3433;
  wire [0:0] vout_canPeek_3433;
  wire [7:0] vout_peek_3433;
  wire [0:0] v_3434;
  wire [0:0] v_3435;
  function [0:0] mux_3435(input [0:0] sel);
    case (sel) 0: mux_3435 = 1'h0; 1: mux_3435 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3436;
  function [0:0] mux_3436(input [0:0] sel);
    case (sel) 0: mux_3436 = 1'h0; 1: mux_3436 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3437;
  wire [0:0] v_3438;
  wire [0:0] v_3439;
  wire [0:0] v_3440;
  wire [0:0] v_3441;
  wire [0:0] v_3442;
  wire [0:0] v_3443;
  function [0:0] mux_3443(input [0:0] sel);
    case (sel) 0: mux_3443 = 1'h0; 1: mux_3443 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3444;
  function [0:0] mux_3444(input [0:0] sel);
    case (sel) 0: mux_3444 = 1'h0; 1: mux_3444 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3445;
  wire [0:0] v_3446;
  wire [0:0] v_3447;
  wire [0:0] v_3448;
  function [0:0] mux_3448(input [0:0] sel);
    case (sel) 0: mux_3448 = 1'h0; 1: mux_3448 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3449;
  function [0:0] mux_3449(input [0:0] sel);
    case (sel) 0: mux_3449 = 1'h0; 1: mux_3449 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3450;
  wire [0:0] v_3451;
  wire [0:0] v_3452;
  wire [0:0] v_3453;
  wire [0:0] v_3454;
  wire [0:0] v_3455;
  function [0:0] mux_3455(input [0:0] sel);
    case (sel) 0: mux_3455 = 1'h0; 1: mux_3455 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3456;
  function [0:0] mux_3456(input [0:0] sel);
    case (sel) 0: mux_3456 = 1'h0; 1: mux_3456 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3457;
  wire [0:0] v_3458;
  wire [0:0] v_3459;
  wire [0:0] v_3460;
  function [0:0] mux_3460(input [0:0] sel);
    case (sel) 0: mux_3460 = 1'h0; 1: mux_3460 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3461;
  function [0:0] mux_3461(input [0:0] sel);
    case (sel) 0: mux_3461 = 1'h0; 1: mux_3461 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3462;
  wire [0:0] v_3463;
  wire [0:0] v_3464;
  wire [0:0] v_3465;
  wire [0:0] v_3466;
  wire [0:0] v_3467;
  function [0:0] mux_3467(input [0:0] sel);
    case (sel) 0: mux_3467 = 1'h0; 1: mux_3467 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3468;
  function [0:0] mux_3468(input [0:0] sel);
    case (sel) 0: mux_3468 = 1'h0; 1: mux_3468 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3469;
  wire [0:0] v_3470;
  wire [0:0] v_3471;
  wire [0:0] v_3472;
  function [0:0] mux_3472(input [0:0] sel);
    case (sel) 0: mux_3472 = 1'h0; 1: mux_3472 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3473;
  function [0:0] mux_3473(input [0:0] sel);
    case (sel) 0: mux_3473 = 1'h0; 1: mux_3473 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3474;
  wire [0:0] v_3475;
  wire [0:0] v_3476;
  wire [0:0] v_3477;
  wire [0:0] v_3478;
  wire [0:0] v_3479;
  function [0:0] mux_3479(input [0:0] sel);
    case (sel) 0: mux_3479 = 1'h0; 1: mux_3479 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3480;
  function [0:0] mux_3480(input [0:0] sel);
    case (sel) 0: mux_3480 = 1'h0; 1: mux_3480 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3481;
  wire [0:0] v_3482;
  wire [0:0] v_3483;
  wire [0:0] v_3484;
  function [0:0] mux_3484(input [0:0] sel);
    case (sel) 0: mux_3484 = 1'h0; 1: mux_3484 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3485;
  function [0:0] mux_3485(input [0:0] sel);
    case (sel) 0: mux_3485 = 1'h0; 1: mux_3485 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3486;
  wire [0:0] v_3487;
  wire [0:0] v_3488;
  wire [0:0] v_3489;
  wire [0:0] v_3490;
  wire [0:0] v_3491;
  function [0:0] mux_3491(input [0:0] sel);
    case (sel) 0: mux_3491 = 1'h0; 1: mux_3491 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3492;
  wire [0:0] v_3493;
  wire [0:0] v_3494;
  wire [0:0] v_3495;
  wire [0:0] v_3496;
  function [0:0] mux_3496(input [0:0] sel);
    case (sel) 0: mux_3496 = 1'h0; 1: mux_3496 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3497;
  wire [0:0] v_3498;
  wire [0:0] v_3499;
  wire [0:0] v_3500;
  function [0:0] mux_3500(input [0:0] sel);
    case (sel) 0: mux_3500 = 1'h0; 1: mux_3500 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3501;
  function [0:0] mux_3501(input [0:0] sel);
    case (sel) 0: mux_3501 = 1'h0; 1: mux_3501 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3502 = 1'h0;
  wire [0:0] v_3503;
  wire [0:0] v_3504;
  wire [0:0] act_3505;
  wire [0:0] v_3506;
  wire [0:0] v_3507;
  wire [0:0] v_3508;
  reg [0:0] v_3509 = 1'h0;
  wire [0:0] v_3510;
  wire [0:0] v_3511;
  wire [0:0] act_3512;
  wire [0:0] v_3513;
  wire [0:0] v_3514;
  wire [0:0] v_3515;
  reg [0:0] v_3516 = 1'h0;
  wire [0:0] v_3517;
  wire [0:0] v_3518;
  wire [0:0] act_3519;
  wire [0:0] v_3520;
  wire [0:0] v_3521;
  wire [0:0] v_3522;
  reg [0:0] v_3523 = 1'h0;
  wire [0:0] v_3524;
  wire [0:0] v_3525;
  wire [0:0] act_3526;
  wire [0:0] v_3527;
  wire [0:0] v_3528;
  wire [0:0] v_3529;
  reg [0:0] v_3530 = 1'h0;
  wire [0:0] v_3531;
  wire [0:0] v_3532;
  wire [0:0] act_3533;
  wire [0:0] v_3534;
  wire [0:0] v_3535;
  wire [0:0] v_3536;
  wire [0:0] vin0_consume_en_3537;
  wire [0:0] vout_canPeek_3537;
  wire [7:0] vout_peek_3537;
  wire [0:0] v_3538;
  wire [0:0] v_3539;
  function [0:0] mux_3539(input [0:0] sel);
    case (sel) 0: mux_3539 = 1'h0; 1: mux_3539 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3540;
  wire [0:0] v_3541;
  wire [0:0] v_3542;
  wire [0:0] v_3543;
  wire [0:0] v_3544;
  function [0:0] mux_3544(input [0:0] sel);
    case (sel) 0: mux_3544 = 1'h0; 1: mux_3544 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3545;
  wire [0:0] vin0_consume_en_3546;
  wire [0:0] vout_canPeek_3546;
  wire [7:0] vout_peek_3546;
  wire [0:0] v_3547;
  wire [0:0] v_3548;
  function [0:0] mux_3548(input [0:0] sel);
    case (sel) 0: mux_3548 = 1'h0; 1: mux_3548 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3549;
  function [0:0] mux_3549(input [0:0] sel);
    case (sel) 0: mux_3549 = 1'h0; 1: mux_3549 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3550;
  wire [0:0] v_3551;
  wire [0:0] v_3552;
  wire [0:0] v_3553;
  wire [0:0] v_3554;
  wire [0:0] v_3555;
  wire [0:0] v_3556;
  function [0:0] mux_3556(input [0:0] sel);
    case (sel) 0: mux_3556 = 1'h0; 1: mux_3556 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3557;
  wire [0:0] v_3558;
  wire [0:0] v_3559;
  wire [0:0] v_3560;
  wire [0:0] v_3561;
  function [0:0] mux_3561(input [0:0] sel);
    case (sel) 0: mux_3561 = 1'h0; 1: mux_3561 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3562;
  wire [0:0] v_3563;
  wire [0:0] v_3564;
  wire [0:0] v_3565;
  function [0:0] mux_3565(input [0:0] sel);
    case (sel) 0: mux_3565 = 1'h0; 1: mux_3565 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3566;
  function [0:0] mux_3566(input [0:0] sel);
    case (sel) 0: mux_3566 = 1'h0; 1: mux_3566 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3567 = 1'h0;
  wire [0:0] v_3568;
  wire [0:0] v_3569;
  wire [0:0] act_3570;
  wire [0:0] v_3571;
  wire [0:0] v_3572;
  wire [0:0] v_3573;
  wire [0:0] vin0_consume_en_3574;
  wire [0:0] vout_canPeek_3574;
  wire [7:0] vout_peek_3574;
  wire [0:0] v_3575;
  wire [0:0] v_3576;
  function [0:0] mux_3576(input [0:0] sel);
    case (sel) 0: mux_3576 = 1'h0; 1: mux_3576 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3577;
  wire [0:0] v_3578;
  wire [0:0] v_3579;
  wire [0:0] v_3580;
  wire [0:0] v_3581;
  function [0:0] mux_3581(input [0:0] sel);
    case (sel) 0: mux_3581 = 1'h0; 1: mux_3581 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3582;
  wire [0:0] vin0_consume_en_3583;
  wire [0:0] vout_canPeek_3583;
  wire [7:0] vout_peek_3583;
  wire [0:0] v_3584;
  wire [0:0] v_3585;
  function [0:0] mux_3585(input [0:0] sel);
    case (sel) 0: mux_3585 = 1'h0; 1: mux_3585 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3586;
  function [0:0] mux_3586(input [0:0] sel);
    case (sel) 0: mux_3586 = 1'h0; 1: mux_3586 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3587;
  wire [0:0] v_3588;
  wire [0:0] v_3589;
  wire [0:0] v_3590;
  wire [0:0] v_3591;
  wire [0:0] v_3592;
  wire [0:0] v_3593;
  function [0:0] mux_3593(input [0:0] sel);
    case (sel) 0: mux_3593 = 1'h0; 1: mux_3593 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3594;
  function [0:0] mux_3594(input [0:0] sel);
    case (sel) 0: mux_3594 = 1'h0; 1: mux_3594 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3595;
  wire [0:0] v_3596;
  wire [0:0] v_3597;
  wire [0:0] v_3598;
  function [0:0] mux_3598(input [0:0] sel);
    case (sel) 0: mux_3598 = 1'h0; 1: mux_3598 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3599;
  function [0:0] mux_3599(input [0:0] sel);
    case (sel) 0: mux_3599 = 1'h0; 1: mux_3599 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3600;
  wire [0:0] v_3601;
  wire [0:0] v_3602;
  wire [0:0] v_3603;
  wire [0:0] v_3604;
  wire [0:0] v_3605;
  function [0:0] mux_3605(input [0:0] sel);
    case (sel) 0: mux_3605 = 1'h0; 1: mux_3605 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3606;
  wire [0:0] v_3607;
  wire [0:0] v_3608;
  wire [0:0] v_3609;
  wire [0:0] v_3610;
  function [0:0] mux_3610(input [0:0] sel);
    case (sel) 0: mux_3610 = 1'h0; 1: mux_3610 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3611;
  wire [0:0] v_3612;
  wire [0:0] v_3613;
  wire [0:0] v_3614;
  function [0:0] mux_3614(input [0:0] sel);
    case (sel) 0: mux_3614 = 1'h0; 1: mux_3614 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3615;
  function [0:0] mux_3615(input [0:0] sel);
    case (sel) 0: mux_3615 = 1'h0; 1: mux_3615 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3616 = 1'h0;
  wire [0:0] v_3617;
  wire [0:0] v_3618;
  wire [0:0] act_3619;
  wire [0:0] v_3620;
  wire [0:0] v_3621;
  wire [0:0] v_3622;
  reg [0:0] v_3623 = 1'h0;
  wire [0:0] v_3624;
  wire [0:0] v_3625;
  wire [0:0] act_3626;
  wire [0:0] v_3627;
  wire [0:0] v_3628;
  wire [0:0] v_3629;
  wire [0:0] vin0_consume_en_3630;
  wire [0:0] vout_canPeek_3630;
  wire [7:0] vout_peek_3630;
  wire [0:0] v_3631;
  wire [0:0] v_3632;
  function [0:0] mux_3632(input [0:0] sel);
    case (sel) 0: mux_3632 = 1'h0; 1: mux_3632 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3633;
  wire [0:0] v_3634;
  wire [0:0] v_3635;
  wire [0:0] v_3636;
  wire [0:0] v_3637;
  function [0:0] mux_3637(input [0:0] sel);
    case (sel) 0: mux_3637 = 1'h0; 1: mux_3637 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3638;
  wire [0:0] vin0_consume_en_3639;
  wire [0:0] vout_canPeek_3639;
  wire [7:0] vout_peek_3639;
  wire [0:0] v_3640;
  wire [0:0] v_3641;
  function [0:0] mux_3641(input [0:0] sel);
    case (sel) 0: mux_3641 = 1'h0; 1: mux_3641 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3642;
  function [0:0] mux_3642(input [0:0] sel);
    case (sel) 0: mux_3642 = 1'h0; 1: mux_3642 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3643;
  wire [0:0] v_3644;
  wire [0:0] v_3645;
  wire [0:0] v_3646;
  wire [0:0] v_3647;
  wire [0:0] v_3648;
  wire [0:0] v_3649;
  function [0:0] mux_3649(input [0:0] sel);
    case (sel) 0: mux_3649 = 1'h0; 1: mux_3649 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3650;
  wire [0:0] v_3651;
  wire [0:0] v_3652;
  wire [0:0] v_3653;
  wire [0:0] v_3654;
  function [0:0] mux_3654(input [0:0] sel);
    case (sel) 0: mux_3654 = 1'h0; 1: mux_3654 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3655;
  wire [0:0] v_3656;
  wire [0:0] v_3657;
  wire [0:0] v_3658;
  function [0:0] mux_3658(input [0:0] sel);
    case (sel) 0: mux_3658 = 1'h0; 1: mux_3658 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3659;
  function [0:0] mux_3659(input [0:0] sel);
    case (sel) 0: mux_3659 = 1'h0; 1: mux_3659 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3660 = 1'h0;
  wire [0:0] v_3661;
  wire [0:0] v_3662;
  wire [0:0] act_3663;
  wire [0:0] v_3664;
  wire [0:0] v_3665;
  wire [0:0] v_3666;
  wire [0:0] vin0_consume_en_3667;
  wire [0:0] vout_canPeek_3667;
  wire [7:0] vout_peek_3667;
  wire [0:0] v_3668;
  wire [0:0] v_3669;
  function [0:0] mux_3669(input [0:0] sel);
    case (sel) 0: mux_3669 = 1'h0; 1: mux_3669 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3670;
  wire [0:0] v_3671;
  wire [0:0] v_3672;
  wire [0:0] v_3673;
  wire [0:0] v_3674;
  function [0:0] mux_3674(input [0:0] sel);
    case (sel) 0: mux_3674 = 1'h0; 1: mux_3674 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3675;
  wire [0:0] vin0_consume_en_3676;
  wire [0:0] vout_canPeek_3676;
  wire [7:0] vout_peek_3676;
  wire [0:0] v_3677;
  wire [0:0] v_3678;
  function [0:0] mux_3678(input [0:0] sel);
    case (sel) 0: mux_3678 = 1'h0; 1: mux_3678 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3679;
  function [0:0] mux_3679(input [0:0] sel);
    case (sel) 0: mux_3679 = 1'h0; 1: mux_3679 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3680;
  wire [0:0] v_3681;
  wire [0:0] v_3682;
  wire [0:0] v_3683;
  wire [0:0] v_3684;
  wire [0:0] v_3685;
  wire [0:0] v_3686;
  function [0:0] mux_3686(input [0:0] sel);
    case (sel) 0: mux_3686 = 1'h0; 1: mux_3686 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3687;
  function [0:0] mux_3687(input [0:0] sel);
    case (sel) 0: mux_3687 = 1'h0; 1: mux_3687 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3688;
  wire [0:0] v_3689;
  wire [0:0] v_3690;
  wire [0:0] v_3691;
  function [0:0] mux_3691(input [0:0] sel);
    case (sel) 0: mux_3691 = 1'h0; 1: mux_3691 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3692;
  function [0:0] mux_3692(input [0:0] sel);
    case (sel) 0: mux_3692 = 1'h0; 1: mux_3692 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3693;
  wire [0:0] v_3694;
  wire [0:0] v_3695;
  wire [0:0] v_3696;
  wire [0:0] v_3697;
  wire [0:0] v_3698;
  function [0:0] mux_3698(input [0:0] sel);
    case (sel) 0: mux_3698 = 1'h0; 1: mux_3698 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3699;
  function [0:0] mux_3699(input [0:0] sel);
    case (sel) 0: mux_3699 = 1'h0; 1: mux_3699 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3700;
  wire [0:0] v_3701;
  wire [0:0] v_3702;
  wire [0:0] v_3703;
  function [0:0] mux_3703(input [0:0] sel);
    case (sel) 0: mux_3703 = 1'h0; 1: mux_3703 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3704;
  function [0:0] mux_3704(input [0:0] sel);
    case (sel) 0: mux_3704 = 1'h0; 1: mux_3704 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3705;
  wire [0:0] v_3706;
  wire [0:0] v_3707;
  wire [0:0] v_3708;
  wire [0:0] v_3709;
  wire [0:0] v_3710;
  function [0:0] mux_3710(input [0:0] sel);
    case (sel) 0: mux_3710 = 1'h0; 1: mux_3710 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3711;
  wire [0:0] v_3712;
  wire [0:0] v_3713;
  wire [0:0] v_3714;
  wire [0:0] v_3715;
  function [0:0] mux_3715(input [0:0] sel);
    case (sel) 0: mux_3715 = 1'h0; 1: mux_3715 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3716;
  wire [0:0] v_3717;
  wire [0:0] v_3718;
  wire [0:0] v_3719;
  function [0:0] mux_3719(input [0:0] sel);
    case (sel) 0: mux_3719 = 1'h0; 1: mux_3719 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3720;
  function [0:0] mux_3720(input [0:0] sel);
    case (sel) 0: mux_3720 = 1'h0; 1: mux_3720 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3721 = 1'h0;
  wire [0:0] v_3722;
  wire [0:0] v_3723;
  wire [0:0] act_3724;
  wire [0:0] v_3725;
  wire [0:0] v_3726;
  wire [0:0] v_3727;
  reg [0:0] v_3728 = 1'h0;
  wire [0:0] v_3729;
  wire [0:0] v_3730;
  wire [0:0] act_3731;
  wire [0:0] v_3732;
  wire [0:0] v_3733;
  wire [0:0] v_3734;
  reg [0:0] v_3735 = 1'h0;
  wire [0:0] v_3736;
  wire [0:0] v_3737;
  wire [0:0] act_3738;
  wire [0:0] v_3739;
  wire [0:0] v_3740;
  wire [0:0] v_3741;
  wire [0:0] vin0_consume_en_3742;
  wire [0:0] vout_canPeek_3742;
  wire [7:0] vout_peek_3742;
  wire [0:0] v_3743;
  wire [0:0] v_3744;
  function [0:0] mux_3744(input [0:0] sel);
    case (sel) 0: mux_3744 = 1'h0; 1: mux_3744 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3745;
  wire [0:0] v_3746;
  wire [0:0] v_3747;
  wire [0:0] v_3748;
  wire [0:0] v_3749;
  function [0:0] mux_3749(input [0:0] sel);
    case (sel) 0: mux_3749 = 1'h0; 1: mux_3749 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3750;
  wire [0:0] vin0_consume_en_3751;
  wire [0:0] vout_canPeek_3751;
  wire [7:0] vout_peek_3751;
  wire [0:0] v_3752;
  wire [0:0] v_3753;
  function [0:0] mux_3753(input [0:0] sel);
    case (sel) 0: mux_3753 = 1'h0; 1: mux_3753 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3754;
  function [0:0] mux_3754(input [0:0] sel);
    case (sel) 0: mux_3754 = 1'h0; 1: mux_3754 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3755;
  wire [0:0] v_3756;
  wire [0:0] v_3757;
  wire [0:0] v_3758;
  wire [0:0] v_3759;
  wire [0:0] v_3760;
  wire [0:0] v_3761;
  function [0:0] mux_3761(input [0:0] sel);
    case (sel) 0: mux_3761 = 1'h0; 1: mux_3761 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3762;
  wire [0:0] v_3763;
  wire [0:0] v_3764;
  wire [0:0] v_3765;
  wire [0:0] v_3766;
  function [0:0] mux_3766(input [0:0] sel);
    case (sel) 0: mux_3766 = 1'h0; 1: mux_3766 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3767;
  wire [0:0] v_3768;
  wire [0:0] v_3769;
  wire [0:0] v_3770;
  function [0:0] mux_3770(input [0:0] sel);
    case (sel) 0: mux_3770 = 1'h0; 1: mux_3770 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3771;
  function [0:0] mux_3771(input [0:0] sel);
    case (sel) 0: mux_3771 = 1'h0; 1: mux_3771 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3772 = 1'h0;
  wire [0:0] v_3773;
  wire [0:0] v_3774;
  wire [0:0] act_3775;
  wire [0:0] v_3776;
  wire [0:0] v_3777;
  wire [0:0] v_3778;
  wire [0:0] vin0_consume_en_3779;
  wire [0:0] vout_canPeek_3779;
  wire [7:0] vout_peek_3779;
  wire [0:0] v_3780;
  wire [0:0] v_3781;
  function [0:0] mux_3781(input [0:0] sel);
    case (sel) 0: mux_3781 = 1'h0; 1: mux_3781 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3782;
  wire [0:0] v_3783;
  wire [0:0] v_3784;
  wire [0:0] v_3785;
  wire [0:0] v_3786;
  function [0:0] mux_3786(input [0:0] sel);
    case (sel) 0: mux_3786 = 1'h0; 1: mux_3786 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3787;
  wire [0:0] vin0_consume_en_3788;
  wire [0:0] vout_canPeek_3788;
  wire [7:0] vout_peek_3788;
  wire [0:0] v_3789;
  wire [0:0] v_3790;
  function [0:0] mux_3790(input [0:0] sel);
    case (sel) 0: mux_3790 = 1'h0; 1: mux_3790 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3791;
  function [0:0] mux_3791(input [0:0] sel);
    case (sel) 0: mux_3791 = 1'h0; 1: mux_3791 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3792;
  wire [0:0] v_3793;
  wire [0:0] v_3794;
  wire [0:0] v_3795;
  wire [0:0] v_3796;
  wire [0:0] v_3797;
  wire [0:0] v_3798;
  function [0:0] mux_3798(input [0:0] sel);
    case (sel) 0: mux_3798 = 1'h0; 1: mux_3798 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3799;
  function [0:0] mux_3799(input [0:0] sel);
    case (sel) 0: mux_3799 = 1'h0; 1: mux_3799 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3800;
  wire [0:0] v_3801;
  wire [0:0] v_3802;
  wire [0:0] v_3803;
  function [0:0] mux_3803(input [0:0] sel);
    case (sel) 0: mux_3803 = 1'h0; 1: mux_3803 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3804;
  function [0:0] mux_3804(input [0:0] sel);
    case (sel) 0: mux_3804 = 1'h0; 1: mux_3804 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3805;
  wire [0:0] v_3806;
  wire [0:0] v_3807;
  wire [0:0] v_3808;
  wire [0:0] v_3809;
  wire [0:0] v_3810;
  function [0:0] mux_3810(input [0:0] sel);
    case (sel) 0: mux_3810 = 1'h0; 1: mux_3810 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3811;
  wire [0:0] v_3812;
  wire [0:0] v_3813;
  wire [0:0] v_3814;
  wire [0:0] v_3815;
  function [0:0] mux_3815(input [0:0] sel);
    case (sel) 0: mux_3815 = 1'h0; 1: mux_3815 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3816;
  wire [0:0] v_3817;
  wire [0:0] v_3818;
  wire [0:0] v_3819;
  function [0:0] mux_3819(input [0:0] sel);
    case (sel) 0: mux_3819 = 1'h0; 1: mux_3819 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3820;
  function [0:0] mux_3820(input [0:0] sel);
    case (sel) 0: mux_3820 = 1'h0; 1: mux_3820 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3821 = 1'h0;
  wire [0:0] v_3822;
  wire [0:0] v_3823;
  wire [0:0] act_3824;
  wire [0:0] v_3825;
  wire [0:0] v_3826;
  wire [0:0] v_3827;
  reg [0:0] v_3828 = 1'h0;
  wire [0:0] v_3829;
  wire [0:0] v_3830;
  wire [0:0] act_3831;
  wire [0:0] v_3832;
  wire [0:0] v_3833;
  wire [0:0] v_3834;
  wire [0:0] vin0_consume_en_3835;
  wire [0:0] vout_canPeek_3835;
  wire [7:0] vout_peek_3835;
  wire [0:0] v_3836;
  wire [0:0] v_3837;
  function [0:0] mux_3837(input [0:0] sel);
    case (sel) 0: mux_3837 = 1'h0; 1: mux_3837 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3838;
  wire [0:0] v_3839;
  wire [0:0] v_3840;
  wire [0:0] v_3841;
  wire [0:0] v_3842;
  function [0:0] mux_3842(input [0:0] sel);
    case (sel) 0: mux_3842 = 1'h0; 1: mux_3842 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3843;
  wire [0:0] vin0_consume_en_3844;
  wire [0:0] vout_canPeek_3844;
  wire [7:0] vout_peek_3844;
  wire [0:0] v_3845;
  wire [0:0] v_3846;
  function [0:0] mux_3846(input [0:0] sel);
    case (sel) 0: mux_3846 = 1'h0; 1: mux_3846 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3847;
  function [0:0] mux_3847(input [0:0] sel);
    case (sel) 0: mux_3847 = 1'h0; 1: mux_3847 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3848;
  wire [0:0] v_3849;
  wire [0:0] v_3850;
  wire [0:0] v_3851;
  wire [0:0] v_3852;
  wire [0:0] v_3853;
  wire [0:0] v_3854;
  function [0:0] mux_3854(input [0:0] sel);
    case (sel) 0: mux_3854 = 1'h0; 1: mux_3854 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3855;
  wire [0:0] v_3856;
  wire [0:0] v_3857;
  wire [0:0] v_3858;
  wire [0:0] v_3859;
  function [0:0] mux_3859(input [0:0] sel);
    case (sel) 0: mux_3859 = 1'h0; 1: mux_3859 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3860;
  wire [0:0] v_3861;
  wire [0:0] v_3862;
  wire [0:0] v_3863;
  function [0:0] mux_3863(input [0:0] sel);
    case (sel) 0: mux_3863 = 1'h0; 1: mux_3863 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3864;
  function [0:0] mux_3864(input [0:0] sel);
    case (sel) 0: mux_3864 = 1'h0; 1: mux_3864 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3865 = 1'h0;
  wire [0:0] v_3866;
  wire [0:0] v_3867;
  wire [0:0] act_3868;
  wire [0:0] v_3869;
  wire [0:0] v_3870;
  wire [0:0] v_3871;
  wire [0:0] vin0_consume_en_3872;
  wire [0:0] vout_canPeek_3872;
  wire [7:0] vout_peek_3872;
  wire [0:0] v_3873;
  wire [0:0] v_3874;
  function [0:0] mux_3874(input [0:0] sel);
    case (sel) 0: mux_3874 = 1'h0; 1: mux_3874 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3875;
  wire [0:0] v_3876;
  wire [0:0] v_3877;
  wire [0:0] v_3878;
  wire [0:0] v_3879;
  function [0:0] mux_3879(input [0:0] sel);
    case (sel) 0: mux_3879 = 1'h0; 1: mux_3879 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3880;
  wire [0:0] vin0_consume_en_3881;
  wire [0:0] vout_canPeek_3881;
  wire [7:0] vout_peek_3881;
  wire [0:0] v_3882;
  wire [0:0] v_3883;
  function [0:0] mux_3883(input [0:0] sel);
    case (sel) 0: mux_3883 = 1'h0; 1: mux_3883 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3884;
  function [0:0] mux_3884(input [0:0] sel);
    case (sel) 0: mux_3884 = 1'h0; 1: mux_3884 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3885;
  wire [0:0] v_3886;
  wire [0:0] v_3887;
  wire [0:0] v_3888;
  wire [0:0] v_3889;
  wire [0:0] v_3890;
  wire [0:0] v_3891;
  function [0:0] mux_3891(input [0:0] sel);
    case (sel) 0: mux_3891 = 1'h0; 1: mux_3891 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3892;
  function [0:0] mux_3892(input [0:0] sel);
    case (sel) 0: mux_3892 = 1'h0; 1: mux_3892 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3893;
  wire [0:0] v_3894;
  wire [0:0] v_3895;
  wire [0:0] v_3896;
  function [0:0] mux_3896(input [0:0] sel);
    case (sel) 0: mux_3896 = 1'h0; 1: mux_3896 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3897;
  function [0:0] mux_3897(input [0:0] sel);
    case (sel) 0: mux_3897 = 1'h0; 1: mux_3897 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3898;
  wire [0:0] v_3899;
  wire [0:0] v_3900;
  wire [0:0] v_3901;
  wire [0:0] v_3902;
  wire [0:0] v_3903;
  function [0:0] mux_3903(input [0:0] sel);
    case (sel) 0: mux_3903 = 1'h0; 1: mux_3903 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3904;
  function [0:0] mux_3904(input [0:0] sel);
    case (sel) 0: mux_3904 = 1'h0; 1: mux_3904 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3905;
  wire [0:0] v_3906;
  wire [0:0] v_3907;
  wire [0:0] v_3908;
  function [0:0] mux_3908(input [0:0] sel);
    case (sel) 0: mux_3908 = 1'h0; 1: mux_3908 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3909;
  function [0:0] mux_3909(input [0:0] sel);
    case (sel) 0: mux_3909 = 1'h0; 1: mux_3909 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3910;
  wire [0:0] v_3911;
  wire [0:0] v_3912;
  wire [0:0] v_3913;
  wire [0:0] v_3914;
  wire [0:0] v_3915;
  function [0:0] mux_3915(input [0:0] sel);
    case (sel) 0: mux_3915 = 1'h0; 1: mux_3915 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3916;
  function [0:0] mux_3916(input [0:0] sel);
    case (sel) 0: mux_3916 = 1'h0; 1: mux_3916 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3917;
  wire [0:0] v_3918;
  wire [0:0] v_3919;
  wire [0:0] v_3920;
  function [0:0] mux_3920(input [0:0] sel);
    case (sel) 0: mux_3920 = 1'h0; 1: mux_3920 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3921;
  function [0:0] mux_3921(input [0:0] sel);
    case (sel) 0: mux_3921 = 1'h0; 1: mux_3921 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3922;
  wire [0:0] v_3923;
  wire [0:0] v_3924;
  wire [0:0] v_3925;
  wire [0:0] v_3926;
  wire [0:0] v_3927;
  function [0:0] mux_3927(input [0:0] sel);
    case (sel) 0: mux_3927 = 1'h0; 1: mux_3927 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3928;
  wire [0:0] v_3929;
  wire [0:0] v_3930;
  wire [0:0] v_3931;
  wire [0:0] v_3932;
  function [0:0] mux_3932(input [0:0] sel);
    case (sel) 0: mux_3932 = 1'h0; 1: mux_3932 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3933;
  wire [0:0] v_3934;
  wire [0:0] v_3935;
  wire [0:0] v_3936;
  function [0:0] mux_3936(input [0:0] sel);
    case (sel) 0: mux_3936 = 1'h0; 1: mux_3936 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3937;
  function [0:0] mux_3937(input [0:0] sel);
    case (sel) 0: mux_3937 = 1'h0; 1: mux_3937 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3938 = 1'h0;
  wire [0:0] v_3939;
  wire [0:0] v_3940;
  wire [0:0] act_3941;
  wire [0:0] v_3942;
  wire [0:0] v_3943;
  wire [0:0] v_3944;
  reg [0:0] v_3945 = 1'h0;
  wire [0:0] v_3946;
  wire [0:0] v_3947;
  wire [0:0] act_3948;
  wire [0:0] v_3949;
  wire [0:0] v_3950;
  wire [0:0] v_3951;
  reg [0:0] v_3952 = 1'h0;
  wire [0:0] v_3953;
  wire [0:0] v_3954;
  wire [0:0] act_3955;
  wire [0:0] v_3956;
  wire [0:0] v_3957;
  wire [0:0] v_3958;
  reg [0:0] v_3959 = 1'h0;
  wire [0:0] v_3960;
  wire [0:0] v_3961;
  wire [0:0] act_3962;
  wire [0:0] v_3963;
  wire [0:0] v_3964;
  wire [0:0] v_3965;
  wire [0:0] vin0_consume_en_3966;
  wire [0:0] vout_canPeek_3966;
  wire [7:0] vout_peek_3966;
  wire [0:0] v_3967;
  wire [0:0] v_3968;
  function [0:0] mux_3968(input [0:0] sel);
    case (sel) 0: mux_3968 = 1'h0; 1: mux_3968 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3969;
  wire [0:0] v_3970;
  wire [0:0] v_3971;
  wire [0:0] v_3972;
  wire [0:0] v_3973;
  function [0:0] mux_3973(input [0:0] sel);
    case (sel) 0: mux_3973 = 1'h0; 1: mux_3973 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3974;
  wire [0:0] vin0_consume_en_3975;
  wire [0:0] vout_canPeek_3975;
  wire [7:0] vout_peek_3975;
  wire [0:0] v_3976;
  wire [0:0] v_3977;
  function [0:0] mux_3977(input [0:0] sel);
    case (sel) 0: mux_3977 = 1'h0; 1: mux_3977 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3978;
  function [0:0] mux_3978(input [0:0] sel);
    case (sel) 0: mux_3978 = 1'h0; 1: mux_3978 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3979;
  wire [0:0] v_3980;
  wire [0:0] v_3981;
  wire [0:0] v_3982;
  wire [0:0] v_3983;
  wire [0:0] v_3984;
  wire [0:0] v_3985;
  function [0:0] mux_3985(input [0:0] sel);
    case (sel) 0: mux_3985 = 1'h0; 1: mux_3985 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3986;
  wire [0:0] v_3987;
  wire [0:0] v_3988;
  wire [0:0] v_3989;
  wire [0:0] v_3990;
  function [0:0] mux_3990(input [0:0] sel);
    case (sel) 0: mux_3990 = 1'h0; 1: mux_3990 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3991;
  wire [0:0] v_3992;
  wire [0:0] v_3993;
  wire [0:0] v_3994;
  function [0:0] mux_3994(input [0:0] sel);
    case (sel) 0: mux_3994 = 1'h0; 1: mux_3994 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3995;
  function [0:0] mux_3995(input [0:0] sel);
    case (sel) 0: mux_3995 = 1'h0; 1: mux_3995 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3996 = 1'h0;
  wire [0:0] v_3997;
  wire [0:0] v_3998;
  wire [0:0] act_3999;
  wire [0:0] v_4000;
  wire [0:0] v_4001;
  wire [0:0] v_4002;
  wire [0:0] vin0_consume_en_4003;
  wire [0:0] vout_canPeek_4003;
  wire [7:0] vout_peek_4003;
  wire [0:0] v_4004;
  wire [0:0] v_4005;
  function [0:0] mux_4005(input [0:0] sel);
    case (sel) 0: mux_4005 = 1'h0; 1: mux_4005 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4006;
  wire [0:0] v_4007;
  wire [0:0] v_4008;
  wire [0:0] v_4009;
  wire [0:0] v_4010;
  function [0:0] mux_4010(input [0:0] sel);
    case (sel) 0: mux_4010 = 1'h0; 1: mux_4010 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4011;
  wire [0:0] vin0_consume_en_4012;
  wire [0:0] vout_canPeek_4012;
  wire [7:0] vout_peek_4012;
  wire [0:0] v_4013;
  wire [0:0] v_4014;
  function [0:0] mux_4014(input [0:0] sel);
    case (sel) 0: mux_4014 = 1'h0; 1: mux_4014 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4015;
  function [0:0] mux_4015(input [0:0] sel);
    case (sel) 0: mux_4015 = 1'h0; 1: mux_4015 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4016;
  wire [0:0] v_4017;
  wire [0:0] v_4018;
  wire [0:0] v_4019;
  wire [0:0] v_4020;
  wire [0:0] v_4021;
  wire [0:0] v_4022;
  function [0:0] mux_4022(input [0:0] sel);
    case (sel) 0: mux_4022 = 1'h0; 1: mux_4022 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4023;
  function [0:0] mux_4023(input [0:0] sel);
    case (sel) 0: mux_4023 = 1'h0; 1: mux_4023 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4024;
  wire [0:0] v_4025;
  wire [0:0] v_4026;
  wire [0:0] v_4027;
  function [0:0] mux_4027(input [0:0] sel);
    case (sel) 0: mux_4027 = 1'h0; 1: mux_4027 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4028;
  function [0:0] mux_4028(input [0:0] sel);
    case (sel) 0: mux_4028 = 1'h0; 1: mux_4028 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4029;
  wire [0:0] v_4030;
  wire [0:0] v_4031;
  wire [0:0] v_4032;
  wire [0:0] v_4033;
  wire [0:0] v_4034;
  function [0:0] mux_4034(input [0:0] sel);
    case (sel) 0: mux_4034 = 1'h0; 1: mux_4034 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4035;
  wire [0:0] v_4036;
  wire [0:0] v_4037;
  wire [0:0] v_4038;
  wire [0:0] v_4039;
  function [0:0] mux_4039(input [0:0] sel);
    case (sel) 0: mux_4039 = 1'h0; 1: mux_4039 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4040;
  wire [0:0] v_4041;
  wire [0:0] v_4042;
  wire [0:0] v_4043;
  function [0:0] mux_4043(input [0:0] sel);
    case (sel) 0: mux_4043 = 1'h0; 1: mux_4043 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4044;
  function [0:0] mux_4044(input [0:0] sel);
    case (sel) 0: mux_4044 = 1'h0; 1: mux_4044 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4045 = 1'h0;
  wire [0:0] v_4046;
  wire [0:0] v_4047;
  wire [0:0] act_4048;
  wire [0:0] v_4049;
  wire [0:0] v_4050;
  wire [0:0] v_4051;
  reg [0:0] v_4052 = 1'h0;
  wire [0:0] v_4053;
  wire [0:0] v_4054;
  wire [0:0] act_4055;
  wire [0:0] v_4056;
  wire [0:0] v_4057;
  wire [0:0] v_4058;
  wire [0:0] vin0_consume_en_4059;
  wire [0:0] vout_canPeek_4059;
  wire [7:0] vout_peek_4059;
  wire [0:0] v_4060;
  wire [0:0] v_4061;
  function [0:0] mux_4061(input [0:0] sel);
    case (sel) 0: mux_4061 = 1'h0; 1: mux_4061 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4062;
  wire [0:0] v_4063;
  wire [0:0] v_4064;
  wire [0:0] v_4065;
  wire [0:0] v_4066;
  function [0:0] mux_4066(input [0:0] sel);
    case (sel) 0: mux_4066 = 1'h0; 1: mux_4066 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4067;
  wire [0:0] vin0_consume_en_4068;
  wire [0:0] vout_canPeek_4068;
  wire [7:0] vout_peek_4068;
  wire [0:0] v_4069;
  wire [0:0] v_4070;
  function [0:0] mux_4070(input [0:0] sel);
    case (sel) 0: mux_4070 = 1'h0; 1: mux_4070 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4071;
  function [0:0] mux_4071(input [0:0] sel);
    case (sel) 0: mux_4071 = 1'h0; 1: mux_4071 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4072;
  wire [0:0] v_4073;
  wire [0:0] v_4074;
  wire [0:0] v_4075;
  wire [0:0] v_4076;
  wire [0:0] v_4077;
  wire [0:0] v_4078;
  function [0:0] mux_4078(input [0:0] sel);
    case (sel) 0: mux_4078 = 1'h0; 1: mux_4078 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4079;
  wire [0:0] v_4080;
  wire [0:0] v_4081;
  wire [0:0] v_4082;
  wire [0:0] v_4083;
  function [0:0] mux_4083(input [0:0] sel);
    case (sel) 0: mux_4083 = 1'h0; 1: mux_4083 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4084;
  wire [0:0] v_4085;
  wire [0:0] v_4086;
  wire [0:0] v_4087;
  function [0:0] mux_4087(input [0:0] sel);
    case (sel) 0: mux_4087 = 1'h0; 1: mux_4087 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4088;
  function [0:0] mux_4088(input [0:0] sel);
    case (sel) 0: mux_4088 = 1'h0; 1: mux_4088 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4089 = 1'h0;
  wire [0:0] v_4090;
  wire [0:0] v_4091;
  wire [0:0] act_4092;
  wire [0:0] v_4093;
  wire [0:0] v_4094;
  wire [0:0] v_4095;
  wire [0:0] vin0_consume_en_4096;
  wire [0:0] vout_canPeek_4096;
  wire [7:0] vout_peek_4096;
  wire [0:0] v_4097;
  wire [0:0] v_4098;
  function [0:0] mux_4098(input [0:0] sel);
    case (sel) 0: mux_4098 = 1'h0; 1: mux_4098 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4099;
  wire [0:0] v_4100;
  wire [0:0] v_4101;
  wire [0:0] v_4102;
  wire [0:0] v_4103;
  function [0:0] mux_4103(input [0:0] sel);
    case (sel) 0: mux_4103 = 1'h0; 1: mux_4103 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4104;
  wire [0:0] vin0_consume_en_4105;
  wire [0:0] vout_canPeek_4105;
  wire [7:0] vout_peek_4105;
  wire [0:0] v_4106;
  wire [0:0] v_4107;
  function [0:0] mux_4107(input [0:0] sel);
    case (sel) 0: mux_4107 = 1'h0; 1: mux_4107 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4108;
  function [0:0] mux_4108(input [0:0] sel);
    case (sel) 0: mux_4108 = 1'h0; 1: mux_4108 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4109;
  wire [0:0] v_4110;
  wire [0:0] v_4111;
  wire [0:0] v_4112;
  wire [0:0] v_4113;
  wire [0:0] v_4114;
  wire [0:0] v_4115;
  function [0:0] mux_4115(input [0:0] sel);
    case (sel) 0: mux_4115 = 1'h0; 1: mux_4115 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4116;
  function [0:0] mux_4116(input [0:0] sel);
    case (sel) 0: mux_4116 = 1'h0; 1: mux_4116 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4117;
  wire [0:0] v_4118;
  wire [0:0] v_4119;
  wire [0:0] v_4120;
  function [0:0] mux_4120(input [0:0] sel);
    case (sel) 0: mux_4120 = 1'h0; 1: mux_4120 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4121;
  function [0:0] mux_4121(input [0:0] sel);
    case (sel) 0: mux_4121 = 1'h0; 1: mux_4121 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4122;
  wire [0:0] v_4123;
  wire [0:0] v_4124;
  wire [0:0] v_4125;
  wire [0:0] v_4126;
  wire [0:0] v_4127;
  function [0:0] mux_4127(input [0:0] sel);
    case (sel) 0: mux_4127 = 1'h0; 1: mux_4127 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4128;
  function [0:0] mux_4128(input [0:0] sel);
    case (sel) 0: mux_4128 = 1'h0; 1: mux_4128 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4129;
  wire [0:0] v_4130;
  wire [0:0] v_4131;
  wire [0:0] v_4132;
  function [0:0] mux_4132(input [0:0] sel);
    case (sel) 0: mux_4132 = 1'h0; 1: mux_4132 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4133;
  function [0:0] mux_4133(input [0:0] sel);
    case (sel) 0: mux_4133 = 1'h0; 1: mux_4133 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4134;
  wire [0:0] v_4135;
  wire [0:0] v_4136;
  wire [0:0] v_4137;
  wire [0:0] v_4138;
  wire [0:0] v_4139;
  function [0:0] mux_4139(input [0:0] sel);
    case (sel) 0: mux_4139 = 1'h0; 1: mux_4139 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4140;
  wire [0:0] v_4141;
  wire [0:0] v_4142;
  wire [0:0] v_4143;
  wire [0:0] v_4144;
  function [0:0] mux_4144(input [0:0] sel);
    case (sel) 0: mux_4144 = 1'h0; 1: mux_4144 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4145;
  wire [0:0] v_4146;
  wire [0:0] v_4147;
  wire [0:0] v_4148;
  function [0:0] mux_4148(input [0:0] sel);
    case (sel) 0: mux_4148 = 1'h0; 1: mux_4148 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4149;
  function [0:0] mux_4149(input [0:0] sel);
    case (sel) 0: mux_4149 = 1'h0; 1: mux_4149 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4150 = 1'h0;
  wire [0:0] v_4151;
  wire [0:0] v_4152;
  wire [0:0] act_4153;
  wire [0:0] v_4154;
  wire [0:0] v_4155;
  wire [0:0] v_4156;
  reg [0:0] v_4157 = 1'h0;
  wire [0:0] v_4158;
  wire [0:0] v_4159;
  wire [0:0] act_4160;
  wire [0:0] v_4161;
  wire [0:0] v_4162;
  wire [0:0] v_4163;
  reg [0:0] v_4164 = 1'h0;
  wire [0:0] v_4165;
  wire [0:0] v_4166;
  wire [0:0] act_4167;
  wire [0:0] v_4168;
  wire [0:0] v_4169;
  wire [0:0] v_4170;
  wire [0:0] vin0_consume_en_4171;
  wire [0:0] vout_canPeek_4171;
  wire [7:0] vout_peek_4171;
  wire [0:0] v_4172;
  wire [0:0] v_4173;
  function [0:0] mux_4173(input [0:0] sel);
    case (sel) 0: mux_4173 = 1'h0; 1: mux_4173 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4174;
  wire [0:0] v_4175;
  wire [0:0] v_4176;
  wire [0:0] v_4177;
  wire [0:0] v_4178;
  function [0:0] mux_4178(input [0:0] sel);
    case (sel) 0: mux_4178 = 1'h0; 1: mux_4178 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4179;
  wire [0:0] vin0_consume_en_4180;
  wire [0:0] vout_canPeek_4180;
  wire [7:0] vout_peek_4180;
  wire [0:0] v_4181;
  wire [0:0] v_4182;
  function [0:0] mux_4182(input [0:0] sel);
    case (sel) 0: mux_4182 = 1'h0; 1: mux_4182 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4183;
  function [0:0] mux_4183(input [0:0] sel);
    case (sel) 0: mux_4183 = 1'h0; 1: mux_4183 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4184;
  wire [0:0] v_4185;
  wire [0:0] v_4186;
  wire [0:0] v_4187;
  wire [0:0] v_4188;
  wire [0:0] v_4189;
  wire [0:0] v_4190;
  function [0:0] mux_4190(input [0:0] sel);
    case (sel) 0: mux_4190 = 1'h0; 1: mux_4190 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4191;
  wire [0:0] v_4192;
  wire [0:0] v_4193;
  wire [0:0] v_4194;
  wire [0:0] v_4195;
  function [0:0] mux_4195(input [0:0] sel);
    case (sel) 0: mux_4195 = 1'h0; 1: mux_4195 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4196;
  wire [0:0] v_4197;
  wire [0:0] v_4198;
  wire [0:0] v_4199;
  function [0:0] mux_4199(input [0:0] sel);
    case (sel) 0: mux_4199 = 1'h0; 1: mux_4199 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4200;
  function [0:0] mux_4200(input [0:0] sel);
    case (sel) 0: mux_4200 = 1'h0; 1: mux_4200 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4201 = 1'h0;
  wire [0:0] v_4202;
  wire [0:0] v_4203;
  wire [0:0] act_4204;
  wire [0:0] v_4205;
  wire [0:0] v_4206;
  wire [0:0] v_4207;
  wire [0:0] vin0_consume_en_4208;
  wire [0:0] vout_canPeek_4208;
  wire [7:0] vout_peek_4208;
  wire [0:0] v_4209;
  wire [0:0] v_4210;
  function [0:0] mux_4210(input [0:0] sel);
    case (sel) 0: mux_4210 = 1'h0; 1: mux_4210 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4211;
  wire [0:0] v_4212;
  wire [0:0] v_4213;
  wire [0:0] v_4214;
  wire [0:0] v_4215;
  function [0:0] mux_4215(input [0:0] sel);
    case (sel) 0: mux_4215 = 1'h0; 1: mux_4215 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4216;
  wire [0:0] vin0_consume_en_4217;
  wire [0:0] vout_canPeek_4217;
  wire [7:0] vout_peek_4217;
  wire [0:0] v_4218;
  wire [0:0] v_4219;
  function [0:0] mux_4219(input [0:0] sel);
    case (sel) 0: mux_4219 = 1'h0; 1: mux_4219 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4220;
  function [0:0] mux_4220(input [0:0] sel);
    case (sel) 0: mux_4220 = 1'h0; 1: mux_4220 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4221;
  wire [0:0] v_4222;
  wire [0:0] v_4223;
  wire [0:0] v_4224;
  wire [0:0] v_4225;
  wire [0:0] v_4226;
  wire [0:0] v_4227;
  function [0:0] mux_4227(input [0:0] sel);
    case (sel) 0: mux_4227 = 1'h0; 1: mux_4227 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4228;
  function [0:0] mux_4228(input [0:0] sel);
    case (sel) 0: mux_4228 = 1'h0; 1: mux_4228 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4229;
  wire [0:0] v_4230;
  wire [0:0] v_4231;
  wire [0:0] v_4232;
  function [0:0] mux_4232(input [0:0] sel);
    case (sel) 0: mux_4232 = 1'h0; 1: mux_4232 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4233;
  function [0:0] mux_4233(input [0:0] sel);
    case (sel) 0: mux_4233 = 1'h0; 1: mux_4233 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4234;
  wire [0:0] v_4235;
  wire [0:0] v_4236;
  wire [0:0] v_4237;
  wire [0:0] v_4238;
  wire [0:0] v_4239;
  function [0:0] mux_4239(input [0:0] sel);
    case (sel) 0: mux_4239 = 1'h0; 1: mux_4239 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4240;
  wire [0:0] v_4241;
  wire [0:0] v_4242;
  wire [0:0] v_4243;
  wire [0:0] v_4244;
  function [0:0] mux_4244(input [0:0] sel);
    case (sel) 0: mux_4244 = 1'h0; 1: mux_4244 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4245;
  wire [0:0] v_4246;
  wire [0:0] v_4247;
  wire [0:0] v_4248;
  function [0:0] mux_4248(input [0:0] sel);
    case (sel) 0: mux_4248 = 1'h0; 1: mux_4248 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4249;
  function [0:0] mux_4249(input [0:0] sel);
    case (sel) 0: mux_4249 = 1'h0; 1: mux_4249 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4250 = 1'h0;
  wire [0:0] v_4251;
  wire [0:0] v_4252;
  wire [0:0] act_4253;
  wire [0:0] v_4254;
  wire [0:0] v_4255;
  wire [0:0] v_4256;
  reg [0:0] v_4257 = 1'h0;
  wire [0:0] v_4258;
  wire [0:0] v_4259;
  wire [0:0] act_4260;
  wire [0:0] v_4261;
  wire [0:0] v_4262;
  wire [0:0] v_4263;
  wire [0:0] vin0_consume_en_4264;
  wire [0:0] vout_canPeek_4264;
  wire [7:0] vout_peek_4264;
  wire [0:0] v_4265;
  wire [0:0] v_4266;
  function [0:0] mux_4266(input [0:0] sel);
    case (sel) 0: mux_4266 = 1'h0; 1: mux_4266 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4267;
  wire [0:0] v_4268;
  wire [0:0] v_4269;
  wire [0:0] v_4270;
  wire [0:0] v_4271;
  function [0:0] mux_4271(input [0:0] sel);
    case (sel) 0: mux_4271 = 1'h0; 1: mux_4271 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4272;
  wire [0:0] vin0_consume_en_4273;
  wire [0:0] vout_canPeek_4273;
  wire [7:0] vout_peek_4273;
  wire [0:0] v_4274;
  wire [0:0] v_4275;
  function [0:0] mux_4275(input [0:0] sel);
    case (sel) 0: mux_4275 = 1'h0; 1: mux_4275 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4276;
  function [0:0] mux_4276(input [0:0] sel);
    case (sel) 0: mux_4276 = 1'h0; 1: mux_4276 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4277;
  wire [0:0] v_4278;
  wire [0:0] v_4279;
  wire [0:0] v_4280;
  wire [0:0] v_4281;
  wire [0:0] v_4282;
  wire [0:0] v_4283;
  function [0:0] mux_4283(input [0:0] sel);
    case (sel) 0: mux_4283 = 1'h0; 1: mux_4283 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4284;
  wire [0:0] v_4285;
  wire [0:0] v_4286;
  wire [0:0] v_4287;
  wire [0:0] v_4288;
  function [0:0] mux_4288(input [0:0] sel);
    case (sel) 0: mux_4288 = 1'h0; 1: mux_4288 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4289;
  wire [0:0] v_4290;
  wire [0:0] v_4291;
  wire [0:0] v_4292;
  function [0:0] mux_4292(input [0:0] sel);
    case (sel) 0: mux_4292 = 1'h0; 1: mux_4292 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4293;
  function [0:0] mux_4293(input [0:0] sel);
    case (sel) 0: mux_4293 = 1'h0; 1: mux_4293 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4294 = 1'h0;
  wire [0:0] v_4295;
  wire [0:0] v_4296;
  wire [0:0] act_4297;
  wire [0:0] v_4298;
  wire [0:0] v_4299;
  wire [0:0] v_4300;
  wire [0:0] vin0_consume_en_4301;
  wire [0:0] vout_canPeek_4301;
  wire [7:0] vout_peek_4301;
  wire [0:0] v_4302;
  wire [0:0] v_4303;
  function [0:0] mux_4303(input [0:0] sel);
    case (sel) 0: mux_4303 = 1'h0; 1: mux_4303 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4304;
  wire [0:0] v_4305;
  wire [0:0] v_4306;
  wire [0:0] v_4307;
  wire [0:0] v_4308;
  function [0:0] mux_4308(input [0:0] sel);
    case (sel) 0: mux_4308 = 1'h0; 1: mux_4308 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4309;
  wire [0:0] vin0_consume_en_4310;
  wire [0:0] vout_canPeek_4310;
  wire [7:0] vout_peek_4310;
  wire [0:0] v_4311;
  wire [0:0] v_4312;
  function [0:0] mux_4312(input [0:0] sel);
    case (sel) 0: mux_4312 = 1'h0; 1: mux_4312 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4313;
  function [0:0] mux_4313(input [0:0] sel);
    case (sel) 0: mux_4313 = 1'h0; 1: mux_4313 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4314;
  wire [0:0] v_4315;
  wire [0:0] v_4316;
  wire [0:0] v_4317;
  wire [0:0] v_4318;
  wire [0:0] v_4319;
  wire [0:0] v_4320;
  function [0:0] mux_4320(input [0:0] sel);
    case (sel) 0: mux_4320 = 1'h0; 1: mux_4320 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4321;
  function [0:0] mux_4321(input [0:0] sel);
    case (sel) 0: mux_4321 = 1'h0; 1: mux_4321 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4322;
  wire [0:0] v_4323;
  wire [0:0] v_4324;
  wire [0:0] v_4325;
  function [0:0] mux_4325(input [0:0] sel);
    case (sel) 0: mux_4325 = 1'h0; 1: mux_4325 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4326;
  function [0:0] mux_4326(input [0:0] sel);
    case (sel) 0: mux_4326 = 1'h0; 1: mux_4326 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4327;
  wire [0:0] v_4328;
  wire [0:0] v_4329;
  wire [0:0] v_4330;
  wire [0:0] v_4331;
  wire [0:0] v_4332;
  function [0:0] mux_4332(input [0:0] sel);
    case (sel) 0: mux_4332 = 1'h0; 1: mux_4332 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4333;
  function [0:0] mux_4333(input [0:0] sel);
    case (sel) 0: mux_4333 = 1'h0; 1: mux_4333 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4334;
  wire [0:0] v_4335;
  wire [0:0] v_4336;
  wire [0:0] v_4337;
  function [0:0] mux_4337(input [0:0] sel);
    case (sel) 0: mux_4337 = 1'h0; 1: mux_4337 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4338;
  function [0:0] mux_4338(input [0:0] sel);
    case (sel) 0: mux_4338 = 1'h0; 1: mux_4338 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4339;
  wire [0:0] v_4340;
  wire [0:0] v_4341;
  wire [0:0] v_4342;
  wire [0:0] v_4343;
  wire [0:0] v_4344;
  function [0:0] mux_4344(input [0:0] sel);
    case (sel) 0: mux_4344 = 1'h0; 1: mux_4344 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4345;
  function [0:0] mux_4345(input [0:0] sel);
    case (sel) 0: mux_4345 = 1'h0; 1: mux_4345 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4346;
  wire [0:0] v_4347;
  wire [0:0] v_4348;
  wire [0:0] v_4349;
  function [0:0] mux_4349(input [0:0] sel);
    case (sel) 0: mux_4349 = 1'h0; 1: mux_4349 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4350;
  function [0:0] mux_4350(input [0:0] sel);
    case (sel) 0: mux_4350 = 1'h0; 1: mux_4350 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4351;
  wire [0:0] v_4352;
  wire [0:0] v_4353;
  wire [0:0] v_4354;
  wire [0:0] v_4355;
  wire [0:0] v_4356;
  function [0:0] mux_4356(input [0:0] sel);
    case (sel) 0: mux_4356 = 1'h0; 1: mux_4356 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4357;
  function [0:0] mux_4357(input [0:0] sel);
    case (sel) 0: mux_4357 = 1'h0; 1: mux_4357 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4358;
  wire [0:0] v_4359;
  wire [0:0] v_4360;
  wire [0:0] v_4361;
  function [0:0] mux_4361(input [0:0] sel);
    case (sel) 0: mux_4361 = 1'h0; 1: mux_4361 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4362;
  function [0:0] mux_4362(input [0:0] sel);
    case (sel) 0: mux_4362 = 1'h0; 1: mux_4362 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4363;
  wire [0:0] v_4364;
  wire [0:0] v_4365;
  wire [0:0] v_4366;
  wire [0:0] v_4367;
  wire [0:0] v_4368;
  function [0:0] mux_4368(input [0:0] sel);
    case (sel) 0: mux_4368 = 1'h0; 1: mux_4368 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4369;
  function [0:0] mux_4369(input [0:0] sel);
    case (sel) 0: mux_4369 = 1'h0; 1: mux_4369 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4370;
  wire [0:0] v_4371;
  wire [0:0] v_4372;
  wire [0:0] v_4373;
  function [0:0] mux_4373(input [0:0] sel);
    case (sel) 0: mux_4373 = 1'h0; 1: mux_4373 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4374;
  function [0:0] mux_4374(input [0:0] sel);
    case (sel) 0: mux_4374 = 1'h0; 1: mux_4374 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4375;
  wire [0:0] v_4376;
  wire [0:0] v_4377;
  wire [0:0] v_4378;
  wire [0:0] v_4379;
  wire [0:0] v_4380;
  function [0:0] mux_4380(input [0:0] sel);
    case (sel) 0: mux_4380 = 1'h0; 1: mux_4380 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4381;
  wire [0:0] v_4382;
  wire [0:0] v_4383;
  wire [0:0] v_4384;
  reg [0:0] v_4385 = 1'h0;
  wire [0:0] v_4386;
  wire [0:0] v_4387;
  wire [0:0] act_4388;
  wire [0:0] v_4389;
  wire [0:0] v_4390;
  wire [0:0] v_4391;
  wire [0:0] v_4392;
  wire [0:0] v_4393;
  wire [0:0] v_4394;
  function [0:0] mux_4394(input [0:0] sel);
    case (sel) 0: mux_4394 = 1'h0; 1: mux_4394 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4395;
  wire [0:0] v_4396;
  wire [0:0] v_4397;
  reg [0:0] v_4398 = 1'h0;
  wire [0:0] v_4399;
  wire [0:0] v_4400;
  wire [0:0] act_4401;
  wire [0:0] v_4402;
  wire [0:0] v_4403;
  wire [0:0] v_4404;
  reg [0:0] v_4405 = 1'h0;
  wire [0:0] v_4406;
  wire [0:0] v_4407;
  wire [0:0] act_4408;
  wire [0:0] v_4409;
  wire [0:0] v_4410;
  wire [0:0] v_4411;
  reg [0:0] v_4412 = 1'h0;
  wire [0:0] v_4413;
  wire [0:0] v_4414;
  wire [0:0] act_4415;
  wire [0:0] v_4416;
  wire [0:0] v_4417;
  wire [0:0] v_4418;
  reg [0:0] v_4419 = 1'h0;
  wire [0:0] v_4420;
  wire [0:0] v_4421;
  wire [0:0] act_4422;
  wire [0:0] v_4423;
  wire [0:0] v_4424;
  wire [0:0] v_4425;
  reg [0:0] v_4426 = 1'h0;
  wire [0:0] v_4427;
  wire [0:0] v_4428;
  wire [0:0] act_4429;
  wire [0:0] v_4430;
  wire [0:0] v_4431;
  wire [0:0] v_4432;
  reg [0:0] v_4433 = 1'h0;
  wire [0:0] v_4434;
  wire [0:0] v_4435;
  wire [0:0] act_4436;
  wire [0:0] v_4437;
  wire [0:0] v_4438;
  wire [0:0] v_4439;
  reg [0:0] v_4440 = 1'h0;
  wire [0:0] v_4441;
  wire [0:0] v_4442;
  wire [0:0] act_4443;
  wire [0:0] v_4444;
  wire [0:0] v_4445;
  wire [0:0] v_4446;
  wire [0:0] vin0_consume_en_4447;
  wire [0:0] vout_canPeek_4447;
  wire [7:0] vout_peek_4447;
  wire [0:0] v_4448;
  wire [0:0] v_4449;
  function [0:0] mux_4449(input [0:0] sel);
    case (sel) 0: mux_4449 = 1'h0; 1: mux_4449 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4450;
  wire [0:0] v_4451;
  wire [0:0] v_4452;
  wire [0:0] v_4453;
  wire [0:0] v_4454;
  function [0:0] mux_4454(input [0:0] sel);
    case (sel) 0: mux_4454 = 1'h0; 1: mux_4454 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4455;
  wire [0:0] vin0_consume_en_4456;
  wire [0:0] vout_canPeek_4456;
  wire [7:0] vout_peek_4456;
  wire [0:0] v_4457;
  wire [0:0] v_4458;
  function [0:0] mux_4458(input [0:0] sel);
    case (sel) 0: mux_4458 = 1'h0; 1: mux_4458 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4459;
  function [0:0] mux_4459(input [0:0] sel);
    case (sel) 0: mux_4459 = 1'h0; 1: mux_4459 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4460;
  wire [0:0] v_4461;
  wire [0:0] v_4462;
  wire [0:0] v_4463;
  wire [0:0] v_4464;
  wire [0:0] v_4465;
  wire [0:0] v_4466;
  function [0:0] mux_4466(input [0:0] sel);
    case (sel) 0: mux_4466 = 1'h0; 1: mux_4466 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4467;
  wire [0:0] v_4468;
  wire [0:0] v_4469;
  wire [0:0] v_4470;
  wire [0:0] v_4471;
  function [0:0] mux_4471(input [0:0] sel);
    case (sel) 0: mux_4471 = 1'h0; 1: mux_4471 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4472;
  wire [0:0] v_4473;
  wire [0:0] v_4474;
  wire [0:0] v_4475;
  function [0:0] mux_4475(input [0:0] sel);
    case (sel) 0: mux_4475 = 1'h0; 1: mux_4475 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4476;
  function [0:0] mux_4476(input [0:0] sel);
    case (sel) 0: mux_4476 = 1'h0; 1: mux_4476 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4477 = 1'h0;
  wire [0:0] v_4478;
  wire [0:0] v_4479;
  wire [0:0] act_4480;
  wire [0:0] v_4481;
  wire [0:0] v_4482;
  wire [0:0] v_4483;
  wire [0:0] vin0_consume_en_4484;
  wire [0:0] vout_canPeek_4484;
  wire [7:0] vout_peek_4484;
  wire [0:0] v_4485;
  wire [0:0] v_4486;
  function [0:0] mux_4486(input [0:0] sel);
    case (sel) 0: mux_4486 = 1'h0; 1: mux_4486 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4487;
  wire [0:0] v_4488;
  wire [0:0] v_4489;
  wire [0:0] v_4490;
  wire [0:0] v_4491;
  function [0:0] mux_4491(input [0:0] sel);
    case (sel) 0: mux_4491 = 1'h0; 1: mux_4491 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4492;
  wire [0:0] vin0_consume_en_4493;
  wire [0:0] vout_canPeek_4493;
  wire [7:0] vout_peek_4493;
  wire [0:0] v_4494;
  wire [0:0] v_4495;
  function [0:0] mux_4495(input [0:0] sel);
    case (sel) 0: mux_4495 = 1'h0; 1: mux_4495 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4496;
  function [0:0] mux_4496(input [0:0] sel);
    case (sel) 0: mux_4496 = 1'h0; 1: mux_4496 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4497;
  wire [0:0] v_4498;
  wire [0:0] v_4499;
  wire [0:0] v_4500;
  wire [0:0] v_4501;
  wire [0:0] v_4502;
  wire [0:0] v_4503;
  function [0:0] mux_4503(input [0:0] sel);
    case (sel) 0: mux_4503 = 1'h0; 1: mux_4503 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4504;
  function [0:0] mux_4504(input [0:0] sel);
    case (sel) 0: mux_4504 = 1'h0; 1: mux_4504 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4505;
  wire [0:0] v_4506;
  wire [0:0] v_4507;
  wire [0:0] v_4508;
  function [0:0] mux_4508(input [0:0] sel);
    case (sel) 0: mux_4508 = 1'h0; 1: mux_4508 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4509;
  function [0:0] mux_4509(input [0:0] sel);
    case (sel) 0: mux_4509 = 1'h0; 1: mux_4509 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4510;
  wire [0:0] v_4511;
  wire [0:0] v_4512;
  wire [0:0] v_4513;
  wire [0:0] v_4514;
  wire [0:0] v_4515;
  function [0:0] mux_4515(input [0:0] sel);
    case (sel) 0: mux_4515 = 1'h0; 1: mux_4515 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4516;
  wire [0:0] v_4517;
  wire [0:0] v_4518;
  wire [0:0] v_4519;
  wire [0:0] v_4520;
  function [0:0] mux_4520(input [0:0] sel);
    case (sel) 0: mux_4520 = 1'h0; 1: mux_4520 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4521;
  wire [0:0] v_4522;
  wire [0:0] v_4523;
  wire [0:0] v_4524;
  function [0:0] mux_4524(input [0:0] sel);
    case (sel) 0: mux_4524 = 1'h0; 1: mux_4524 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4525;
  function [0:0] mux_4525(input [0:0] sel);
    case (sel) 0: mux_4525 = 1'h0; 1: mux_4525 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4526 = 1'h0;
  wire [0:0] v_4527;
  wire [0:0] v_4528;
  wire [0:0] act_4529;
  wire [0:0] v_4530;
  wire [0:0] v_4531;
  wire [0:0] v_4532;
  reg [0:0] v_4533 = 1'h0;
  wire [0:0] v_4534;
  wire [0:0] v_4535;
  wire [0:0] act_4536;
  wire [0:0] v_4537;
  wire [0:0] v_4538;
  wire [0:0] v_4539;
  wire [0:0] vin0_consume_en_4540;
  wire [0:0] vout_canPeek_4540;
  wire [7:0] vout_peek_4540;
  wire [0:0] v_4541;
  wire [0:0] v_4542;
  function [0:0] mux_4542(input [0:0] sel);
    case (sel) 0: mux_4542 = 1'h0; 1: mux_4542 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4543;
  wire [0:0] v_4544;
  wire [0:0] v_4545;
  wire [0:0] v_4546;
  wire [0:0] v_4547;
  function [0:0] mux_4547(input [0:0] sel);
    case (sel) 0: mux_4547 = 1'h0; 1: mux_4547 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4548;
  wire [0:0] vin0_consume_en_4549;
  wire [0:0] vout_canPeek_4549;
  wire [7:0] vout_peek_4549;
  wire [0:0] v_4550;
  wire [0:0] v_4551;
  function [0:0] mux_4551(input [0:0] sel);
    case (sel) 0: mux_4551 = 1'h0; 1: mux_4551 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4552;
  function [0:0] mux_4552(input [0:0] sel);
    case (sel) 0: mux_4552 = 1'h0; 1: mux_4552 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4553;
  wire [0:0] v_4554;
  wire [0:0] v_4555;
  wire [0:0] v_4556;
  wire [0:0] v_4557;
  wire [0:0] v_4558;
  wire [0:0] v_4559;
  function [0:0] mux_4559(input [0:0] sel);
    case (sel) 0: mux_4559 = 1'h0; 1: mux_4559 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4560;
  wire [0:0] v_4561;
  wire [0:0] v_4562;
  wire [0:0] v_4563;
  wire [0:0] v_4564;
  function [0:0] mux_4564(input [0:0] sel);
    case (sel) 0: mux_4564 = 1'h0; 1: mux_4564 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4565;
  wire [0:0] v_4566;
  wire [0:0] v_4567;
  wire [0:0] v_4568;
  function [0:0] mux_4568(input [0:0] sel);
    case (sel) 0: mux_4568 = 1'h0; 1: mux_4568 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4569;
  function [0:0] mux_4569(input [0:0] sel);
    case (sel) 0: mux_4569 = 1'h0; 1: mux_4569 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4570 = 1'h0;
  wire [0:0] v_4571;
  wire [0:0] v_4572;
  wire [0:0] act_4573;
  wire [0:0] v_4574;
  wire [0:0] v_4575;
  wire [0:0] v_4576;
  wire [0:0] vin0_consume_en_4577;
  wire [0:0] vout_canPeek_4577;
  wire [7:0] vout_peek_4577;
  wire [0:0] v_4578;
  wire [0:0] v_4579;
  function [0:0] mux_4579(input [0:0] sel);
    case (sel) 0: mux_4579 = 1'h0; 1: mux_4579 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4580;
  wire [0:0] v_4581;
  wire [0:0] v_4582;
  wire [0:0] v_4583;
  wire [0:0] v_4584;
  function [0:0] mux_4584(input [0:0] sel);
    case (sel) 0: mux_4584 = 1'h0; 1: mux_4584 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4585;
  wire [0:0] vin0_consume_en_4586;
  wire [0:0] vout_canPeek_4586;
  wire [7:0] vout_peek_4586;
  wire [0:0] v_4587;
  wire [0:0] v_4588;
  function [0:0] mux_4588(input [0:0] sel);
    case (sel) 0: mux_4588 = 1'h0; 1: mux_4588 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4589;
  function [0:0] mux_4589(input [0:0] sel);
    case (sel) 0: mux_4589 = 1'h0; 1: mux_4589 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4590;
  wire [0:0] v_4591;
  wire [0:0] v_4592;
  wire [0:0] v_4593;
  wire [0:0] v_4594;
  wire [0:0] v_4595;
  wire [0:0] v_4596;
  function [0:0] mux_4596(input [0:0] sel);
    case (sel) 0: mux_4596 = 1'h0; 1: mux_4596 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4597;
  function [0:0] mux_4597(input [0:0] sel);
    case (sel) 0: mux_4597 = 1'h0; 1: mux_4597 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4598;
  wire [0:0] v_4599;
  wire [0:0] v_4600;
  wire [0:0] v_4601;
  function [0:0] mux_4601(input [0:0] sel);
    case (sel) 0: mux_4601 = 1'h0; 1: mux_4601 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4602;
  function [0:0] mux_4602(input [0:0] sel);
    case (sel) 0: mux_4602 = 1'h0; 1: mux_4602 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4603;
  wire [0:0] v_4604;
  wire [0:0] v_4605;
  wire [0:0] v_4606;
  wire [0:0] v_4607;
  wire [0:0] v_4608;
  function [0:0] mux_4608(input [0:0] sel);
    case (sel) 0: mux_4608 = 1'h0; 1: mux_4608 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4609;
  function [0:0] mux_4609(input [0:0] sel);
    case (sel) 0: mux_4609 = 1'h0; 1: mux_4609 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4610;
  wire [0:0] v_4611;
  wire [0:0] v_4612;
  wire [0:0] v_4613;
  function [0:0] mux_4613(input [0:0] sel);
    case (sel) 0: mux_4613 = 1'h0; 1: mux_4613 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4614;
  function [0:0] mux_4614(input [0:0] sel);
    case (sel) 0: mux_4614 = 1'h0; 1: mux_4614 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4615;
  wire [0:0] v_4616;
  wire [0:0] v_4617;
  wire [0:0] v_4618;
  wire [0:0] v_4619;
  wire [0:0] v_4620;
  function [0:0] mux_4620(input [0:0] sel);
    case (sel) 0: mux_4620 = 1'h0; 1: mux_4620 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4621;
  wire [0:0] v_4622;
  wire [0:0] v_4623;
  wire [0:0] v_4624;
  wire [0:0] v_4625;
  function [0:0] mux_4625(input [0:0] sel);
    case (sel) 0: mux_4625 = 1'h0; 1: mux_4625 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4626;
  wire [0:0] v_4627;
  wire [0:0] v_4628;
  wire [0:0] v_4629;
  function [0:0] mux_4629(input [0:0] sel);
    case (sel) 0: mux_4629 = 1'h0; 1: mux_4629 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4630;
  function [0:0] mux_4630(input [0:0] sel);
    case (sel) 0: mux_4630 = 1'h0; 1: mux_4630 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4631 = 1'h0;
  wire [0:0] v_4632;
  wire [0:0] v_4633;
  wire [0:0] act_4634;
  wire [0:0] v_4635;
  wire [0:0] v_4636;
  wire [0:0] v_4637;
  reg [0:0] v_4638 = 1'h0;
  wire [0:0] v_4639;
  wire [0:0] v_4640;
  wire [0:0] act_4641;
  wire [0:0] v_4642;
  wire [0:0] v_4643;
  wire [0:0] v_4644;
  reg [0:0] v_4645 = 1'h0;
  wire [0:0] v_4646;
  wire [0:0] v_4647;
  wire [0:0] act_4648;
  wire [0:0] v_4649;
  wire [0:0] v_4650;
  wire [0:0] v_4651;
  wire [0:0] vin0_consume_en_4652;
  wire [0:0] vout_canPeek_4652;
  wire [7:0] vout_peek_4652;
  wire [0:0] v_4653;
  wire [0:0] v_4654;
  function [0:0] mux_4654(input [0:0] sel);
    case (sel) 0: mux_4654 = 1'h0; 1: mux_4654 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4655;
  wire [0:0] v_4656;
  wire [0:0] v_4657;
  wire [0:0] v_4658;
  wire [0:0] v_4659;
  function [0:0] mux_4659(input [0:0] sel);
    case (sel) 0: mux_4659 = 1'h0; 1: mux_4659 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4660;
  wire [0:0] vin0_consume_en_4661;
  wire [0:0] vout_canPeek_4661;
  wire [7:0] vout_peek_4661;
  wire [0:0] v_4662;
  wire [0:0] v_4663;
  function [0:0] mux_4663(input [0:0] sel);
    case (sel) 0: mux_4663 = 1'h0; 1: mux_4663 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4664;
  function [0:0] mux_4664(input [0:0] sel);
    case (sel) 0: mux_4664 = 1'h0; 1: mux_4664 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4665;
  wire [0:0] v_4666;
  wire [0:0] v_4667;
  wire [0:0] v_4668;
  wire [0:0] v_4669;
  wire [0:0] v_4670;
  wire [0:0] v_4671;
  function [0:0] mux_4671(input [0:0] sel);
    case (sel) 0: mux_4671 = 1'h0; 1: mux_4671 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4672;
  wire [0:0] v_4673;
  wire [0:0] v_4674;
  wire [0:0] v_4675;
  wire [0:0] v_4676;
  function [0:0] mux_4676(input [0:0] sel);
    case (sel) 0: mux_4676 = 1'h0; 1: mux_4676 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4677;
  wire [0:0] v_4678;
  wire [0:0] v_4679;
  wire [0:0] v_4680;
  function [0:0] mux_4680(input [0:0] sel);
    case (sel) 0: mux_4680 = 1'h0; 1: mux_4680 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4681;
  function [0:0] mux_4681(input [0:0] sel);
    case (sel) 0: mux_4681 = 1'h0; 1: mux_4681 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4682 = 1'h0;
  wire [0:0] v_4683;
  wire [0:0] v_4684;
  wire [0:0] act_4685;
  wire [0:0] v_4686;
  wire [0:0] v_4687;
  wire [0:0] v_4688;
  wire [0:0] vin0_consume_en_4689;
  wire [0:0] vout_canPeek_4689;
  wire [7:0] vout_peek_4689;
  wire [0:0] v_4690;
  wire [0:0] v_4691;
  function [0:0] mux_4691(input [0:0] sel);
    case (sel) 0: mux_4691 = 1'h0; 1: mux_4691 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4692;
  wire [0:0] v_4693;
  wire [0:0] v_4694;
  wire [0:0] v_4695;
  wire [0:0] v_4696;
  function [0:0] mux_4696(input [0:0] sel);
    case (sel) 0: mux_4696 = 1'h0; 1: mux_4696 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4697;
  wire [0:0] vin0_consume_en_4698;
  wire [0:0] vout_canPeek_4698;
  wire [7:0] vout_peek_4698;
  wire [0:0] v_4699;
  wire [0:0] v_4700;
  function [0:0] mux_4700(input [0:0] sel);
    case (sel) 0: mux_4700 = 1'h0; 1: mux_4700 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4701;
  function [0:0] mux_4701(input [0:0] sel);
    case (sel) 0: mux_4701 = 1'h0; 1: mux_4701 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4702;
  wire [0:0] v_4703;
  wire [0:0] v_4704;
  wire [0:0] v_4705;
  wire [0:0] v_4706;
  wire [0:0] v_4707;
  wire [0:0] v_4708;
  function [0:0] mux_4708(input [0:0] sel);
    case (sel) 0: mux_4708 = 1'h0; 1: mux_4708 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4709;
  function [0:0] mux_4709(input [0:0] sel);
    case (sel) 0: mux_4709 = 1'h0; 1: mux_4709 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4710;
  wire [0:0] v_4711;
  wire [0:0] v_4712;
  wire [0:0] v_4713;
  function [0:0] mux_4713(input [0:0] sel);
    case (sel) 0: mux_4713 = 1'h0; 1: mux_4713 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4714;
  function [0:0] mux_4714(input [0:0] sel);
    case (sel) 0: mux_4714 = 1'h0; 1: mux_4714 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4715;
  wire [0:0] v_4716;
  wire [0:0] v_4717;
  wire [0:0] v_4718;
  wire [0:0] v_4719;
  wire [0:0] v_4720;
  function [0:0] mux_4720(input [0:0] sel);
    case (sel) 0: mux_4720 = 1'h0; 1: mux_4720 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4721;
  wire [0:0] v_4722;
  wire [0:0] v_4723;
  wire [0:0] v_4724;
  wire [0:0] v_4725;
  function [0:0] mux_4725(input [0:0] sel);
    case (sel) 0: mux_4725 = 1'h0; 1: mux_4725 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4726;
  wire [0:0] v_4727;
  wire [0:0] v_4728;
  wire [0:0] v_4729;
  function [0:0] mux_4729(input [0:0] sel);
    case (sel) 0: mux_4729 = 1'h0; 1: mux_4729 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4730;
  function [0:0] mux_4730(input [0:0] sel);
    case (sel) 0: mux_4730 = 1'h0; 1: mux_4730 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4731 = 1'h0;
  wire [0:0] v_4732;
  wire [0:0] v_4733;
  wire [0:0] act_4734;
  wire [0:0] v_4735;
  wire [0:0] v_4736;
  wire [0:0] v_4737;
  reg [0:0] v_4738 = 1'h0;
  wire [0:0] v_4739;
  wire [0:0] v_4740;
  wire [0:0] act_4741;
  wire [0:0] v_4742;
  wire [0:0] v_4743;
  wire [0:0] v_4744;
  wire [0:0] vin0_consume_en_4745;
  wire [0:0] vout_canPeek_4745;
  wire [7:0] vout_peek_4745;
  wire [0:0] v_4746;
  wire [0:0] v_4747;
  function [0:0] mux_4747(input [0:0] sel);
    case (sel) 0: mux_4747 = 1'h0; 1: mux_4747 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4748;
  wire [0:0] v_4749;
  wire [0:0] v_4750;
  wire [0:0] v_4751;
  wire [0:0] v_4752;
  function [0:0] mux_4752(input [0:0] sel);
    case (sel) 0: mux_4752 = 1'h0; 1: mux_4752 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4753;
  wire [0:0] vin0_consume_en_4754;
  wire [0:0] vout_canPeek_4754;
  wire [7:0] vout_peek_4754;
  wire [0:0] v_4755;
  wire [0:0] v_4756;
  function [0:0] mux_4756(input [0:0] sel);
    case (sel) 0: mux_4756 = 1'h0; 1: mux_4756 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4757;
  function [0:0] mux_4757(input [0:0] sel);
    case (sel) 0: mux_4757 = 1'h0; 1: mux_4757 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4758;
  wire [0:0] v_4759;
  wire [0:0] v_4760;
  wire [0:0] v_4761;
  wire [0:0] v_4762;
  wire [0:0] v_4763;
  wire [0:0] v_4764;
  function [0:0] mux_4764(input [0:0] sel);
    case (sel) 0: mux_4764 = 1'h0; 1: mux_4764 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4765;
  wire [0:0] v_4766;
  wire [0:0] v_4767;
  wire [0:0] v_4768;
  wire [0:0] v_4769;
  function [0:0] mux_4769(input [0:0] sel);
    case (sel) 0: mux_4769 = 1'h0; 1: mux_4769 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4770;
  wire [0:0] v_4771;
  wire [0:0] v_4772;
  wire [0:0] v_4773;
  function [0:0] mux_4773(input [0:0] sel);
    case (sel) 0: mux_4773 = 1'h0; 1: mux_4773 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4774;
  function [0:0] mux_4774(input [0:0] sel);
    case (sel) 0: mux_4774 = 1'h0; 1: mux_4774 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4775 = 1'h0;
  wire [0:0] v_4776;
  wire [0:0] v_4777;
  wire [0:0] act_4778;
  wire [0:0] v_4779;
  wire [0:0] v_4780;
  wire [0:0] v_4781;
  wire [0:0] vin0_consume_en_4782;
  wire [0:0] vout_canPeek_4782;
  wire [7:0] vout_peek_4782;
  wire [0:0] v_4783;
  wire [0:0] v_4784;
  function [0:0] mux_4784(input [0:0] sel);
    case (sel) 0: mux_4784 = 1'h0; 1: mux_4784 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4785;
  wire [0:0] v_4786;
  wire [0:0] v_4787;
  wire [0:0] v_4788;
  wire [0:0] v_4789;
  function [0:0] mux_4789(input [0:0] sel);
    case (sel) 0: mux_4789 = 1'h0; 1: mux_4789 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4790;
  wire [0:0] vin0_consume_en_4791;
  wire [0:0] vout_canPeek_4791;
  wire [7:0] vout_peek_4791;
  wire [0:0] v_4792;
  wire [0:0] v_4793;
  function [0:0] mux_4793(input [0:0] sel);
    case (sel) 0: mux_4793 = 1'h0; 1: mux_4793 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4794;
  function [0:0] mux_4794(input [0:0] sel);
    case (sel) 0: mux_4794 = 1'h0; 1: mux_4794 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4795;
  wire [0:0] v_4796;
  wire [0:0] v_4797;
  wire [0:0] v_4798;
  wire [0:0] v_4799;
  wire [0:0] v_4800;
  wire [0:0] v_4801;
  function [0:0] mux_4801(input [0:0] sel);
    case (sel) 0: mux_4801 = 1'h0; 1: mux_4801 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4802;
  function [0:0] mux_4802(input [0:0] sel);
    case (sel) 0: mux_4802 = 1'h0; 1: mux_4802 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4803;
  wire [0:0] v_4804;
  wire [0:0] v_4805;
  wire [0:0] v_4806;
  function [0:0] mux_4806(input [0:0] sel);
    case (sel) 0: mux_4806 = 1'h0; 1: mux_4806 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4807;
  function [0:0] mux_4807(input [0:0] sel);
    case (sel) 0: mux_4807 = 1'h0; 1: mux_4807 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4808;
  wire [0:0] v_4809;
  wire [0:0] v_4810;
  wire [0:0] v_4811;
  wire [0:0] v_4812;
  wire [0:0] v_4813;
  function [0:0] mux_4813(input [0:0] sel);
    case (sel) 0: mux_4813 = 1'h0; 1: mux_4813 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4814;
  function [0:0] mux_4814(input [0:0] sel);
    case (sel) 0: mux_4814 = 1'h0; 1: mux_4814 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4815;
  wire [0:0] v_4816;
  wire [0:0] v_4817;
  wire [0:0] v_4818;
  function [0:0] mux_4818(input [0:0] sel);
    case (sel) 0: mux_4818 = 1'h0; 1: mux_4818 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4819;
  function [0:0] mux_4819(input [0:0] sel);
    case (sel) 0: mux_4819 = 1'h0; 1: mux_4819 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4820;
  wire [0:0] v_4821;
  wire [0:0] v_4822;
  wire [0:0] v_4823;
  wire [0:0] v_4824;
  wire [0:0] v_4825;
  function [0:0] mux_4825(input [0:0] sel);
    case (sel) 0: mux_4825 = 1'h0; 1: mux_4825 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4826;
  function [0:0] mux_4826(input [0:0] sel);
    case (sel) 0: mux_4826 = 1'h0; 1: mux_4826 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4827;
  wire [0:0] v_4828;
  wire [0:0] v_4829;
  wire [0:0] v_4830;
  function [0:0] mux_4830(input [0:0] sel);
    case (sel) 0: mux_4830 = 1'h0; 1: mux_4830 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4831;
  function [0:0] mux_4831(input [0:0] sel);
    case (sel) 0: mux_4831 = 1'h0; 1: mux_4831 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4832;
  wire [0:0] v_4833;
  wire [0:0] v_4834;
  wire [0:0] v_4835;
  wire [0:0] v_4836;
  wire [0:0] v_4837;
  function [0:0] mux_4837(input [0:0] sel);
    case (sel) 0: mux_4837 = 1'h0; 1: mux_4837 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4838;
  wire [0:0] v_4839;
  wire [0:0] v_4840;
  wire [0:0] v_4841;
  wire [0:0] v_4842;
  function [0:0] mux_4842(input [0:0] sel);
    case (sel) 0: mux_4842 = 1'h0; 1: mux_4842 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4843;
  wire [0:0] v_4844;
  wire [0:0] v_4845;
  wire [0:0] v_4846;
  function [0:0] mux_4846(input [0:0] sel);
    case (sel) 0: mux_4846 = 1'h0; 1: mux_4846 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4847;
  function [0:0] mux_4847(input [0:0] sel);
    case (sel) 0: mux_4847 = 1'h0; 1: mux_4847 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4848 = 1'h0;
  wire [0:0] v_4849;
  wire [0:0] v_4850;
  wire [0:0] act_4851;
  wire [0:0] v_4852;
  wire [0:0] v_4853;
  wire [0:0] v_4854;
  reg [0:0] v_4855 = 1'h0;
  wire [0:0] v_4856;
  wire [0:0] v_4857;
  wire [0:0] act_4858;
  wire [0:0] v_4859;
  wire [0:0] v_4860;
  wire [0:0] v_4861;
  reg [0:0] v_4862 = 1'h0;
  wire [0:0] v_4863;
  wire [0:0] v_4864;
  wire [0:0] act_4865;
  wire [0:0] v_4866;
  wire [0:0] v_4867;
  wire [0:0] v_4868;
  reg [0:0] v_4869 = 1'h0;
  wire [0:0] v_4870;
  wire [0:0] v_4871;
  wire [0:0] act_4872;
  wire [0:0] v_4873;
  wire [0:0] v_4874;
  wire [0:0] v_4875;
  wire [0:0] vin0_consume_en_4876;
  wire [0:0] vout_canPeek_4876;
  wire [7:0] vout_peek_4876;
  wire [0:0] v_4877;
  wire [0:0] v_4878;
  function [0:0] mux_4878(input [0:0] sel);
    case (sel) 0: mux_4878 = 1'h0; 1: mux_4878 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4879;
  wire [0:0] v_4880;
  wire [0:0] v_4881;
  wire [0:0] v_4882;
  wire [0:0] v_4883;
  function [0:0] mux_4883(input [0:0] sel);
    case (sel) 0: mux_4883 = 1'h0; 1: mux_4883 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4884;
  wire [0:0] vin0_consume_en_4885;
  wire [0:0] vout_canPeek_4885;
  wire [7:0] vout_peek_4885;
  wire [0:0] v_4886;
  wire [0:0] v_4887;
  function [0:0] mux_4887(input [0:0] sel);
    case (sel) 0: mux_4887 = 1'h0; 1: mux_4887 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4888;
  function [0:0] mux_4888(input [0:0] sel);
    case (sel) 0: mux_4888 = 1'h0; 1: mux_4888 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4889;
  wire [0:0] v_4890;
  wire [0:0] v_4891;
  wire [0:0] v_4892;
  wire [0:0] v_4893;
  wire [0:0] v_4894;
  wire [0:0] v_4895;
  function [0:0] mux_4895(input [0:0] sel);
    case (sel) 0: mux_4895 = 1'h0; 1: mux_4895 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4896;
  wire [0:0] v_4897;
  wire [0:0] v_4898;
  wire [0:0] v_4899;
  wire [0:0] v_4900;
  function [0:0] mux_4900(input [0:0] sel);
    case (sel) 0: mux_4900 = 1'h0; 1: mux_4900 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4901;
  wire [0:0] v_4902;
  wire [0:0] v_4903;
  wire [0:0] v_4904;
  function [0:0] mux_4904(input [0:0] sel);
    case (sel) 0: mux_4904 = 1'h0; 1: mux_4904 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4905;
  function [0:0] mux_4905(input [0:0] sel);
    case (sel) 0: mux_4905 = 1'h0; 1: mux_4905 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4906 = 1'h0;
  wire [0:0] v_4907;
  wire [0:0] v_4908;
  wire [0:0] act_4909;
  wire [0:0] v_4910;
  wire [0:0] v_4911;
  wire [0:0] v_4912;
  wire [0:0] vin0_consume_en_4913;
  wire [0:0] vout_canPeek_4913;
  wire [7:0] vout_peek_4913;
  wire [0:0] v_4914;
  wire [0:0] v_4915;
  function [0:0] mux_4915(input [0:0] sel);
    case (sel) 0: mux_4915 = 1'h0; 1: mux_4915 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4916;
  wire [0:0] v_4917;
  wire [0:0] v_4918;
  wire [0:0] v_4919;
  wire [0:0] v_4920;
  function [0:0] mux_4920(input [0:0] sel);
    case (sel) 0: mux_4920 = 1'h0; 1: mux_4920 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4921;
  wire [0:0] vin0_consume_en_4922;
  wire [0:0] vout_canPeek_4922;
  wire [7:0] vout_peek_4922;
  wire [0:0] v_4923;
  wire [0:0] v_4924;
  function [0:0] mux_4924(input [0:0] sel);
    case (sel) 0: mux_4924 = 1'h0; 1: mux_4924 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4925;
  function [0:0] mux_4925(input [0:0] sel);
    case (sel) 0: mux_4925 = 1'h0; 1: mux_4925 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4926;
  wire [0:0] v_4927;
  wire [0:0] v_4928;
  wire [0:0] v_4929;
  wire [0:0] v_4930;
  wire [0:0] v_4931;
  wire [0:0] v_4932;
  function [0:0] mux_4932(input [0:0] sel);
    case (sel) 0: mux_4932 = 1'h0; 1: mux_4932 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4933;
  function [0:0] mux_4933(input [0:0] sel);
    case (sel) 0: mux_4933 = 1'h0; 1: mux_4933 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4934;
  wire [0:0] v_4935;
  wire [0:0] v_4936;
  wire [0:0] v_4937;
  function [0:0] mux_4937(input [0:0] sel);
    case (sel) 0: mux_4937 = 1'h0; 1: mux_4937 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4938;
  function [0:0] mux_4938(input [0:0] sel);
    case (sel) 0: mux_4938 = 1'h0; 1: mux_4938 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4939;
  wire [0:0] v_4940;
  wire [0:0] v_4941;
  wire [0:0] v_4942;
  wire [0:0] v_4943;
  wire [0:0] v_4944;
  function [0:0] mux_4944(input [0:0] sel);
    case (sel) 0: mux_4944 = 1'h0; 1: mux_4944 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4945;
  wire [0:0] v_4946;
  wire [0:0] v_4947;
  wire [0:0] v_4948;
  wire [0:0] v_4949;
  function [0:0] mux_4949(input [0:0] sel);
    case (sel) 0: mux_4949 = 1'h0; 1: mux_4949 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4950;
  wire [0:0] v_4951;
  wire [0:0] v_4952;
  wire [0:0] v_4953;
  function [0:0] mux_4953(input [0:0] sel);
    case (sel) 0: mux_4953 = 1'h0; 1: mux_4953 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4954;
  function [0:0] mux_4954(input [0:0] sel);
    case (sel) 0: mux_4954 = 1'h0; 1: mux_4954 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4955 = 1'h0;
  wire [0:0] v_4956;
  wire [0:0] v_4957;
  wire [0:0] act_4958;
  wire [0:0] v_4959;
  wire [0:0] v_4960;
  wire [0:0] v_4961;
  reg [0:0] v_4962 = 1'h0;
  wire [0:0] v_4963;
  wire [0:0] v_4964;
  wire [0:0] act_4965;
  wire [0:0] v_4966;
  wire [0:0] v_4967;
  wire [0:0] v_4968;
  wire [0:0] vin0_consume_en_4969;
  wire [0:0] vout_canPeek_4969;
  wire [7:0] vout_peek_4969;
  wire [0:0] v_4970;
  wire [0:0] v_4971;
  function [0:0] mux_4971(input [0:0] sel);
    case (sel) 0: mux_4971 = 1'h0; 1: mux_4971 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4972;
  wire [0:0] v_4973;
  wire [0:0] v_4974;
  wire [0:0] v_4975;
  wire [0:0] v_4976;
  function [0:0] mux_4976(input [0:0] sel);
    case (sel) 0: mux_4976 = 1'h0; 1: mux_4976 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4977;
  wire [0:0] vin0_consume_en_4978;
  wire [0:0] vout_canPeek_4978;
  wire [7:0] vout_peek_4978;
  wire [0:0] v_4979;
  wire [0:0] v_4980;
  function [0:0] mux_4980(input [0:0] sel);
    case (sel) 0: mux_4980 = 1'h0; 1: mux_4980 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4981;
  function [0:0] mux_4981(input [0:0] sel);
    case (sel) 0: mux_4981 = 1'h0; 1: mux_4981 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4982;
  wire [0:0] v_4983;
  wire [0:0] v_4984;
  wire [0:0] v_4985;
  wire [0:0] v_4986;
  wire [0:0] v_4987;
  wire [0:0] v_4988;
  function [0:0] mux_4988(input [0:0] sel);
    case (sel) 0: mux_4988 = 1'h0; 1: mux_4988 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4989;
  wire [0:0] v_4990;
  wire [0:0] v_4991;
  wire [0:0] v_4992;
  wire [0:0] v_4993;
  function [0:0] mux_4993(input [0:0] sel);
    case (sel) 0: mux_4993 = 1'h0; 1: mux_4993 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4994;
  wire [0:0] v_4995;
  wire [0:0] v_4996;
  wire [0:0] v_4997;
  function [0:0] mux_4997(input [0:0] sel);
    case (sel) 0: mux_4997 = 1'h0; 1: mux_4997 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4998;
  function [0:0] mux_4998(input [0:0] sel);
    case (sel) 0: mux_4998 = 1'h0; 1: mux_4998 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4999 = 1'h0;
  wire [0:0] v_5000;
  wire [0:0] v_5001;
  wire [0:0] act_5002;
  wire [0:0] v_5003;
  wire [0:0] v_5004;
  wire [0:0] v_5005;
  wire [0:0] vin0_consume_en_5006;
  wire [0:0] vout_canPeek_5006;
  wire [7:0] vout_peek_5006;
  wire [0:0] v_5007;
  wire [0:0] v_5008;
  function [0:0] mux_5008(input [0:0] sel);
    case (sel) 0: mux_5008 = 1'h0; 1: mux_5008 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5009;
  wire [0:0] v_5010;
  wire [0:0] v_5011;
  wire [0:0] v_5012;
  wire [0:0] v_5013;
  function [0:0] mux_5013(input [0:0] sel);
    case (sel) 0: mux_5013 = 1'h0; 1: mux_5013 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5014;
  wire [0:0] vin0_consume_en_5015;
  wire [0:0] vout_canPeek_5015;
  wire [7:0] vout_peek_5015;
  wire [0:0] v_5016;
  wire [0:0] v_5017;
  function [0:0] mux_5017(input [0:0] sel);
    case (sel) 0: mux_5017 = 1'h0; 1: mux_5017 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5018;
  function [0:0] mux_5018(input [0:0] sel);
    case (sel) 0: mux_5018 = 1'h0; 1: mux_5018 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5019;
  wire [0:0] v_5020;
  wire [0:0] v_5021;
  wire [0:0] v_5022;
  wire [0:0] v_5023;
  wire [0:0] v_5024;
  wire [0:0] v_5025;
  function [0:0] mux_5025(input [0:0] sel);
    case (sel) 0: mux_5025 = 1'h0; 1: mux_5025 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5026;
  function [0:0] mux_5026(input [0:0] sel);
    case (sel) 0: mux_5026 = 1'h0; 1: mux_5026 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5027;
  wire [0:0] v_5028;
  wire [0:0] v_5029;
  wire [0:0] v_5030;
  function [0:0] mux_5030(input [0:0] sel);
    case (sel) 0: mux_5030 = 1'h0; 1: mux_5030 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5031;
  function [0:0] mux_5031(input [0:0] sel);
    case (sel) 0: mux_5031 = 1'h0; 1: mux_5031 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5032;
  wire [0:0] v_5033;
  wire [0:0] v_5034;
  wire [0:0] v_5035;
  wire [0:0] v_5036;
  wire [0:0] v_5037;
  function [0:0] mux_5037(input [0:0] sel);
    case (sel) 0: mux_5037 = 1'h0; 1: mux_5037 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5038;
  function [0:0] mux_5038(input [0:0] sel);
    case (sel) 0: mux_5038 = 1'h0; 1: mux_5038 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5039;
  wire [0:0] v_5040;
  wire [0:0] v_5041;
  wire [0:0] v_5042;
  function [0:0] mux_5042(input [0:0] sel);
    case (sel) 0: mux_5042 = 1'h0; 1: mux_5042 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5043;
  function [0:0] mux_5043(input [0:0] sel);
    case (sel) 0: mux_5043 = 1'h0; 1: mux_5043 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5044;
  wire [0:0] v_5045;
  wire [0:0] v_5046;
  wire [0:0] v_5047;
  wire [0:0] v_5048;
  wire [0:0] v_5049;
  function [0:0] mux_5049(input [0:0] sel);
    case (sel) 0: mux_5049 = 1'h0; 1: mux_5049 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5050;
  wire [0:0] v_5051;
  wire [0:0] v_5052;
  wire [0:0] v_5053;
  wire [0:0] v_5054;
  function [0:0] mux_5054(input [0:0] sel);
    case (sel) 0: mux_5054 = 1'h0; 1: mux_5054 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5055;
  wire [0:0] v_5056;
  wire [0:0] v_5057;
  wire [0:0] v_5058;
  function [0:0] mux_5058(input [0:0] sel);
    case (sel) 0: mux_5058 = 1'h0; 1: mux_5058 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5059;
  function [0:0] mux_5059(input [0:0] sel);
    case (sel) 0: mux_5059 = 1'h0; 1: mux_5059 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5060 = 1'h0;
  wire [0:0] v_5061;
  wire [0:0] v_5062;
  wire [0:0] act_5063;
  wire [0:0] v_5064;
  wire [0:0] v_5065;
  wire [0:0] v_5066;
  reg [0:0] v_5067 = 1'h0;
  wire [0:0] v_5068;
  wire [0:0] v_5069;
  wire [0:0] act_5070;
  wire [0:0] v_5071;
  wire [0:0] v_5072;
  wire [0:0] v_5073;
  reg [0:0] v_5074 = 1'h0;
  wire [0:0] v_5075;
  wire [0:0] v_5076;
  wire [0:0] act_5077;
  wire [0:0] v_5078;
  wire [0:0] v_5079;
  wire [0:0] v_5080;
  wire [0:0] vin0_consume_en_5081;
  wire [0:0] vout_canPeek_5081;
  wire [7:0] vout_peek_5081;
  wire [0:0] v_5082;
  wire [0:0] v_5083;
  function [0:0] mux_5083(input [0:0] sel);
    case (sel) 0: mux_5083 = 1'h0; 1: mux_5083 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5084;
  wire [0:0] v_5085;
  wire [0:0] v_5086;
  wire [0:0] v_5087;
  wire [0:0] v_5088;
  function [0:0] mux_5088(input [0:0] sel);
    case (sel) 0: mux_5088 = 1'h0; 1: mux_5088 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5089;
  wire [0:0] vin0_consume_en_5090;
  wire [0:0] vout_canPeek_5090;
  wire [7:0] vout_peek_5090;
  wire [0:0] v_5091;
  wire [0:0] v_5092;
  function [0:0] mux_5092(input [0:0] sel);
    case (sel) 0: mux_5092 = 1'h0; 1: mux_5092 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5093;
  function [0:0] mux_5093(input [0:0] sel);
    case (sel) 0: mux_5093 = 1'h0; 1: mux_5093 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5094;
  wire [0:0] v_5095;
  wire [0:0] v_5096;
  wire [0:0] v_5097;
  wire [0:0] v_5098;
  wire [0:0] v_5099;
  wire [0:0] v_5100;
  function [0:0] mux_5100(input [0:0] sel);
    case (sel) 0: mux_5100 = 1'h0; 1: mux_5100 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5101;
  wire [0:0] v_5102;
  wire [0:0] v_5103;
  wire [0:0] v_5104;
  wire [0:0] v_5105;
  function [0:0] mux_5105(input [0:0] sel);
    case (sel) 0: mux_5105 = 1'h0; 1: mux_5105 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5106;
  wire [0:0] v_5107;
  wire [0:0] v_5108;
  wire [0:0] v_5109;
  function [0:0] mux_5109(input [0:0] sel);
    case (sel) 0: mux_5109 = 1'h0; 1: mux_5109 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5110;
  function [0:0] mux_5110(input [0:0] sel);
    case (sel) 0: mux_5110 = 1'h0; 1: mux_5110 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5111 = 1'h0;
  wire [0:0] v_5112;
  wire [0:0] v_5113;
  wire [0:0] act_5114;
  wire [0:0] v_5115;
  wire [0:0] v_5116;
  wire [0:0] v_5117;
  wire [0:0] vin0_consume_en_5118;
  wire [0:0] vout_canPeek_5118;
  wire [7:0] vout_peek_5118;
  wire [0:0] v_5119;
  wire [0:0] v_5120;
  function [0:0] mux_5120(input [0:0] sel);
    case (sel) 0: mux_5120 = 1'h0; 1: mux_5120 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5121;
  wire [0:0] v_5122;
  wire [0:0] v_5123;
  wire [0:0] v_5124;
  wire [0:0] v_5125;
  function [0:0] mux_5125(input [0:0] sel);
    case (sel) 0: mux_5125 = 1'h0; 1: mux_5125 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5126;
  wire [0:0] vin0_consume_en_5127;
  wire [0:0] vout_canPeek_5127;
  wire [7:0] vout_peek_5127;
  wire [0:0] v_5128;
  wire [0:0] v_5129;
  function [0:0] mux_5129(input [0:0] sel);
    case (sel) 0: mux_5129 = 1'h0; 1: mux_5129 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5130;
  function [0:0] mux_5130(input [0:0] sel);
    case (sel) 0: mux_5130 = 1'h0; 1: mux_5130 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5131;
  wire [0:0] v_5132;
  wire [0:0] v_5133;
  wire [0:0] v_5134;
  wire [0:0] v_5135;
  wire [0:0] v_5136;
  wire [0:0] v_5137;
  function [0:0] mux_5137(input [0:0] sel);
    case (sel) 0: mux_5137 = 1'h0; 1: mux_5137 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5138;
  function [0:0] mux_5138(input [0:0] sel);
    case (sel) 0: mux_5138 = 1'h0; 1: mux_5138 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5139;
  wire [0:0] v_5140;
  wire [0:0] v_5141;
  wire [0:0] v_5142;
  function [0:0] mux_5142(input [0:0] sel);
    case (sel) 0: mux_5142 = 1'h0; 1: mux_5142 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5143;
  function [0:0] mux_5143(input [0:0] sel);
    case (sel) 0: mux_5143 = 1'h0; 1: mux_5143 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5144;
  wire [0:0] v_5145;
  wire [0:0] v_5146;
  wire [0:0] v_5147;
  wire [0:0] v_5148;
  wire [0:0] v_5149;
  function [0:0] mux_5149(input [0:0] sel);
    case (sel) 0: mux_5149 = 1'h0; 1: mux_5149 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5150;
  wire [0:0] v_5151;
  wire [0:0] v_5152;
  wire [0:0] v_5153;
  wire [0:0] v_5154;
  function [0:0] mux_5154(input [0:0] sel);
    case (sel) 0: mux_5154 = 1'h0; 1: mux_5154 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5155;
  wire [0:0] v_5156;
  wire [0:0] v_5157;
  wire [0:0] v_5158;
  function [0:0] mux_5158(input [0:0] sel);
    case (sel) 0: mux_5158 = 1'h0; 1: mux_5158 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5159;
  function [0:0] mux_5159(input [0:0] sel);
    case (sel) 0: mux_5159 = 1'h0; 1: mux_5159 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5160 = 1'h0;
  wire [0:0] v_5161;
  wire [0:0] v_5162;
  wire [0:0] act_5163;
  wire [0:0] v_5164;
  wire [0:0] v_5165;
  wire [0:0] v_5166;
  reg [0:0] v_5167 = 1'h0;
  wire [0:0] v_5168;
  wire [0:0] v_5169;
  wire [0:0] act_5170;
  wire [0:0] v_5171;
  wire [0:0] v_5172;
  wire [0:0] v_5173;
  wire [0:0] vin0_consume_en_5174;
  wire [0:0] vout_canPeek_5174;
  wire [7:0] vout_peek_5174;
  wire [0:0] v_5175;
  wire [0:0] v_5176;
  function [0:0] mux_5176(input [0:0] sel);
    case (sel) 0: mux_5176 = 1'h0; 1: mux_5176 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5177;
  wire [0:0] v_5178;
  wire [0:0] v_5179;
  wire [0:0] v_5180;
  wire [0:0] v_5181;
  function [0:0] mux_5181(input [0:0] sel);
    case (sel) 0: mux_5181 = 1'h0; 1: mux_5181 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5182;
  wire [0:0] vin0_consume_en_5183;
  wire [0:0] vout_canPeek_5183;
  wire [7:0] vout_peek_5183;
  wire [0:0] v_5184;
  wire [0:0] v_5185;
  function [0:0] mux_5185(input [0:0] sel);
    case (sel) 0: mux_5185 = 1'h0; 1: mux_5185 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5186;
  function [0:0] mux_5186(input [0:0] sel);
    case (sel) 0: mux_5186 = 1'h0; 1: mux_5186 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5187;
  wire [0:0] v_5188;
  wire [0:0] v_5189;
  wire [0:0] v_5190;
  wire [0:0] v_5191;
  wire [0:0] v_5192;
  wire [0:0] v_5193;
  function [0:0] mux_5193(input [0:0] sel);
    case (sel) 0: mux_5193 = 1'h0; 1: mux_5193 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5194;
  wire [0:0] v_5195;
  wire [0:0] v_5196;
  wire [0:0] v_5197;
  wire [0:0] v_5198;
  function [0:0] mux_5198(input [0:0] sel);
    case (sel) 0: mux_5198 = 1'h0; 1: mux_5198 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5199;
  wire [0:0] v_5200;
  wire [0:0] v_5201;
  wire [0:0] v_5202;
  function [0:0] mux_5202(input [0:0] sel);
    case (sel) 0: mux_5202 = 1'h0; 1: mux_5202 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5203;
  function [0:0] mux_5203(input [0:0] sel);
    case (sel) 0: mux_5203 = 1'h0; 1: mux_5203 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5204 = 1'h0;
  wire [0:0] v_5205;
  wire [0:0] v_5206;
  wire [0:0] act_5207;
  wire [0:0] v_5208;
  wire [0:0] v_5209;
  wire [0:0] v_5210;
  wire [0:0] vin0_consume_en_5211;
  wire [0:0] vout_canPeek_5211;
  wire [7:0] vout_peek_5211;
  wire [0:0] v_5212;
  wire [0:0] v_5213;
  function [0:0] mux_5213(input [0:0] sel);
    case (sel) 0: mux_5213 = 1'h0; 1: mux_5213 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5214;
  wire [0:0] v_5215;
  wire [0:0] v_5216;
  wire [0:0] v_5217;
  wire [0:0] v_5218;
  function [0:0] mux_5218(input [0:0] sel);
    case (sel) 0: mux_5218 = 1'h0; 1: mux_5218 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5219;
  wire [0:0] vin0_consume_en_5220;
  wire [0:0] vout_canPeek_5220;
  wire [7:0] vout_peek_5220;
  wire [0:0] v_5221;
  wire [0:0] v_5222;
  function [0:0] mux_5222(input [0:0] sel);
    case (sel) 0: mux_5222 = 1'h0; 1: mux_5222 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5223;
  function [0:0] mux_5223(input [0:0] sel);
    case (sel) 0: mux_5223 = 1'h0; 1: mux_5223 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5224;
  wire [0:0] v_5225;
  wire [0:0] v_5226;
  wire [0:0] v_5227;
  wire [0:0] v_5228;
  wire [0:0] v_5229;
  wire [0:0] v_5230;
  function [0:0] mux_5230(input [0:0] sel);
    case (sel) 0: mux_5230 = 1'h0; 1: mux_5230 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5231;
  function [0:0] mux_5231(input [0:0] sel);
    case (sel) 0: mux_5231 = 1'h0; 1: mux_5231 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5232;
  wire [0:0] v_5233;
  wire [0:0] v_5234;
  wire [0:0] v_5235;
  function [0:0] mux_5235(input [0:0] sel);
    case (sel) 0: mux_5235 = 1'h0; 1: mux_5235 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5236;
  function [0:0] mux_5236(input [0:0] sel);
    case (sel) 0: mux_5236 = 1'h0; 1: mux_5236 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5237;
  wire [0:0] v_5238;
  wire [0:0] v_5239;
  wire [0:0] v_5240;
  wire [0:0] v_5241;
  wire [0:0] v_5242;
  function [0:0] mux_5242(input [0:0] sel);
    case (sel) 0: mux_5242 = 1'h0; 1: mux_5242 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5243;
  function [0:0] mux_5243(input [0:0] sel);
    case (sel) 0: mux_5243 = 1'h0; 1: mux_5243 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5244;
  wire [0:0] v_5245;
  wire [0:0] v_5246;
  wire [0:0] v_5247;
  function [0:0] mux_5247(input [0:0] sel);
    case (sel) 0: mux_5247 = 1'h0; 1: mux_5247 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5248;
  function [0:0] mux_5248(input [0:0] sel);
    case (sel) 0: mux_5248 = 1'h0; 1: mux_5248 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5249;
  wire [0:0] v_5250;
  wire [0:0] v_5251;
  wire [0:0] v_5252;
  wire [0:0] v_5253;
  wire [0:0] v_5254;
  function [0:0] mux_5254(input [0:0] sel);
    case (sel) 0: mux_5254 = 1'h0; 1: mux_5254 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5255;
  function [0:0] mux_5255(input [0:0] sel);
    case (sel) 0: mux_5255 = 1'h0; 1: mux_5255 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5256;
  wire [0:0] v_5257;
  wire [0:0] v_5258;
  wire [0:0] v_5259;
  function [0:0] mux_5259(input [0:0] sel);
    case (sel) 0: mux_5259 = 1'h0; 1: mux_5259 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5260;
  function [0:0] mux_5260(input [0:0] sel);
    case (sel) 0: mux_5260 = 1'h0; 1: mux_5260 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5261;
  wire [0:0] v_5262;
  wire [0:0] v_5263;
  wire [0:0] v_5264;
  wire [0:0] v_5265;
  wire [0:0] v_5266;
  function [0:0] mux_5266(input [0:0] sel);
    case (sel) 0: mux_5266 = 1'h0; 1: mux_5266 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5267;
  function [0:0] mux_5267(input [0:0] sel);
    case (sel) 0: mux_5267 = 1'h0; 1: mux_5267 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5268;
  wire [0:0] v_5269;
  wire [0:0] v_5270;
  wire [0:0] v_5271;
  function [0:0] mux_5271(input [0:0] sel);
    case (sel) 0: mux_5271 = 1'h0; 1: mux_5271 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5272;
  function [0:0] mux_5272(input [0:0] sel);
    case (sel) 0: mux_5272 = 1'h0; 1: mux_5272 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5273;
  wire [0:0] v_5274;
  wire [0:0] v_5275;
  wire [0:0] v_5276;
  wire [0:0] v_5277;
  wire [0:0] v_5278;
  function [0:0] mux_5278(input [0:0] sel);
    case (sel) 0: mux_5278 = 1'h0; 1: mux_5278 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5279;
  wire [0:0] v_5280;
  wire [0:0] v_5281;
  wire [0:0] v_5282;
  wire [0:0] v_5283;
  function [0:0] mux_5283(input [0:0] sel);
    case (sel) 0: mux_5283 = 1'h0; 1: mux_5283 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5284;
  wire [0:0] v_5285;
  wire [0:0] v_5286;
  wire [0:0] v_5287;
  function [0:0] mux_5287(input [0:0] sel);
    case (sel) 0: mux_5287 = 1'h0; 1: mux_5287 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5288;
  function [0:0] mux_5288(input [0:0] sel);
    case (sel) 0: mux_5288 = 1'h0; 1: mux_5288 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5289 = 1'h0;
  wire [0:0] v_5290;
  wire [0:0] v_5291;
  wire [0:0] act_5292;
  wire [0:0] v_5293;
  wire [0:0] v_5294;
  wire [0:0] v_5295;
  reg [0:0] v_5296 = 1'h0;
  wire [0:0] v_5297;
  wire [0:0] v_5298;
  wire [0:0] act_5299;
  wire [0:0] v_5300;
  wire [0:0] v_5301;
  wire [0:0] v_5302;
  reg [0:0] v_5303 = 1'h0;
  wire [0:0] v_5304;
  wire [0:0] v_5305;
  wire [0:0] act_5306;
  wire [0:0] v_5307;
  wire [0:0] v_5308;
  wire [0:0] v_5309;
  reg [0:0] v_5310 = 1'h0;
  wire [0:0] v_5311;
  wire [0:0] v_5312;
  wire [0:0] act_5313;
  wire [0:0] v_5314;
  wire [0:0] v_5315;
  wire [0:0] v_5316;
  reg [0:0] v_5317 = 1'h0;
  wire [0:0] v_5318;
  wire [0:0] v_5319;
  wire [0:0] act_5320;
  wire [0:0] v_5321;
  wire [0:0] v_5322;
  wire [0:0] v_5323;
  wire [0:0] vin0_consume_en_5324;
  wire [0:0] vout_canPeek_5324;
  wire [7:0] vout_peek_5324;
  wire [0:0] v_5325;
  wire [0:0] v_5326;
  function [0:0] mux_5326(input [0:0] sel);
    case (sel) 0: mux_5326 = 1'h0; 1: mux_5326 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5327;
  wire [0:0] v_5328;
  wire [0:0] v_5329;
  wire [0:0] v_5330;
  wire [0:0] v_5331;
  function [0:0] mux_5331(input [0:0] sel);
    case (sel) 0: mux_5331 = 1'h0; 1: mux_5331 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5332;
  wire [0:0] vin0_consume_en_5333;
  wire [0:0] vout_canPeek_5333;
  wire [7:0] vout_peek_5333;
  wire [0:0] v_5334;
  wire [0:0] v_5335;
  function [0:0] mux_5335(input [0:0] sel);
    case (sel) 0: mux_5335 = 1'h0; 1: mux_5335 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5336;
  function [0:0] mux_5336(input [0:0] sel);
    case (sel) 0: mux_5336 = 1'h0; 1: mux_5336 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5337;
  wire [0:0] v_5338;
  wire [0:0] v_5339;
  wire [0:0] v_5340;
  wire [0:0] v_5341;
  wire [0:0] v_5342;
  wire [0:0] v_5343;
  function [0:0] mux_5343(input [0:0] sel);
    case (sel) 0: mux_5343 = 1'h0; 1: mux_5343 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5344;
  wire [0:0] v_5345;
  wire [0:0] v_5346;
  wire [0:0] v_5347;
  wire [0:0] v_5348;
  function [0:0] mux_5348(input [0:0] sel);
    case (sel) 0: mux_5348 = 1'h0; 1: mux_5348 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5349;
  wire [0:0] v_5350;
  wire [0:0] v_5351;
  wire [0:0] v_5352;
  function [0:0] mux_5352(input [0:0] sel);
    case (sel) 0: mux_5352 = 1'h0; 1: mux_5352 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5353;
  function [0:0] mux_5353(input [0:0] sel);
    case (sel) 0: mux_5353 = 1'h0; 1: mux_5353 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5354 = 1'h0;
  wire [0:0] v_5355;
  wire [0:0] v_5356;
  wire [0:0] act_5357;
  wire [0:0] v_5358;
  wire [0:0] v_5359;
  wire [0:0] v_5360;
  wire [0:0] vin0_consume_en_5361;
  wire [0:0] vout_canPeek_5361;
  wire [7:0] vout_peek_5361;
  wire [0:0] v_5362;
  wire [0:0] v_5363;
  function [0:0] mux_5363(input [0:0] sel);
    case (sel) 0: mux_5363 = 1'h0; 1: mux_5363 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5364;
  wire [0:0] v_5365;
  wire [0:0] v_5366;
  wire [0:0] v_5367;
  wire [0:0] v_5368;
  function [0:0] mux_5368(input [0:0] sel);
    case (sel) 0: mux_5368 = 1'h0; 1: mux_5368 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5369;
  wire [0:0] vin0_consume_en_5370;
  wire [0:0] vout_canPeek_5370;
  wire [7:0] vout_peek_5370;
  wire [0:0] v_5371;
  wire [0:0] v_5372;
  function [0:0] mux_5372(input [0:0] sel);
    case (sel) 0: mux_5372 = 1'h0; 1: mux_5372 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5373;
  function [0:0] mux_5373(input [0:0] sel);
    case (sel) 0: mux_5373 = 1'h0; 1: mux_5373 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5374;
  wire [0:0] v_5375;
  wire [0:0] v_5376;
  wire [0:0] v_5377;
  wire [0:0] v_5378;
  wire [0:0] v_5379;
  wire [0:0] v_5380;
  function [0:0] mux_5380(input [0:0] sel);
    case (sel) 0: mux_5380 = 1'h0; 1: mux_5380 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5381;
  function [0:0] mux_5381(input [0:0] sel);
    case (sel) 0: mux_5381 = 1'h0; 1: mux_5381 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5382;
  wire [0:0] v_5383;
  wire [0:0] v_5384;
  wire [0:0] v_5385;
  function [0:0] mux_5385(input [0:0] sel);
    case (sel) 0: mux_5385 = 1'h0; 1: mux_5385 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5386;
  function [0:0] mux_5386(input [0:0] sel);
    case (sel) 0: mux_5386 = 1'h0; 1: mux_5386 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5387;
  wire [0:0] v_5388;
  wire [0:0] v_5389;
  wire [0:0] v_5390;
  wire [0:0] v_5391;
  wire [0:0] v_5392;
  function [0:0] mux_5392(input [0:0] sel);
    case (sel) 0: mux_5392 = 1'h0; 1: mux_5392 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5393;
  wire [0:0] v_5394;
  wire [0:0] v_5395;
  wire [0:0] v_5396;
  wire [0:0] v_5397;
  function [0:0] mux_5397(input [0:0] sel);
    case (sel) 0: mux_5397 = 1'h0; 1: mux_5397 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5398;
  wire [0:0] v_5399;
  wire [0:0] v_5400;
  wire [0:0] v_5401;
  function [0:0] mux_5401(input [0:0] sel);
    case (sel) 0: mux_5401 = 1'h0; 1: mux_5401 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5402;
  function [0:0] mux_5402(input [0:0] sel);
    case (sel) 0: mux_5402 = 1'h0; 1: mux_5402 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5403 = 1'h0;
  wire [0:0] v_5404;
  wire [0:0] v_5405;
  wire [0:0] act_5406;
  wire [0:0] v_5407;
  wire [0:0] v_5408;
  wire [0:0] v_5409;
  reg [0:0] v_5410 = 1'h0;
  wire [0:0] v_5411;
  wire [0:0] v_5412;
  wire [0:0] act_5413;
  wire [0:0] v_5414;
  wire [0:0] v_5415;
  wire [0:0] v_5416;
  wire [0:0] vin0_consume_en_5417;
  wire [0:0] vout_canPeek_5417;
  wire [7:0] vout_peek_5417;
  wire [0:0] v_5418;
  wire [0:0] v_5419;
  function [0:0] mux_5419(input [0:0] sel);
    case (sel) 0: mux_5419 = 1'h0; 1: mux_5419 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5420;
  wire [0:0] v_5421;
  wire [0:0] v_5422;
  wire [0:0] v_5423;
  wire [0:0] v_5424;
  function [0:0] mux_5424(input [0:0] sel);
    case (sel) 0: mux_5424 = 1'h0; 1: mux_5424 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5425;
  wire [0:0] vin0_consume_en_5426;
  wire [0:0] vout_canPeek_5426;
  wire [7:0] vout_peek_5426;
  wire [0:0] v_5427;
  wire [0:0] v_5428;
  function [0:0] mux_5428(input [0:0] sel);
    case (sel) 0: mux_5428 = 1'h0; 1: mux_5428 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5429;
  function [0:0] mux_5429(input [0:0] sel);
    case (sel) 0: mux_5429 = 1'h0; 1: mux_5429 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5430;
  wire [0:0] v_5431;
  wire [0:0] v_5432;
  wire [0:0] v_5433;
  wire [0:0] v_5434;
  wire [0:0] v_5435;
  wire [0:0] v_5436;
  function [0:0] mux_5436(input [0:0] sel);
    case (sel) 0: mux_5436 = 1'h0; 1: mux_5436 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5437;
  wire [0:0] v_5438;
  wire [0:0] v_5439;
  wire [0:0] v_5440;
  wire [0:0] v_5441;
  function [0:0] mux_5441(input [0:0] sel);
    case (sel) 0: mux_5441 = 1'h0; 1: mux_5441 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5442;
  wire [0:0] v_5443;
  wire [0:0] v_5444;
  wire [0:0] v_5445;
  function [0:0] mux_5445(input [0:0] sel);
    case (sel) 0: mux_5445 = 1'h0; 1: mux_5445 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5446;
  function [0:0] mux_5446(input [0:0] sel);
    case (sel) 0: mux_5446 = 1'h0; 1: mux_5446 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5447 = 1'h0;
  wire [0:0] v_5448;
  wire [0:0] v_5449;
  wire [0:0] act_5450;
  wire [0:0] v_5451;
  wire [0:0] v_5452;
  wire [0:0] v_5453;
  wire [0:0] vin0_consume_en_5454;
  wire [0:0] vout_canPeek_5454;
  wire [7:0] vout_peek_5454;
  wire [0:0] v_5455;
  wire [0:0] v_5456;
  function [0:0] mux_5456(input [0:0] sel);
    case (sel) 0: mux_5456 = 1'h0; 1: mux_5456 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5457;
  wire [0:0] v_5458;
  wire [0:0] v_5459;
  wire [0:0] v_5460;
  wire [0:0] v_5461;
  function [0:0] mux_5461(input [0:0] sel);
    case (sel) 0: mux_5461 = 1'h0; 1: mux_5461 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5462;
  wire [0:0] vin0_consume_en_5463;
  wire [0:0] vout_canPeek_5463;
  wire [7:0] vout_peek_5463;
  wire [0:0] v_5464;
  wire [0:0] v_5465;
  function [0:0] mux_5465(input [0:0] sel);
    case (sel) 0: mux_5465 = 1'h0; 1: mux_5465 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5466;
  function [0:0] mux_5466(input [0:0] sel);
    case (sel) 0: mux_5466 = 1'h0; 1: mux_5466 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5467;
  wire [0:0] v_5468;
  wire [0:0] v_5469;
  wire [0:0] v_5470;
  wire [0:0] v_5471;
  wire [0:0] v_5472;
  wire [0:0] v_5473;
  function [0:0] mux_5473(input [0:0] sel);
    case (sel) 0: mux_5473 = 1'h0; 1: mux_5473 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5474;
  function [0:0] mux_5474(input [0:0] sel);
    case (sel) 0: mux_5474 = 1'h0; 1: mux_5474 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5475;
  wire [0:0] v_5476;
  wire [0:0] v_5477;
  wire [0:0] v_5478;
  function [0:0] mux_5478(input [0:0] sel);
    case (sel) 0: mux_5478 = 1'h0; 1: mux_5478 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5479;
  function [0:0] mux_5479(input [0:0] sel);
    case (sel) 0: mux_5479 = 1'h0; 1: mux_5479 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5480;
  wire [0:0] v_5481;
  wire [0:0] v_5482;
  wire [0:0] v_5483;
  wire [0:0] v_5484;
  wire [0:0] v_5485;
  function [0:0] mux_5485(input [0:0] sel);
    case (sel) 0: mux_5485 = 1'h0; 1: mux_5485 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5486;
  function [0:0] mux_5486(input [0:0] sel);
    case (sel) 0: mux_5486 = 1'h0; 1: mux_5486 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5487;
  wire [0:0] v_5488;
  wire [0:0] v_5489;
  wire [0:0] v_5490;
  function [0:0] mux_5490(input [0:0] sel);
    case (sel) 0: mux_5490 = 1'h0; 1: mux_5490 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5491;
  function [0:0] mux_5491(input [0:0] sel);
    case (sel) 0: mux_5491 = 1'h0; 1: mux_5491 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5492;
  wire [0:0] v_5493;
  wire [0:0] v_5494;
  wire [0:0] v_5495;
  wire [0:0] v_5496;
  wire [0:0] v_5497;
  function [0:0] mux_5497(input [0:0] sel);
    case (sel) 0: mux_5497 = 1'h0; 1: mux_5497 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5498;
  wire [0:0] v_5499;
  wire [0:0] v_5500;
  wire [0:0] v_5501;
  wire [0:0] v_5502;
  function [0:0] mux_5502(input [0:0] sel);
    case (sel) 0: mux_5502 = 1'h0; 1: mux_5502 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5503;
  wire [0:0] v_5504;
  wire [0:0] v_5505;
  wire [0:0] v_5506;
  function [0:0] mux_5506(input [0:0] sel);
    case (sel) 0: mux_5506 = 1'h0; 1: mux_5506 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5507;
  function [0:0] mux_5507(input [0:0] sel);
    case (sel) 0: mux_5507 = 1'h0; 1: mux_5507 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5508 = 1'h0;
  wire [0:0] v_5509;
  wire [0:0] v_5510;
  wire [0:0] act_5511;
  wire [0:0] v_5512;
  wire [0:0] v_5513;
  wire [0:0] v_5514;
  reg [0:0] v_5515 = 1'h0;
  wire [0:0] v_5516;
  wire [0:0] v_5517;
  wire [0:0] act_5518;
  wire [0:0] v_5519;
  wire [0:0] v_5520;
  wire [0:0] v_5521;
  reg [0:0] v_5522 = 1'h0;
  wire [0:0] v_5523;
  wire [0:0] v_5524;
  wire [0:0] act_5525;
  wire [0:0] v_5526;
  wire [0:0] v_5527;
  wire [0:0] v_5528;
  wire [0:0] vin0_consume_en_5529;
  wire [0:0] vout_canPeek_5529;
  wire [7:0] vout_peek_5529;
  wire [0:0] v_5530;
  wire [0:0] v_5531;
  function [0:0] mux_5531(input [0:0] sel);
    case (sel) 0: mux_5531 = 1'h0; 1: mux_5531 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5532;
  wire [0:0] v_5533;
  wire [0:0] v_5534;
  wire [0:0] v_5535;
  wire [0:0] v_5536;
  function [0:0] mux_5536(input [0:0] sel);
    case (sel) 0: mux_5536 = 1'h0; 1: mux_5536 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5537;
  wire [0:0] vin0_consume_en_5538;
  wire [0:0] vout_canPeek_5538;
  wire [7:0] vout_peek_5538;
  wire [0:0] v_5539;
  wire [0:0] v_5540;
  function [0:0] mux_5540(input [0:0] sel);
    case (sel) 0: mux_5540 = 1'h0; 1: mux_5540 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5541;
  function [0:0] mux_5541(input [0:0] sel);
    case (sel) 0: mux_5541 = 1'h0; 1: mux_5541 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5542;
  wire [0:0] v_5543;
  wire [0:0] v_5544;
  wire [0:0] v_5545;
  wire [0:0] v_5546;
  wire [0:0] v_5547;
  wire [0:0] v_5548;
  function [0:0] mux_5548(input [0:0] sel);
    case (sel) 0: mux_5548 = 1'h0; 1: mux_5548 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5549;
  wire [0:0] v_5550;
  wire [0:0] v_5551;
  wire [0:0] v_5552;
  wire [0:0] v_5553;
  function [0:0] mux_5553(input [0:0] sel);
    case (sel) 0: mux_5553 = 1'h0; 1: mux_5553 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5554;
  wire [0:0] v_5555;
  wire [0:0] v_5556;
  wire [0:0] v_5557;
  function [0:0] mux_5557(input [0:0] sel);
    case (sel) 0: mux_5557 = 1'h0; 1: mux_5557 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5558;
  function [0:0] mux_5558(input [0:0] sel);
    case (sel) 0: mux_5558 = 1'h0; 1: mux_5558 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5559 = 1'h0;
  wire [0:0] v_5560;
  wire [0:0] v_5561;
  wire [0:0] act_5562;
  wire [0:0] v_5563;
  wire [0:0] v_5564;
  wire [0:0] v_5565;
  wire [0:0] vin0_consume_en_5566;
  wire [0:0] vout_canPeek_5566;
  wire [7:0] vout_peek_5566;
  wire [0:0] v_5567;
  wire [0:0] v_5568;
  function [0:0] mux_5568(input [0:0] sel);
    case (sel) 0: mux_5568 = 1'h0; 1: mux_5568 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5569;
  wire [0:0] v_5570;
  wire [0:0] v_5571;
  wire [0:0] v_5572;
  wire [0:0] v_5573;
  function [0:0] mux_5573(input [0:0] sel);
    case (sel) 0: mux_5573 = 1'h0; 1: mux_5573 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5574;
  wire [0:0] vin0_consume_en_5575;
  wire [0:0] vout_canPeek_5575;
  wire [7:0] vout_peek_5575;
  wire [0:0] v_5576;
  wire [0:0] v_5577;
  function [0:0] mux_5577(input [0:0] sel);
    case (sel) 0: mux_5577 = 1'h0; 1: mux_5577 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5578;
  function [0:0] mux_5578(input [0:0] sel);
    case (sel) 0: mux_5578 = 1'h0; 1: mux_5578 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5579;
  wire [0:0] v_5580;
  wire [0:0] v_5581;
  wire [0:0] v_5582;
  wire [0:0] v_5583;
  wire [0:0] v_5584;
  wire [0:0] v_5585;
  function [0:0] mux_5585(input [0:0] sel);
    case (sel) 0: mux_5585 = 1'h0; 1: mux_5585 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5586;
  function [0:0] mux_5586(input [0:0] sel);
    case (sel) 0: mux_5586 = 1'h0; 1: mux_5586 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5587;
  wire [0:0] v_5588;
  wire [0:0] v_5589;
  wire [0:0] v_5590;
  function [0:0] mux_5590(input [0:0] sel);
    case (sel) 0: mux_5590 = 1'h0; 1: mux_5590 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5591;
  function [0:0] mux_5591(input [0:0] sel);
    case (sel) 0: mux_5591 = 1'h0; 1: mux_5591 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5592;
  wire [0:0] v_5593;
  wire [0:0] v_5594;
  wire [0:0] v_5595;
  wire [0:0] v_5596;
  wire [0:0] v_5597;
  function [0:0] mux_5597(input [0:0] sel);
    case (sel) 0: mux_5597 = 1'h0; 1: mux_5597 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5598;
  wire [0:0] v_5599;
  wire [0:0] v_5600;
  wire [0:0] v_5601;
  wire [0:0] v_5602;
  function [0:0] mux_5602(input [0:0] sel);
    case (sel) 0: mux_5602 = 1'h0; 1: mux_5602 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5603;
  wire [0:0] v_5604;
  wire [0:0] v_5605;
  wire [0:0] v_5606;
  function [0:0] mux_5606(input [0:0] sel);
    case (sel) 0: mux_5606 = 1'h0; 1: mux_5606 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5607;
  function [0:0] mux_5607(input [0:0] sel);
    case (sel) 0: mux_5607 = 1'h0; 1: mux_5607 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5608 = 1'h0;
  wire [0:0] v_5609;
  wire [0:0] v_5610;
  wire [0:0] act_5611;
  wire [0:0] v_5612;
  wire [0:0] v_5613;
  wire [0:0] v_5614;
  reg [0:0] v_5615 = 1'h0;
  wire [0:0] v_5616;
  wire [0:0] v_5617;
  wire [0:0] act_5618;
  wire [0:0] v_5619;
  wire [0:0] v_5620;
  wire [0:0] v_5621;
  wire [0:0] vin0_consume_en_5622;
  wire [0:0] vout_canPeek_5622;
  wire [7:0] vout_peek_5622;
  wire [0:0] v_5623;
  wire [0:0] v_5624;
  function [0:0] mux_5624(input [0:0] sel);
    case (sel) 0: mux_5624 = 1'h0; 1: mux_5624 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5625;
  wire [0:0] v_5626;
  wire [0:0] v_5627;
  wire [0:0] v_5628;
  wire [0:0] v_5629;
  function [0:0] mux_5629(input [0:0] sel);
    case (sel) 0: mux_5629 = 1'h0; 1: mux_5629 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5630;
  wire [0:0] vin0_consume_en_5631;
  wire [0:0] vout_canPeek_5631;
  wire [7:0] vout_peek_5631;
  wire [0:0] v_5632;
  wire [0:0] v_5633;
  function [0:0] mux_5633(input [0:0] sel);
    case (sel) 0: mux_5633 = 1'h0; 1: mux_5633 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5634;
  function [0:0] mux_5634(input [0:0] sel);
    case (sel) 0: mux_5634 = 1'h0; 1: mux_5634 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5635;
  wire [0:0] v_5636;
  wire [0:0] v_5637;
  wire [0:0] v_5638;
  wire [0:0] v_5639;
  wire [0:0] v_5640;
  wire [0:0] v_5641;
  function [0:0] mux_5641(input [0:0] sel);
    case (sel) 0: mux_5641 = 1'h0; 1: mux_5641 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5642;
  wire [0:0] v_5643;
  wire [0:0] v_5644;
  wire [0:0] v_5645;
  wire [0:0] v_5646;
  function [0:0] mux_5646(input [0:0] sel);
    case (sel) 0: mux_5646 = 1'h0; 1: mux_5646 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5647;
  wire [0:0] v_5648;
  wire [0:0] v_5649;
  wire [0:0] v_5650;
  function [0:0] mux_5650(input [0:0] sel);
    case (sel) 0: mux_5650 = 1'h0; 1: mux_5650 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5651;
  function [0:0] mux_5651(input [0:0] sel);
    case (sel) 0: mux_5651 = 1'h0; 1: mux_5651 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5652 = 1'h0;
  wire [0:0] v_5653;
  wire [0:0] v_5654;
  wire [0:0] act_5655;
  wire [0:0] v_5656;
  wire [0:0] v_5657;
  wire [0:0] v_5658;
  wire [0:0] vin0_consume_en_5659;
  wire [0:0] vout_canPeek_5659;
  wire [7:0] vout_peek_5659;
  wire [0:0] v_5660;
  wire [0:0] v_5661;
  function [0:0] mux_5661(input [0:0] sel);
    case (sel) 0: mux_5661 = 1'h0; 1: mux_5661 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5662;
  wire [0:0] v_5663;
  wire [0:0] v_5664;
  wire [0:0] v_5665;
  wire [0:0] v_5666;
  function [0:0] mux_5666(input [0:0] sel);
    case (sel) 0: mux_5666 = 1'h0; 1: mux_5666 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5667;
  wire [0:0] vin0_consume_en_5668;
  wire [0:0] vout_canPeek_5668;
  wire [7:0] vout_peek_5668;
  wire [0:0] v_5669;
  wire [0:0] v_5670;
  function [0:0] mux_5670(input [0:0] sel);
    case (sel) 0: mux_5670 = 1'h0; 1: mux_5670 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5671;
  function [0:0] mux_5671(input [0:0] sel);
    case (sel) 0: mux_5671 = 1'h0; 1: mux_5671 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5672;
  wire [0:0] v_5673;
  wire [0:0] v_5674;
  wire [0:0] v_5675;
  wire [0:0] v_5676;
  wire [0:0] v_5677;
  wire [0:0] v_5678;
  function [0:0] mux_5678(input [0:0] sel);
    case (sel) 0: mux_5678 = 1'h0; 1: mux_5678 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5679;
  function [0:0] mux_5679(input [0:0] sel);
    case (sel) 0: mux_5679 = 1'h0; 1: mux_5679 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5680;
  wire [0:0] v_5681;
  wire [0:0] v_5682;
  wire [0:0] v_5683;
  function [0:0] mux_5683(input [0:0] sel);
    case (sel) 0: mux_5683 = 1'h0; 1: mux_5683 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5684;
  function [0:0] mux_5684(input [0:0] sel);
    case (sel) 0: mux_5684 = 1'h0; 1: mux_5684 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5685;
  wire [0:0] v_5686;
  wire [0:0] v_5687;
  wire [0:0] v_5688;
  wire [0:0] v_5689;
  wire [0:0] v_5690;
  function [0:0] mux_5690(input [0:0] sel);
    case (sel) 0: mux_5690 = 1'h0; 1: mux_5690 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5691;
  function [0:0] mux_5691(input [0:0] sel);
    case (sel) 0: mux_5691 = 1'h0; 1: mux_5691 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5692;
  wire [0:0] v_5693;
  wire [0:0] v_5694;
  wire [0:0] v_5695;
  function [0:0] mux_5695(input [0:0] sel);
    case (sel) 0: mux_5695 = 1'h0; 1: mux_5695 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5696;
  function [0:0] mux_5696(input [0:0] sel);
    case (sel) 0: mux_5696 = 1'h0; 1: mux_5696 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5697;
  wire [0:0] v_5698;
  wire [0:0] v_5699;
  wire [0:0] v_5700;
  wire [0:0] v_5701;
  wire [0:0] v_5702;
  function [0:0] mux_5702(input [0:0] sel);
    case (sel) 0: mux_5702 = 1'h0; 1: mux_5702 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5703;
  function [0:0] mux_5703(input [0:0] sel);
    case (sel) 0: mux_5703 = 1'h0; 1: mux_5703 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5704;
  wire [0:0] v_5705;
  wire [0:0] v_5706;
  wire [0:0] v_5707;
  function [0:0] mux_5707(input [0:0] sel);
    case (sel) 0: mux_5707 = 1'h0; 1: mux_5707 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5708;
  function [0:0] mux_5708(input [0:0] sel);
    case (sel) 0: mux_5708 = 1'h0; 1: mux_5708 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5709;
  wire [0:0] v_5710;
  wire [0:0] v_5711;
  wire [0:0] v_5712;
  wire [0:0] v_5713;
  wire [0:0] v_5714;
  function [0:0] mux_5714(input [0:0] sel);
    case (sel) 0: mux_5714 = 1'h0; 1: mux_5714 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5715;
  wire [0:0] v_5716;
  wire [0:0] v_5717;
  wire [0:0] v_5718;
  wire [0:0] v_5719;
  function [0:0] mux_5719(input [0:0] sel);
    case (sel) 0: mux_5719 = 1'h0; 1: mux_5719 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5720;
  wire [0:0] v_5721;
  wire [0:0] v_5722;
  wire [0:0] v_5723;
  function [0:0] mux_5723(input [0:0] sel);
    case (sel) 0: mux_5723 = 1'h0; 1: mux_5723 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5724;
  function [0:0] mux_5724(input [0:0] sel);
    case (sel) 0: mux_5724 = 1'h0; 1: mux_5724 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5725 = 1'h0;
  wire [0:0] v_5726;
  wire [0:0] v_5727;
  wire [0:0] act_5728;
  wire [0:0] v_5729;
  wire [0:0] v_5730;
  wire [0:0] v_5731;
  reg [0:0] v_5732 = 1'h0;
  wire [0:0] v_5733;
  wire [0:0] v_5734;
  wire [0:0] act_5735;
  wire [0:0] v_5736;
  wire [0:0] v_5737;
  wire [0:0] v_5738;
  reg [0:0] v_5739 = 1'h0;
  wire [0:0] v_5740;
  wire [0:0] v_5741;
  wire [0:0] act_5742;
  wire [0:0] v_5743;
  wire [0:0] v_5744;
  wire [0:0] v_5745;
  reg [0:0] v_5746 = 1'h0;
  wire [0:0] v_5747;
  wire [0:0] v_5748;
  wire [0:0] act_5749;
  wire [0:0] v_5750;
  wire [0:0] v_5751;
  wire [0:0] v_5752;
  wire [0:0] vin0_consume_en_5753;
  wire [0:0] vout_canPeek_5753;
  wire [7:0] vout_peek_5753;
  wire [0:0] v_5754;
  wire [0:0] v_5755;
  function [0:0] mux_5755(input [0:0] sel);
    case (sel) 0: mux_5755 = 1'h0; 1: mux_5755 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5756;
  wire [0:0] v_5757;
  wire [0:0] v_5758;
  wire [0:0] v_5759;
  wire [0:0] v_5760;
  function [0:0] mux_5760(input [0:0] sel);
    case (sel) 0: mux_5760 = 1'h0; 1: mux_5760 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5761;
  wire [0:0] vin0_consume_en_5762;
  wire [0:0] vout_canPeek_5762;
  wire [7:0] vout_peek_5762;
  wire [0:0] v_5763;
  wire [0:0] v_5764;
  function [0:0] mux_5764(input [0:0] sel);
    case (sel) 0: mux_5764 = 1'h0; 1: mux_5764 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5765;
  function [0:0] mux_5765(input [0:0] sel);
    case (sel) 0: mux_5765 = 1'h0; 1: mux_5765 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5766;
  wire [0:0] v_5767;
  wire [0:0] v_5768;
  wire [0:0] v_5769;
  wire [0:0] v_5770;
  wire [0:0] v_5771;
  wire [0:0] v_5772;
  function [0:0] mux_5772(input [0:0] sel);
    case (sel) 0: mux_5772 = 1'h0; 1: mux_5772 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5773;
  wire [0:0] v_5774;
  wire [0:0] v_5775;
  wire [0:0] v_5776;
  wire [0:0] v_5777;
  function [0:0] mux_5777(input [0:0] sel);
    case (sel) 0: mux_5777 = 1'h0; 1: mux_5777 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5778;
  wire [0:0] v_5779;
  wire [0:0] v_5780;
  wire [0:0] v_5781;
  function [0:0] mux_5781(input [0:0] sel);
    case (sel) 0: mux_5781 = 1'h0; 1: mux_5781 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5782;
  function [0:0] mux_5782(input [0:0] sel);
    case (sel) 0: mux_5782 = 1'h0; 1: mux_5782 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5783 = 1'h0;
  wire [0:0] v_5784;
  wire [0:0] v_5785;
  wire [0:0] act_5786;
  wire [0:0] v_5787;
  wire [0:0] v_5788;
  wire [0:0] v_5789;
  wire [0:0] vin0_consume_en_5790;
  wire [0:0] vout_canPeek_5790;
  wire [7:0] vout_peek_5790;
  wire [0:0] v_5791;
  wire [0:0] v_5792;
  function [0:0] mux_5792(input [0:0] sel);
    case (sel) 0: mux_5792 = 1'h0; 1: mux_5792 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5793;
  wire [0:0] v_5794;
  wire [0:0] v_5795;
  wire [0:0] v_5796;
  wire [0:0] v_5797;
  function [0:0] mux_5797(input [0:0] sel);
    case (sel) 0: mux_5797 = 1'h0; 1: mux_5797 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5798;
  wire [0:0] vin0_consume_en_5799;
  wire [0:0] vout_canPeek_5799;
  wire [7:0] vout_peek_5799;
  wire [0:0] v_5800;
  wire [0:0] v_5801;
  function [0:0] mux_5801(input [0:0] sel);
    case (sel) 0: mux_5801 = 1'h0; 1: mux_5801 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5802;
  function [0:0] mux_5802(input [0:0] sel);
    case (sel) 0: mux_5802 = 1'h0; 1: mux_5802 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5803;
  wire [0:0] v_5804;
  wire [0:0] v_5805;
  wire [0:0] v_5806;
  wire [0:0] v_5807;
  wire [0:0] v_5808;
  wire [0:0] v_5809;
  function [0:0] mux_5809(input [0:0] sel);
    case (sel) 0: mux_5809 = 1'h0; 1: mux_5809 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5810;
  function [0:0] mux_5810(input [0:0] sel);
    case (sel) 0: mux_5810 = 1'h0; 1: mux_5810 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5811;
  wire [0:0] v_5812;
  wire [0:0] v_5813;
  wire [0:0] v_5814;
  function [0:0] mux_5814(input [0:0] sel);
    case (sel) 0: mux_5814 = 1'h0; 1: mux_5814 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5815;
  function [0:0] mux_5815(input [0:0] sel);
    case (sel) 0: mux_5815 = 1'h0; 1: mux_5815 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5816;
  wire [0:0] v_5817;
  wire [0:0] v_5818;
  wire [0:0] v_5819;
  wire [0:0] v_5820;
  wire [0:0] v_5821;
  function [0:0] mux_5821(input [0:0] sel);
    case (sel) 0: mux_5821 = 1'h0; 1: mux_5821 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5822;
  wire [0:0] v_5823;
  wire [0:0] v_5824;
  wire [0:0] v_5825;
  wire [0:0] v_5826;
  function [0:0] mux_5826(input [0:0] sel);
    case (sel) 0: mux_5826 = 1'h0; 1: mux_5826 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5827;
  wire [0:0] v_5828;
  wire [0:0] v_5829;
  wire [0:0] v_5830;
  function [0:0] mux_5830(input [0:0] sel);
    case (sel) 0: mux_5830 = 1'h0; 1: mux_5830 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5831;
  function [0:0] mux_5831(input [0:0] sel);
    case (sel) 0: mux_5831 = 1'h0; 1: mux_5831 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5832 = 1'h0;
  wire [0:0] v_5833;
  wire [0:0] v_5834;
  wire [0:0] act_5835;
  wire [0:0] v_5836;
  wire [0:0] v_5837;
  wire [0:0] v_5838;
  reg [0:0] v_5839 = 1'h0;
  wire [0:0] v_5840;
  wire [0:0] v_5841;
  wire [0:0] act_5842;
  wire [0:0] v_5843;
  wire [0:0] v_5844;
  wire [0:0] v_5845;
  wire [0:0] vin0_consume_en_5846;
  wire [0:0] vout_canPeek_5846;
  wire [7:0] vout_peek_5846;
  wire [0:0] v_5847;
  wire [0:0] v_5848;
  function [0:0] mux_5848(input [0:0] sel);
    case (sel) 0: mux_5848 = 1'h0; 1: mux_5848 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5849;
  wire [0:0] v_5850;
  wire [0:0] v_5851;
  wire [0:0] v_5852;
  wire [0:0] v_5853;
  function [0:0] mux_5853(input [0:0] sel);
    case (sel) 0: mux_5853 = 1'h0; 1: mux_5853 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5854;
  wire [0:0] vin0_consume_en_5855;
  wire [0:0] vout_canPeek_5855;
  wire [7:0] vout_peek_5855;
  wire [0:0] v_5856;
  wire [0:0] v_5857;
  function [0:0] mux_5857(input [0:0] sel);
    case (sel) 0: mux_5857 = 1'h0; 1: mux_5857 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5858;
  function [0:0] mux_5858(input [0:0] sel);
    case (sel) 0: mux_5858 = 1'h0; 1: mux_5858 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5859;
  wire [0:0] v_5860;
  wire [0:0] v_5861;
  wire [0:0] v_5862;
  wire [0:0] v_5863;
  wire [0:0] v_5864;
  wire [0:0] v_5865;
  function [0:0] mux_5865(input [0:0] sel);
    case (sel) 0: mux_5865 = 1'h0; 1: mux_5865 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5866;
  wire [0:0] v_5867;
  wire [0:0] v_5868;
  wire [0:0] v_5869;
  wire [0:0] v_5870;
  function [0:0] mux_5870(input [0:0] sel);
    case (sel) 0: mux_5870 = 1'h0; 1: mux_5870 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5871;
  wire [0:0] v_5872;
  wire [0:0] v_5873;
  wire [0:0] v_5874;
  function [0:0] mux_5874(input [0:0] sel);
    case (sel) 0: mux_5874 = 1'h0; 1: mux_5874 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5875;
  function [0:0] mux_5875(input [0:0] sel);
    case (sel) 0: mux_5875 = 1'h0; 1: mux_5875 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5876 = 1'h0;
  wire [0:0] v_5877;
  wire [0:0] v_5878;
  wire [0:0] act_5879;
  wire [0:0] v_5880;
  wire [0:0] v_5881;
  wire [0:0] v_5882;
  wire [0:0] vin0_consume_en_5883;
  wire [0:0] vout_canPeek_5883;
  wire [7:0] vout_peek_5883;
  wire [0:0] v_5884;
  wire [0:0] v_5885;
  function [0:0] mux_5885(input [0:0] sel);
    case (sel) 0: mux_5885 = 1'h0; 1: mux_5885 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5886;
  wire [0:0] v_5887;
  wire [0:0] v_5888;
  wire [0:0] v_5889;
  wire [0:0] v_5890;
  function [0:0] mux_5890(input [0:0] sel);
    case (sel) 0: mux_5890 = 1'h0; 1: mux_5890 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5891;
  wire [0:0] vin0_consume_en_5892;
  wire [0:0] vout_canPeek_5892;
  wire [7:0] vout_peek_5892;
  wire [0:0] v_5893;
  wire [0:0] v_5894;
  function [0:0] mux_5894(input [0:0] sel);
    case (sel) 0: mux_5894 = 1'h0; 1: mux_5894 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5895;
  function [0:0] mux_5895(input [0:0] sel);
    case (sel) 0: mux_5895 = 1'h0; 1: mux_5895 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5896;
  wire [0:0] v_5897;
  wire [0:0] v_5898;
  wire [0:0] v_5899;
  wire [0:0] v_5900;
  wire [0:0] v_5901;
  wire [0:0] v_5902;
  function [0:0] mux_5902(input [0:0] sel);
    case (sel) 0: mux_5902 = 1'h0; 1: mux_5902 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5903;
  function [0:0] mux_5903(input [0:0] sel);
    case (sel) 0: mux_5903 = 1'h0; 1: mux_5903 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5904;
  wire [0:0] v_5905;
  wire [0:0] v_5906;
  wire [0:0] v_5907;
  function [0:0] mux_5907(input [0:0] sel);
    case (sel) 0: mux_5907 = 1'h0; 1: mux_5907 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5908;
  function [0:0] mux_5908(input [0:0] sel);
    case (sel) 0: mux_5908 = 1'h0; 1: mux_5908 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5909;
  wire [0:0] v_5910;
  wire [0:0] v_5911;
  wire [0:0] v_5912;
  wire [0:0] v_5913;
  wire [0:0] v_5914;
  function [0:0] mux_5914(input [0:0] sel);
    case (sel) 0: mux_5914 = 1'h0; 1: mux_5914 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5915;
  function [0:0] mux_5915(input [0:0] sel);
    case (sel) 0: mux_5915 = 1'h0; 1: mux_5915 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5916;
  wire [0:0] v_5917;
  wire [0:0] v_5918;
  wire [0:0] v_5919;
  function [0:0] mux_5919(input [0:0] sel);
    case (sel) 0: mux_5919 = 1'h0; 1: mux_5919 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5920;
  function [0:0] mux_5920(input [0:0] sel);
    case (sel) 0: mux_5920 = 1'h0; 1: mux_5920 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5921;
  wire [0:0] v_5922;
  wire [0:0] v_5923;
  wire [0:0] v_5924;
  wire [0:0] v_5925;
  wire [0:0] v_5926;
  function [0:0] mux_5926(input [0:0] sel);
    case (sel) 0: mux_5926 = 1'h0; 1: mux_5926 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5927;
  wire [0:0] v_5928;
  wire [0:0] v_5929;
  wire [0:0] v_5930;
  wire [0:0] v_5931;
  function [0:0] mux_5931(input [0:0] sel);
    case (sel) 0: mux_5931 = 1'h0; 1: mux_5931 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5932;
  wire [0:0] v_5933;
  wire [0:0] v_5934;
  wire [0:0] v_5935;
  function [0:0] mux_5935(input [0:0] sel);
    case (sel) 0: mux_5935 = 1'h0; 1: mux_5935 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5936;
  function [0:0] mux_5936(input [0:0] sel);
    case (sel) 0: mux_5936 = 1'h0; 1: mux_5936 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5937 = 1'h0;
  wire [0:0] v_5938;
  wire [0:0] v_5939;
  wire [0:0] act_5940;
  wire [0:0] v_5941;
  wire [0:0] v_5942;
  wire [0:0] v_5943;
  reg [0:0] v_5944 = 1'h0;
  wire [0:0] v_5945;
  wire [0:0] v_5946;
  wire [0:0] act_5947;
  wire [0:0] v_5948;
  wire [0:0] v_5949;
  wire [0:0] v_5950;
  reg [0:0] v_5951 = 1'h0;
  wire [0:0] v_5952;
  wire [0:0] v_5953;
  wire [0:0] act_5954;
  wire [0:0] v_5955;
  wire [0:0] v_5956;
  wire [0:0] v_5957;
  wire [0:0] vin0_consume_en_5958;
  wire [0:0] vout_canPeek_5958;
  wire [7:0] vout_peek_5958;
  wire [0:0] v_5959;
  wire [0:0] v_5960;
  function [0:0] mux_5960(input [0:0] sel);
    case (sel) 0: mux_5960 = 1'h0; 1: mux_5960 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5961;
  wire [0:0] v_5962;
  wire [0:0] v_5963;
  wire [0:0] v_5964;
  wire [0:0] v_5965;
  function [0:0] mux_5965(input [0:0] sel);
    case (sel) 0: mux_5965 = 1'h0; 1: mux_5965 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5966;
  wire [0:0] vin0_consume_en_5967;
  wire [0:0] vout_canPeek_5967;
  wire [7:0] vout_peek_5967;
  wire [0:0] v_5968;
  wire [0:0] v_5969;
  function [0:0] mux_5969(input [0:0] sel);
    case (sel) 0: mux_5969 = 1'h0; 1: mux_5969 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5970;
  function [0:0] mux_5970(input [0:0] sel);
    case (sel) 0: mux_5970 = 1'h0; 1: mux_5970 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5971;
  wire [0:0] v_5972;
  wire [0:0] v_5973;
  wire [0:0] v_5974;
  wire [0:0] v_5975;
  wire [0:0] v_5976;
  wire [0:0] v_5977;
  function [0:0] mux_5977(input [0:0] sel);
    case (sel) 0: mux_5977 = 1'h0; 1: mux_5977 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5978;
  wire [0:0] v_5979;
  wire [0:0] v_5980;
  wire [0:0] v_5981;
  wire [0:0] v_5982;
  function [0:0] mux_5982(input [0:0] sel);
    case (sel) 0: mux_5982 = 1'h0; 1: mux_5982 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5983;
  wire [0:0] v_5984;
  wire [0:0] v_5985;
  wire [0:0] v_5986;
  function [0:0] mux_5986(input [0:0] sel);
    case (sel) 0: mux_5986 = 1'h0; 1: mux_5986 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5987;
  function [0:0] mux_5987(input [0:0] sel);
    case (sel) 0: mux_5987 = 1'h0; 1: mux_5987 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5988 = 1'h0;
  wire [0:0] v_5989;
  wire [0:0] v_5990;
  wire [0:0] act_5991;
  wire [0:0] v_5992;
  wire [0:0] v_5993;
  wire [0:0] v_5994;
  wire [0:0] vin0_consume_en_5995;
  wire [0:0] vout_canPeek_5995;
  wire [7:0] vout_peek_5995;
  wire [0:0] v_5996;
  wire [0:0] v_5997;
  function [0:0] mux_5997(input [0:0] sel);
    case (sel) 0: mux_5997 = 1'h0; 1: mux_5997 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5998;
  wire [0:0] v_5999;
  wire [0:0] v_6000;
  wire [0:0] v_6001;
  wire [0:0] v_6002;
  function [0:0] mux_6002(input [0:0] sel);
    case (sel) 0: mux_6002 = 1'h0; 1: mux_6002 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6003;
  wire [0:0] vin0_consume_en_6004;
  wire [0:0] vout_canPeek_6004;
  wire [7:0] vout_peek_6004;
  wire [0:0] v_6005;
  wire [0:0] v_6006;
  function [0:0] mux_6006(input [0:0] sel);
    case (sel) 0: mux_6006 = 1'h0; 1: mux_6006 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6007;
  function [0:0] mux_6007(input [0:0] sel);
    case (sel) 0: mux_6007 = 1'h0; 1: mux_6007 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6008;
  wire [0:0] v_6009;
  wire [0:0] v_6010;
  wire [0:0] v_6011;
  wire [0:0] v_6012;
  wire [0:0] v_6013;
  wire [0:0] v_6014;
  function [0:0] mux_6014(input [0:0] sel);
    case (sel) 0: mux_6014 = 1'h0; 1: mux_6014 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6015;
  function [0:0] mux_6015(input [0:0] sel);
    case (sel) 0: mux_6015 = 1'h0; 1: mux_6015 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6016;
  wire [0:0] v_6017;
  wire [0:0] v_6018;
  wire [0:0] v_6019;
  function [0:0] mux_6019(input [0:0] sel);
    case (sel) 0: mux_6019 = 1'h0; 1: mux_6019 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6020;
  function [0:0] mux_6020(input [0:0] sel);
    case (sel) 0: mux_6020 = 1'h0; 1: mux_6020 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6021;
  wire [0:0] v_6022;
  wire [0:0] v_6023;
  wire [0:0] v_6024;
  wire [0:0] v_6025;
  wire [0:0] v_6026;
  function [0:0] mux_6026(input [0:0] sel);
    case (sel) 0: mux_6026 = 1'h0; 1: mux_6026 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6027;
  wire [0:0] v_6028;
  wire [0:0] v_6029;
  wire [0:0] v_6030;
  wire [0:0] v_6031;
  function [0:0] mux_6031(input [0:0] sel);
    case (sel) 0: mux_6031 = 1'h0; 1: mux_6031 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6032;
  wire [0:0] v_6033;
  wire [0:0] v_6034;
  wire [0:0] v_6035;
  function [0:0] mux_6035(input [0:0] sel);
    case (sel) 0: mux_6035 = 1'h0; 1: mux_6035 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6036;
  function [0:0] mux_6036(input [0:0] sel);
    case (sel) 0: mux_6036 = 1'h0; 1: mux_6036 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6037 = 1'h0;
  wire [0:0] v_6038;
  wire [0:0] v_6039;
  wire [0:0] act_6040;
  wire [0:0] v_6041;
  wire [0:0] v_6042;
  wire [0:0] v_6043;
  reg [0:0] v_6044 = 1'h0;
  wire [0:0] v_6045;
  wire [0:0] v_6046;
  wire [0:0] act_6047;
  wire [0:0] v_6048;
  wire [0:0] v_6049;
  wire [0:0] v_6050;
  wire [0:0] vin0_consume_en_6051;
  wire [0:0] vout_canPeek_6051;
  wire [7:0] vout_peek_6051;
  wire [0:0] v_6052;
  wire [0:0] v_6053;
  function [0:0] mux_6053(input [0:0] sel);
    case (sel) 0: mux_6053 = 1'h0; 1: mux_6053 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6054;
  wire [0:0] v_6055;
  wire [0:0] v_6056;
  wire [0:0] v_6057;
  wire [0:0] v_6058;
  function [0:0] mux_6058(input [0:0] sel);
    case (sel) 0: mux_6058 = 1'h0; 1: mux_6058 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6059;
  wire [0:0] vin0_consume_en_6060;
  wire [0:0] vout_canPeek_6060;
  wire [7:0] vout_peek_6060;
  wire [0:0] v_6061;
  wire [0:0] v_6062;
  function [0:0] mux_6062(input [0:0] sel);
    case (sel) 0: mux_6062 = 1'h0; 1: mux_6062 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6063;
  function [0:0] mux_6063(input [0:0] sel);
    case (sel) 0: mux_6063 = 1'h0; 1: mux_6063 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6064;
  wire [0:0] v_6065;
  wire [0:0] v_6066;
  wire [0:0] v_6067;
  wire [0:0] v_6068;
  wire [0:0] v_6069;
  wire [0:0] v_6070;
  function [0:0] mux_6070(input [0:0] sel);
    case (sel) 0: mux_6070 = 1'h0; 1: mux_6070 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6071;
  wire [0:0] v_6072;
  wire [0:0] v_6073;
  wire [0:0] v_6074;
  wire [0:0] v_6075;
  function [0:0] mux_6075(input [0:0] sel);
    case (sel) 0: mux_6075 = 1'h0; 1: mux_6075 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6076;
  wire [0:0] v_6077;
  wire [0:0] v_6078;
  wire [0:0] v_6079;
  function [0:0] mux_6079(input [0:0] sel);
    case (sel) 0: mux_6079 = 1'h0; 1: mux_6079 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6080;
  function [0:0] mux_6080(input [0:0] sel);
    case (sel) 0: mux_6080 = 1'h0; 1: mux_6080 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6081 = 1'h0;
  wire [0:0] v_6082;
  wire [0:0] v_6083;
  wire [0:0] act_6084;
  wire [0:0] v_6085;
  wire [0:0] v_6086;
  wire [0:0] v_6087;
  wire [0:0] vin0_consume_en_6088;
  wire [0:0] vout_canPeek_6088;
  wire [7:0] vout_peek_6088;
  wire [0:0] v_6089;
  wire [0:0] v_6090;
  function [0:0] mux_6090(input [0:0] sel);
    case (sel) 0: mux_6090 = 1'h0; 1: mux_6090 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6091;
  wire [0:0] v_6092;
  wire [0:0] v_6093;
  wire [0:0] v_6094;
  wire [0:0] v_6095;
  function [0:0] mux_6095(input [0:0] sel);
    case (sel) 0: mux_6095 = 1'h0; 1: mux_6095 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6096;
  wire [0:0] vin0_consume_en_6097;
  wire [0:0] vout_canPeek_6097;
  wire [7:0] vout_peek_6097;
  wire [0:0] v_6098;
  wire [0:0] v_6099;
  function [0:0] mux_6099(input [0:0] sel);
    case (sel) 0: mux_6099 = 1'h0; 1: mux_6099 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6100;
  function [0:0] mux_6100(input [0:0] sel);
    case (sel) 0: mux_6100 = 1'h0; 1: mux_6100 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6101;
  wire [0:0] v_6102;
  wire [0:0] v_6103;
  wire [0:0] v_6104;
  wire [0:0] v_6105;
  wire [0:0] v_6106;
  wire [0:0] v_6107;
  function [0:0] mux_6107(input [0:0] sel);
    case (sel) 0: mux_6107 = 1'h0; 1: mux_6107 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6108;
  function [0:0] mux_6108(input [0:0] sel);
    case (sel) 0: mux_6108 = 1'h0; 1: mux_6108 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6109;
  wire [0:0] v_6110;
  wire [0:0] v_6111;
  wire [0:0] v_6112;
  function [0:0] mux_6112(input [0:0] sel);
    case (sel) 0: mux_6112 = 1'h0; 1: mux_6112 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6113;
  function [0:0] mux_6113(input [0:0] sel);
    case (sel) 0: mux_6113 = 1'h0; 1: mux_6113 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6114;
  wire [0:0] v_6115;
  wire [0:0] v_6116;
  wire [0:0] v_6117;
  wire [0:0] v_6118;
  wire [0:0] v_6119;
  function [0:0] mux_6119(input [0:0] sel);
    case (sel) 0: mux_6119 = 1'h0; 1: mux_6119 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6120;
  function [0:0] mux_6120(input [0:0] sel);
    case (sel) 0: mux_6120 = 1'h0; 1: mux_6120 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6121;
  wire [0:0] v_6122;
  wire [0:0] v_6123;
  wire [0:0] v_6124;
  function [0:0] mux_6124(input [0:0] sel);
    case (sel) 0: mux_6124 = 1'h0; 1: mux_6124 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6125;
  function [0:0] mux_6125(input [0:0] sel);
    case (sel) 0: mux_6125 = 1'h0; 1: mux_6125 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6126;
  wire [0:0] v_6127;
  wire [0:0] v_6128;
  wire [0:0] v_6129;
  wire [0:0] v_6130;
  wire [0:0] v_6131;
  function [0:0] mux_6131(input [0:0] sel);
    case (sel) 0: mux_6131 = 1'h0; 1: mux_6131 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6132;
  function [0:0] mux_6132(input [0:0] sel);
    case (sel) 0: mux_6132 = 1'h0; 1: mux_6132 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6133;
  wire [0:0] v_6134;
  wire [0:0] v_6135;
  wire [0:0] v_6136;
  function [0:0] mux_6136(input [0:0] sel);
    case (sel) 0: mux_6136 = 1'h0; 1: mux_6136 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6137;
  function [0:0] mux_6137(input [0:0] sel);
    case (sel) 0: mux_6137 = 1'h0; 1: mux_6137 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6138;
  wire [0:0] v_6139;
  wire [0:0] v_6140;
  wire [0:0] v_6141;
  wire [0:0] v_6142;
  wire [0:0] v_6143;
  function [0:0] mux_6143(input [0:0] sel);
    case (sel) 0: mux_6143 = 1'h0; 1: mux_6143 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6144;
  function [0:0] mux_6144(input [0:0] sel);
    case (sel) 0: mux_6144 = 1'h0; 1: mux_6144 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6145;
  wire [0:0] v_6146;
  wire [0:0] v_6147;
  wire [0:0] v_6148;
  function [0:0] mux_6148(input [0:0] sel);
    case (sel) 0: mux_6148 = 1'h0; 1: mux_6148 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6149;
  function [0:0] mux_6149(input [0:0] sel);
    case (sel) 0: mux_6149 = 1'h0; 1: mux_6149 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6150;
  wire [0:0] v_6151;
  wire [0:0] v_6152;
  wire [0:0] v_6153;
  wire [0:0] v_6154;
  wire [0:0] v_6155;
  function [0:0] mux_6155(input [0:0] sel);
    case (sel) 0: mux_6155 = 1'h0; 1: mux_6155 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6156;
  function [0:0] mux_6156(input [0:0] sel);
    case (sel) 0: mux_6156 = 1'h0; 1: mux_6156 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6157;
  wire [0:0] v_6158;
  wire [0:0] v_6159;
  wire [0:0] v_6160;
  function [0:0] mux_6160(input [0:0] sel);
    case (sel) 0: mux_6160 = 1'h0; 1: mux_6160 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6161;
  function [0:0] mux_6161(input [0:0] sel);
    case (sel) 0: mux_6161 = 1'h0; 1: mux_6161 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6162;
  wire [0:0] v_6163;
  wire [0:0] v_6164;
  wire [0:0] v_6165;
  wire [0:0] v_6166;
  wire [0:0] v_6167;
  function [0:0] mux_6167(input [0:0] sel);
    case (sel) 0: mux_6167 = 1'h0; 1: mux_6167 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6168;
  wire [0:0] v_6169;
  wire [0:0] v_6170;
  wire [0:0] v_6171;
  wire [0:0] v_6172;
  function [0:0] mux_6172(input [0:0] sel);
    case (sel) 0: mux_6172 = 1'h0; 1: mux_6172 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6173;
  wire [0:0] v_6174;
  wire [0:0] v_6175;
  wire [0:0] v_6176;
  function [0:0] mux_6176(input [0:0] sel);
    case (sel) 0: mux_6176 = 1'h0; 1: mux_6176 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6177;
  function [0:0] mux_6177(input [0:0] sel);
    case (sel) 0: mux_6177 = 1'h0; 1: mux_6177 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6178 = 1'h0;
  wire [0:0] v_6179;
  wire [0:0] v_6180;
  wire [0:0] act_6181;
  wire [0:0] v_6182;
  wire [0:0] v_6183;
  wire [0:0] v_6184;
  reg [0:0] v_6185 = 1'h0;
  wire [0:0] v_6186;
  wire [0:0] v_6187;
  wire [0:0] act_6188;
  wire [0:0] v_6189;
  wire [0:0] v_6190;
  wire [0:0] v_6191;
  reg [0:0] v_6192 = 1'h0;
  wire [0:0] v_6193;
  wire [0:0] v_6194;
  wire [0:0] act_6195;
  wire [0:0] v_6196;
  wire [0:0] v_6197;
  wire [0:0] v_6198;
  reg [0:0] v_6199 = 1'h0;
  wire [0:0] v_6200;
  wire [0:0] v_6201;
  wire [0:0] act_6202;
  wire [0:0] v_6203;
  wire [0:0] v_6204;
  wire [0:0] v_6205;
  reg [0:0] v_6206 = 1'h0;
  wire [0:0] v_6207;
  wire [0:0] v_6208;
  wire [0:0] act_6209;
  wire [0:0] v_6210;
  wire [0:0] v_6211;
  wire [0:0] v_6212;
  reg [0:0] v_6213 = 1'h0;
  wire [0:0] v_6214;
  wire [0:0] v_6215;
  wire [0:0] act_6216;
  wire [0:0] v_6217;
  wire [0:0] v_6218;
  wire [0:0] v_6219;
  wire [0:0] vin0_consume_en_6220;
  wire [0:0] vout_canPeek_6220;
  wire [7:0] vout_peek_6220;
  wire [0:0] v_6221;
  wire [0:0] v_6222;
  function [0:0] mux_6222(input [0:0] sel);
    case (sel) 0: mux_6222 = 1'h0; 1: mux_6222 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6223;
  wire [0:0] v_6224;
  wire [0:0] v_6225;
  wire [0:0] v_6226;
  wire [0:0] v_6227;
  function [0:0] mux_6227(input [0:0] sel);
    case (sel) 0: mux_6227 = 1'h0; 1: mux_6227 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6228;
  wire [0:0] vin0_consume_en_6229;
  wire [0:0] vout_canPeek_6229;
  wire [7:0] vout_peek_6229;
  wire [0:0] v_6230;
  wire [0:0] v_6231;
  function [0:0] mux_6231(input [0:0] sel);
    case (sel) 0: mux_6231 = 1'h0; 1: mux_6231 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6232;
  function [0:0] mux_6232(input [0:0] sel);
    case (sel) 0: mux_6232 = 1'h0; 1: mux_6232 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6233;
  wire [0:0] v_6234;
  wire [0:0] v_6235;
  wire [0:0] v_6236;
  wire [0:0] v_6237;
  wire [0:0] v_6238;
  wire [0:0] v_6239;
  function [0:0] mux_6239(input [0:0] sel);
    case (sel) 0: mux_6239 = 1'h0; 1: mux_6239 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6240;
  wire [0:0] v_6241;
  wire [0:0] v_6242;
  wire [0:0] v_6243;
  wire [0:0] v_6244;
  function [0:0] mux_6244(input [0:0] sel);
    case (sel) 0: mux_6244 = 1'h0; 1: mux_6244 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6245;
  wire [0:0] v_6246;
  wire [0:0] v_6247;
  wire [0:0] v_6248;
  function [0:0] mux_6248(input [0:0] sel);
    case (sel) 0: mux_6248 = 1'h0; 1: mux_6248 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6249;
  function [0:0] mux_6249(input [0:0] sel);
    case (sel) 0: mux_6249 = 1'h0; 1: mux_6249 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6250 = 1'h0;
  wire [0:0] v_6251;
  wire [0:0] v_6252;
  wire [0:0] act_6253;
  wire [0:0] v_6254;
  wire [0:0] v_6255;
  wire [0:0] v_6256;
  wire [0:0] vin0_consume_en_6257;
  wire [0:0] vout_canPeek_6257;
  wire [7:0] vout_peek_6257;
  wire [0:0] v_6258;
  wire [0:0] v_6259;
  function [0:0] mux_6259(input [0:0] sel);
    case (sel) 0: mux_6259 = 1'h0; 1: mux_6259 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6260;
  wire [0:0] v_6261;
  wire [0:0] v_6262;
  wire [0:0] v_6263;
  wire [0:0] v_6264;
  function [0:0] mux_6264(input [0:0] sel);
    case (sel) 0: mux_6264 = 1'h0; 1: mux_6264 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6265;
  wire [0:0] vin0_consume_en_6266;
  wire [0:0] vout_canPeek_6266;
  wire [7:0] vout_peek_6266;
  wire [0:0] v_6267;
  wire [0:0] v_6268;
  function [0:0] mux_6268(input [0:0] sel);
    case (sel) 0: mux_6268 = 1'h0; 1: mux_6268 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6269;
  function [0:0] mux_6269(input [0:0] sel);
    case (sel) 0: mux_6269 = 1'h0; 1: mux_6269 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6270;
  wire [0:0] v_6271;
  wire [0:0] v_6272;
  wire [0:0] v_6273;
  wire [0:0] v_6274;
  wire [0:0] v_6275;
  wire [0:0] v_6276;
  function [0:0] mux_6276(input [0:0] sel);
    case (sel) 0: mux_6276 = 1'h0; 1: mux_6276 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6277;
  function [0:0] mux_6277(input [0:0] sel);
    case (sel) 0: mux_6277 = 1'h0; 1: mux_6277 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6278;
  wire [0:0] v_6279;
  wire [0:0] v_6280;
  wire [0:0] v_6281;
  function [0:0] mux_6281(input [0:0] sel);
    case (sel) 0: mux_6281 = 1'h0; 1: mux_6281 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6282;
  function [0:0] mux_6282(input [0:0] sel);
    case (sel) 0: mux_6282 = 1'h0; 1: mux_6282 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6283;
  wire [0:0] v_6284;
  wire [0:0] v_6285;
  wire [0:0] v_6286;
  wire [0:0] v_6287;
  wire [0:0] v_6288;
  function [0:0] mux_6288(input [0:0] sel);
    case (sel) 0: mux_6288 = 1'h0; 1: mux_6288 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6289;
  wire [0:0] v_6290;
  wire [0:0] v_6291;
  wire [0:0] v_6292;
  wire [0:0] v_6293;
  function [0:0] mux_6293(input [0:0] sel);
    case (sel) 0: mux_6293 = 1'h0; 1: mux_6293 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6294;
  wire [0:0] v_6295;
  wire [0:0] v_6296;
  wire [0:0] v_6297;
  function [0:0] mux_6297(input [0:0] sel);
    case (sel) 0: mux_6297 = 1'h0; 1: mux_6297 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6298;
  function [0:0] mux_6298(input [0:0] sel);
    case (sel) 0: mux_6298 = 1'h0; 1: mux_6298 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6299 = 1'h0;
  wire [0:0] v_6300;
  wire [0:0] v_6301;
  wire [0:0] act_6302;
  wire [0:0] v_6303;
  wire [0:0] v_6304;
  wire [0:0] v_6305;
  reg [0:0] v_6306 = 1'h0;
  wire [0:0] v_6307;
  wire [0:0] v_6308;
  wire [0:0] act_6309;
  wire [0:0] v_6310;
  wire [0:0] v_6311;
  wire [0:0] v_6312;
  wire [0:0] vin0_consume_en_6313;
  wire [0:0] vout_canPeek_6313;
  wire [7:0] vout_peek_6313;
  wire [0:0] v_6314;
  wire [0:0] v_6315;
  function [0:0] mux_6315(input [0:0] sel);
    case (sel) 0: mux_6315 = 1'h0; 1: mux_6315 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6316;
  wire [0:0] v_6317;
  wire [0:0] v_6318;
  wire [0:0] v_6319;
  wire [0:0] v_6320;
  function [0:0] mux_6320(input [0:0] sel);
    case (sel) 0: mux_6320 = 1'h0; 1: mux_6320 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6321;
  wire [0:0] vin0_consume_en_6322;
  wire [0:0] vout_canPeek_6322;
  wire [7:0] vout_peek_6322;
  wire [0:0] v_6323;
  wire [0:0] v_6324;
  function [0:0] mux_6324(input [0:0] sel);
    case (sel) 0: mux_6324 = 1'h0; 1: mux_6324 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6325;
  function [0:0] mux_6325(input [0:0] sel);
    case (sel) 0: mux_6325 = 1'h0; 1: mux_6325 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6326;
  wire [0:0] v_6327;
  wire [0:0] v_6328;
  wire [0:0] v_6329;
  wire [0:0] v_6330;
  wire [0:0] v_6331;
  wire [0:0] v_6332;
  function [0:0] mux_6332(input [0:0] sel);
    case (sel) 0: mux_6332 = 1'h0; 1: mux_6332 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6333;
  wire [0:0] v_6334;
  wire [0:0] v_6335;
  wire [0:0] v_6336;
  wire [0:0] v_6337;
  function [0:0] mux_6337(input [0:0] sel);
    case (sel) 0: mux_6337 = 1'h0; 1: mux_6337 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6338;
  wire [0:0] v_6339;
  wire [0:0] v_6340;
  wire [0:0] v_6341;
  function [0:0] mux_6341(input [0:0] sel);
    case (sel) 0: mux_6341 = 1'h0; 1: mux_6341 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6342;
  function [0:0] mux_6342(input [0:0] sel);
    case (sel) 0: mux_6342 = 1'h0; 1: mux_6342 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6343 = 1'h0;
  wire [0:0] v_6344;
  wire [0:0] v_6345;
  wire [0:0] act_6346;
  wire [0:0] v_6347;
  wire [0:0] v_6348;
  wire [0:0] v_6349;
  wire [0:0] vin0_consume_en_6350;
  wire [0:0] vout_canPeek_6350;
  wire [7:0] vout_peek_6350;
  wire [0:0] v_6351;
  wire [0:0] v_6352;
  function [0:0] mux_6352(input [0:0] sel);
    case (sel) 0: mux_6352 = 1'h0; 1: mux_6352 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6353;
  wire [0:0] v_6354;
  wire [0:0] v_6355;
  wire [0:0] v_6356;
  wire [0:0] v_6357;
  function [0:0] mux_6357(input [0:0] sel);
    case (sel) 0: mux_6357 = 1'h0; 1: mux_6357 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6358;
  wire [0:0] vin0_consume_en_6359;
  wire [0:0] vout_canPeek_6359;
  wire [7:0] vout_peek_6359;
  wire [0:0] v_6360;
  wire [0:0] v_6361;
  function [0:0] mux_6361(input [0:0] sel);
    case (sel) 0: mux_6361 = 1'h0; 1: mux_6361 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6362;
  function [0:0] mux_6362(input [0:0] sel);
    case (sel) 0: mux_6362 = 1'h0; 1: mux_6362 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6363;
  wire [0:0] v_6364;
  wire [0:0] v_6365;
  wire [0:0] v_6366;
  wire [0:0] v_6367;
  wire [0:0] v_6368;
  wire [0:0] v_6369;
  function [0:0] mux_6369(input [0:0] sel);
    case (sel) 0: mux_6369 = 1'h0; 1: mux_6369 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6370;
  function [0:0] mux_6370(input [0:0] sel);
    case (sel) 0: mux_6370 = 1'h0; 1: mux_6370 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6371;
  wire [0:0] v_6372;
  wire [0:0] v_6373;
  wire [0:0] v_6374;
  function [0:0] mux_6374(input [0:0] sel);
    case (sel) 0: mux_6374 = 1'h0; 1: mux_6374 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6375;
  function [0:0] mux_6375(input [0:0] sel);
    case (sel) 0: mux_6375 = 1'h0; 1: mux_6375 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6376;
  wire [0:0] v_6377;
  wire [0:0] v_6378;
  wire [0:0] v_6379;
  wire [0:0] v_6380;
  wire [0:0] v_6381;
  function [0:0] mux_6381(input [0:0] sel);
    case (sel) 0: mux_6381 = 1'h0; 1: mux_6381 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6382;
  function [0:0] mux_6382(input [0:0] sel);
    case (sel) 0: mux_6382 = 1'h0; 1: mux_6382 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6383;
  wire [0:0] v_6384;
  wire [0:0] v_6385;
  wire [0:0] v_6386;
  function [0:0] mux_6386(input [0:0] sel);
    case (sel) 0: mux_6386 = 1'h0; 1: mux_6386 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6387;
  function [0:0] mux_6387(input [0:0] sel);
    case (sel) 0: mux_6387 = 1'h0; 1: mux_6387 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6388;
  wire [0:0] v_6389;
  wire [0:0] v_6390;
  wire [0:0] v_6391;
  wire [0:0] v_6392;
  wire [0:0] v_6393;
  function [0:0] mux_6393(input [0:0] sel);
    case (sel) 0: mux_6393 = 1'h0; 1: mux_6393 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6394;
  wire [0:0] v_6395;
  wire [0:0] v_6396;
  wire [0:0] v_6397;
  wire [0:0] v_6398;
  function [0:0] mux_6398(input [0:0] sel);
    case (sel) 0: mux_6398 = 1'h0; 1: mux_6398 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6399;
  wire [0:0] v_6400;
  wire [0:0] v_6401;
  wire [0:0] v_6402;
  function [0:0] mux_6402(input [0:0] sel);
    case (sel) 0: mux_6402 = 1'h0; 1: mux_6402 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6403;
  function [0:0] mux_6403(input [0:0] sel);
    case (sel) 0: mux_6403 = 1'h0; 1: mux_6403 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6404 = 1'h0;
  wire [0:0] v_6405;
  wire [0:0] v_6406;
  wire [0:0] act_6407;
  wire [0:0] v_6408;
  wire [0:0] v_6409;
  wire [0:0] v_6410;
  reg [0:0] v_6411 = 1'h0;
  wire [0:0] v_6412;
  wire [0:0] v_6413;
  wire [0:0] act_6414;
  wire [0:0] v_6415;
  wire [0:0] v_6416;
  wire [0:0] v_6417;
  reg [0:0] v_6418 = 1'h0;
  wire [0:0] v_6419;
  wire [0:0] v_6420;
  wire [0:0] act_6421;
  wire [0:0] v_6422;
  wire [0:0] v_6423;
  wire [0:0] v_6424;
  wire [0:0] vin0_consume_en_6425;
  wire [0:0] vout_canPeek_6425;
  wire [7:0] vout_peek_6425;
  wire [0:0] v_6426;
  wire [0:0] v_6427;
  function [0:0] mux_6427(input [0:0] sel);
    case (sel) 0: mux_6427 = 1'h0; 1: mux_6427 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6428;
  wire [0:0] v_6429;
  wire [0:0] v_6430;
  wire [0:0] v_6431;
  wire [0:0] v_6432;
  function [0:0] mux_6432(input [0:0] sel);
    case (sel) 0: mux_6432 = 1'h0; 1: mux_6432 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6433;
  wire [0:0] vin0_consume_en_6434;
  wire [0:0] vout_canPeek_6434;
  wire [7:0] vout_peek_6434;
  wire [0:0] v_6435;
  wire [0:0] v_6436;
  function [0:0] mux_6436(input [0:0] sel);
    case (sel) 0: mux_6436 = 1'h0; 1: mux_6436 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6437;
  function [0:0] mux_6437(input [0:0] sel);
    case (sel) 0: mux_6437 = 1'h0; 1: mux_6437 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6438;
  wire [0:0] v_6439;
  wire [0:0] v_6440;
  wire [0:0] v_6441;
  wire [0:0] v_6442;
  wire [0:0] v_6443;
  wire [0:0] v_6444;
  function [0:0] mux_6444(input [0:0] sel);
    case (sel) 0: mux_6444 = 1'h0; 1: mux_6444 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6445;
  wire [0:0] v_6446;
  wire [0:0] v_6447;
  wire [0:0] v_6448;
  wire [0:0] v_6449;
  function [0:0] mux_6449(input [0:0] sel);
    case (sel) 0: mux_6449 = 1'h0; 1: mux_6449 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6450;
  wire [0:0] v_6451;
  wire [0:0] v_6452;
  wire [0:0] v_6453;
  function [0:0] mux_6453(input [0:0] sel);
    case (sel) 0: mux_6453 = 1'h0; 1: mux_6453 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6454;
  function [0:0] mux_6454(input [0:0] sel);
    case (sel) 0: mux_6454 = 1'h0; 1: mux_6454 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6455 = 1'h0;
  wire [0:0] v_6456;
  wire [0:0] v_6457;
  wire [0:0] act_6458;
  wire [0:0] v_6459;
  wire [0:0] v_6460;
  wire [0:0] v_6461;
  wire [0:0] vin0_consume_en_6462;
  wire [0:0] vout_canPeek_6462;
  wire [7:0] vout_peek_6462;
  wire [0:0] v_6463;
  wire [0:0] v_6464;
  function [0:0] mux_6464(input [0:0] sel);
    case (sel) 0: mux_6464 = 1'h0; 1: mux_6464 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6465;
  wire [0:0] v_6466;
  wire [0:0] v_6467;
  wire [0:0] v_6468;
  wire [0:0] v_6469;
  function [0:0] mux_6469(input [0:0] sel);
    case (sel) 0: mux_6469 = 1'h0; 1: mux_6469 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6470;
  wire [0:0] vin0_consume_en_6471;
  wire [0:0] vout_canPeek_6471;
  wire [7:0] vout_peek_6471;
  wire [0:0] v_6472;
  wire [0:0] v_6473;
  function [0:0] mux_6473(input [0:0] sel);
    case (sel) 0: mux_6473 = 1'h0; 1: mux_6473 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6474;
  function [0:0] mux_6474(input [0:0] sel);
    case (sel) 0: mux_6474 = 1'h0; 1: mux_6474 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6475;
  wire [0:0] v_6476;
  wire [0:0] v_6477;
  wire [0:0] v_6478;
  wire [0:0] v_6479;
  wire [0:0] v_6480;
  wire [0:0] v_6481;
  function [0:0] mux_6481(input [0:0] sel);
    case (sel) 0: mux_6481 = 1'h0; 1: mux_6481 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6482;
  function [0:0] mux_6482(input [0:0] sel);
    case (sel) 0: mux_6482 = 1'h0; 1: mux_6482 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6483;
  wire [0:0] v_6484;
  wire [0:0] v_6485;
  wire [0:0] v_6486;
  function [0:0] mux_6486(input [0:0] sel);
    case (sel) 0: mux_6486 = 1'h0; 1: mux_6486 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6487;
  function [0:0] mux_6487(input [0:0] sel);
    case (sel) 0: mux_6487 = 1'h0; 1: mux_6487 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6488;
  wire [0:0] v_6489;
  wire [0:0] v_6490;
  wire [0:0] v_6491;
  wire [0:0] v_6492;
  wire [0:0] v_6493;
  function [0:0] mux_6493(input [0:0] sel);
    case (sel) 0: mux_6493 = 1'h0; 1: mux_6493 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6494;
  wire [0:0] v_6495;
  wire [0:0] v_6496;
  wire [0:0] v_6497;
  wire [0:0] v_6498;
  function [0:0] mux_6498(input [0:0] sel);
    case (sel) 0: mux_6498 = 1'h0; 1: mux_6498 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6499;
  wire [0:0] v_6500;
  wire [0:0] v_6501;
  wire [0:0] v_6502;
  function [0:0] mux_6502(input [0:0] sel);
    case (sel) 0: mux_6502 = 1'h0; 1: mux_6502 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6503;
  function [0:0] mux_6503(input [0:0] sel);
    case (sel) 0: mux_6503 = 1'h0; 1: mux_6503 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6504 = 1'h0;
  wire [0:0] v_6505;
  wire [0:0] v_6506;
  wire [0:0] act_6507;
  wire [0:0] v_6508;
  wire [0:0] v_6509;
  wire [0:0] v_6510;
  reg [0:0] v_6511 = 1'h0;
  wire [0:0] v_6512;
  wire [0:0] v_6513;
  wire [0:0] act_6514;
  wire [0:0] v_6515;
  wire [0:0] v_6516;
  wire [0:0] v_6517;
  wire [0:0] vin0_consume_en_6518;
  wire [0:0] vout_canPeek_6518;
  wire [7:0] vout_peek_6518;
  wire [0:0] v_6519;
  wire [0:0] v_6520;
  function [0:0] mux_6520(input [0:0] sel);
    case (sel) 0: mux_6520 = 1'h0; 1: mux_6520 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6521;
  wire [0:0] v_6522;
  wire [0:0] v_6523;
  wire [0:0] v_6524;
  wire [0:0] v_6525;
  function [0:0] mux_6525(input [0:0] sel);
    case (sel) 0: mux_6525 = 1'h0; 1: mux_6525 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6526;
  wire [0:0] vin0_consume_en_6527;
  wire [0:0] vout_canPeek_6527;
  wire [7:0] vout_peek_6527;
  wire [0:0] v_6528;
  wire [0:0] v_6529;
  function [0:0] mux_6529(input [0:0] sel);
    case (sel) 0: mux_6529 = 1'h0; 1: mux_6529 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6530;
  function [0:0] mux_6530(input [0:0] sel);
    case (sel) 0: mux_6530 = 1'h0; 1: mux_6530 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6531;
  wire [0:0] v_6532;
  wire [0:0] v_6533;
  wire [0:0] v_6534;
  wire [0:0] v_6535;
  wire [0:0] v_6536;
  wire [0:0] v_6537;
  function [0:0] mux_6537(input [0:0] sel);
    case (sel) 0: mux_6537 = 1'h0; 1: mux_6537 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6538;
  wire [0:0] v_6539;
  wire [0:0] v_6540;
  wire [0:0] v_6541;
  wire [0:0] v_6542;
  function [0:0] mux_6542(input [0:0] sel);
    case (sel) 0: mux_6542 = 1'h0; 1: mux_6542 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6543;
  wire [0:0] v_6544;
  wire [0:0] v_6545;
  wire [0:0] v_6546;
  function [0:0] mux_6546(input [0:0] sel);
    case (sel) 0: mux_6546 = 1'h0; 1: mux_6546 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6547;
  function [0:0] mux_6547(input [0:0] sel);
    case (sel) 0: mux_6547 = 1'h0; 1: mux_6547 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6548 = 1'h0;
  wire [0:0] v_6549;
  wire [0:0] v_6550;
  wire [0:0] act_6551;
  wire [0:0] v_6552;
  wire [0:0] v_6553;
  wire [0:0] v_6554;
  wire [0:0] vin0_consume_en_6555;
  wire [0:0] vout_canPeek_6555;
  wire [7:0] vout_peek_6555;
  wire [0:0] v_6556;
  wire [0:0] v_6557;
  function [0:0] mux_6557(input [0:0] sel);
    case (sel) 0: mux_6557 = 1'h0; 1: mux_6557 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6558;
  wire [0:0] v_6559;
  wire [0:0] v_6560;
  wire [0:0] v_6561;
  wire [0:0] v_6562;
  function [0:0] mux_6562(input [0:0] sel);
    case (sel) 0: mux_6562 = 1'h0; 1: mux_6562 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6563;
  wire [0:0] vin0_consume_en_6564;
  wire [0:0] vout_canPeek_6564;
  wire [7:0] vout_peek_6564;
  wire [0:0] v_6565;
  wire [0:0] v_6566;
  function [0:0] mux_6566(input [0:0] sel);
    case (sel) 0: mux_6566 = 1'h0; 1: mux_6566 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6567;
  function [0:0] mux_6567(input [0:0] sel);
    case (sel) 0: mux_6567 = 1'h0; 1: mux_6567 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6568;
  wire [0:0] v_6569;
  wire [0:0] v_6570;
  wire [0:0] v_6571;
  wire [0:0] v_6572;
  wire [0:0] v_6573;
  wire [0:0] v_6574;
  function [0:0] mux_6574(input [0:0] sel);
    case (sel) 0: mux_6574 = 1'h0; 1: mux_6574 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6575;
  function [0:0] mux_6575(input [0:0] sel);
    case (sel) 0: mux_6575 = 1'h0; 1: mux_6575 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6576;
  wire [0:0] v_6577;
  wire [0:0] v_6578;
  wire [0:0] v_6579;
  function [0:0] mux_6579(input [0:0] sel);
    case (sel) 0: mux_6579 = 1'h0; 1: mux_6579 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6580;
  function [0:0] mux_6580(input [0:0] sel);
    case (sel) 0: mux_6580 = 1'h0; 1: mux_6580 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6581;
  wire [0:0] v_6582;
  wire [0:0] v_6583;
  wire [0:0] v_6584;
  wire [0:0] v_6585;
  wire [0:0] v_6586;
  function [0:0] mux_6586(input [0:0] sel);
    case (sel) 0: mux_6586 = 1'h0; 1: mux_6586 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6587;
  function [0:0] mux_6587(input [0:0] sel);
    case (sel) 0: mux_6587 = 1'h0; 1: mux_6587 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6588;
  wire [0:0] v_6589;
  wire [0:0] v_6590;
  wire [0:0] v_6591;
  function [0:0] mux_6591(input [0:0] sel);
    case (sel) 0: mux_6591 = 1'h0; 1: mux_6591 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6592;
  function [0:0] mux_6592(input [0:0] sel);
    case (sel) 0: mux_6592 = 1'h0; 1: mux_6592 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6593;
  wire [0:0] v_6594;
  wire [0:0] v_6595;
  wire [0:0] v_6596;
  wire [0:0] v_6597;
  wire [0:0] v_6598;
  function [0:0] mux_6598(input [0:0] sel);
    case (sel) 0: mux_6598 = 1'h0; 1: mux_6598 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6599;
  function [0:0] mux_6599(input [0:0] sel);
    case (sel) 0: mux_6599 = 1'h0; 1: mux_6599 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6600;
  wire [0:0] v_6601;
  wire [0:0] v_6602;
  wire [0:0] v_6603;
  function [0:0] mux_6603(input [0:0] sel);
    case (sel) 0: mux_6603 = 1'h0; 1: mux_6603 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6604;
  function [0:0] mux_6604(input [0:0] sel);
    case (sel) 0: mux_6604 = 1'h0; 1: mux_6604 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6605;
  wire [0:0] v_6606;
  wire [0:0] v_6607;
  wire [0:0] v_6608;
  wire [0:0] v_6609;
  wire [0:0] v_6610;
  function [0:0] mux_6610(input [0:0] sel);
    case (sel) 0: mux_6610 = 1'h0; 1: mux_6610 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6611;
  wire [0:0] v_6612;
  wire [0:0] v_6613;
  wire [0:0] v_6614;
  wire [0:0] v_6615;
  function [0:0] mux_6615(input [0:0] sel);
    case (sel) 0: mux_6615 = 1'h0; 1: mux_6615 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6616;
  wire [0:0] v_6617;
  wire [0:0] v_6618;
  wire [0:0] v_6619;
  function [0:0] mux_6619(input [0:0] sel);
    case (sel) 0: mux_6619 = 1'h0; 1: mux_6619 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6620;
  function [0:0] mux_6620(input [0:0] sel);
    case (sel) 0: mux_6620 = 1'h0; 1: mux_6620 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6621 = 1'h0;
  wire [0:0] v_6622;
  wire [0:0] v_6623;
  wire [0:0] act_6624;
  wire [0:0] v_6625;
  wire [0:0] v_6626;
  wire [0:0] v_6627;
  reg [0:0] v_6628 = 1'h0;
  wire [0:0] v_6629;
  wire [0:0] v_6630;
  wire [0:0] act_6631;
  wire [0:0] v_6632;
  wire [0:0] v_6633;
  wire [0:0] v_6634;
  reg [0:0] v_6635 = 1'h0;
  wire [0:0] v_6636;
  wire [0:0] v_6637;
  wire [0:0] act_6638;
  wire [0:0] v_6639;
  wire [0:0] v_6640;
  wire [0:0] v_6641;
  reg [0:0] v_6642 = 1'h0;
  wire [0:0] v_6643;
  wire [0:0] v_6644;
  wire [0:0] act_6645;
  wire [0:0] v_6646;
  wire [0:0] v_6647;
  wire [0:0] v_6648;
  wire [0:0] vin0_consume_en_6649;
  wire [0:0] vout_canPeek_6649;
  wire [7:0] vout_peek_6649;
  wire [0:0] v_6650;
  wire [0:0] v_6651;
  function [0:0] mux_6651(input [0:0] sel);
    case (sel) 0: mux_6651 = 1'h0; 1: mux_6651 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6652;
  wire [0:0] v_6653;
  wire [0:0] v_6654;
  wire [0:0] v_6655;
  wire [0:0] v_6656;
  function [0:0] mux_6656(input [0:0] sel);
    case (sel) 0: mux_6656 = 1'h0; 1: mux_6656 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6657;
  wire [0:0] vin0_consume_en_6658;
  wire [0:0] vout_canPeek_6658;
  wire [7:0] vout_peek_6658;
  wire [0:0] v_6659;
  wire [0:0] v_6660;
  function [0:0] mux_6660(input [0:0] sel);
    case (sel) 0: mux_6660 = 1'h0; 1: mux_6660 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6661;
  function [0:0] mux_6661(input [0:0] sel);
    case (sel) 0: mux_6661 = 1'h0; 1: mux_6661 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6662;
  wire [0:0] v_6663;
  wire [0:0] v_6664;
  wire [0:0] v_6665;
  wire [0:0] v_6666;
  wire [0:0] v_6667;
  wire [0:0] v_6668;
  function [0:0] mux_6668(input [0:0] sel);
    case (sel) 0: mux_6668 = 1'h0; 1: mux_6668 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6669;
  wire [0:0] v_6670;
  wire [0:0] v_6671;
  wire [0:0] v_6672;
  wire [0:0] v_6673;
  function [0:0] mux_6673(input [0:0] sel);
    case (sel) 0: mux_6673 = 1'h0; 1: mux_6673 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6674;
  wire [0:0] v_6675;
  wire [0:0] v_6676;
  wire [0:0] v_6677;
  function [0:0] mux_6677(input [0:0] sel);
    case (sel) 0: mux_6677 = 1'h0; 1: mux_6677 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6678;
  function [0:0] mux_6678(input [0:0] sel);
    case (sel) 0: mux_6678 = 1'h0; 1: mux_6678 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6679 = 1'h0;
  wire [0:0] v_6680;
  wire [0:0] v_6681;
  wire [0:0] act_6682;
  wire [0:0] v_6683;
  wire [0:0] v_6684;
  wire [0:0] v_6685;
  wire [0:0] vin0_consume_en_6686;
  wire [0:0] vout_canPeek_6686;
  wire [7:0] vout_peek_6686;
  wire [0:0] v_6687;
  wire [0:0] v_6688;
  function [0:0] mux_6688(input [0:0] sel);
    case (sel) 0: mux_6688 = 1'h0; 1: mux_6688 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6689;
  wire [0:0] v_6690;
  wire [0:0] v_6691;
  wire [0:0] v_6692;
  wire [0:0] v_6693;
  function [0:0] mux_6693(input [0:0] sel);
    case (sel) 0: mux_6693 = 1'h0; 1: mux_6693 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6694;
  wire [0:0] vin0_consume_en_6695;
  wire [0:0] vout_canPeek_6695;
  wire [7:0] vout_peek_6695;
  wire [0:0] v_6696;
  wire [0:0] v_6697;
  function [0:0] mux_6697(input [0:0] sel);
    case (sel) 0: mux_6697 = 1'h0; 1: mux_6697 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6698;
  function [0:0] mux_6698(input [0:0] sel);
    case (sel) 0: mux_6698 = 1'h0; 1: mux_6698 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6699;
  wire [0:0] v_6700;
  wire [0:0] v_6701;
  wire [0:0] v_6702;
  wire [0:0] v_6703;
  wire [0:0] v_6704;
  wire [0:0] v_6705;
  function [0:0] mux_6705(input [0:0] sel);
    case (sel) 0: mux_6705 = 1'h0; 1: mux_6705 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6706;
  function [0:0] mux_6706(input [0:0] sel);
    case (sel) 0: mux_6706 = 1'h0; 1: mux_6706 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6707;
  wire [0:0] v_6708;
  wire [0:0] v_6709;
  wire [0:0] v_6710;
  function [0:0] mux_6710(input [0:0] sel);
    case (sel) 0: mux_6710 = 1'h0; 1: mux_6710 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6711;
  function [0:0] mux_6711(input [0:0] sel);
    case (sel) 0: mux_6711 = 1'h0; 1: mux_6711 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6712;
  wire [0:0] v_6713;
  wire [0:0] v_6714;
  wire [0:0] v_6715;
  wire [0:0] v_6716;
  wire [0:0] v_6717;
  function [0:0] mux_6717(input [0:0] sel);
    case (sel) 0: mux_6717 = 1'h0; 1: mux_6717 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6718;
  wire [0:0] v_6719;
  wire [0:0] v_6720;
  wire [0:0] v_6721;
  wire [0:0] v_6722;
  function [0:0] mux_6722(input [0:0] sel);
    case (sel) 0: mux_6722 = 1'h0; 1: mux_6722 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6723;
  wire [0:0] v_6724;
  wire [0:0] v_6725;
  wire [0:0] v_6726;
  function [0:0] mux_6726(input [0:0] sel);
    case (sel) 0: mux_6726 = 1'h0; 1: mux_6726 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6727;
  function [0:0] mux_6727(input [0:0] sel);
    case (sel) 0: mux_6727 = 1'h0; 1: mux_6727 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6728 = 1'h0;
  wire [0:0] v_6729;
  wire [0:0] v_6730;
  wire [0:0] act_6731;
  wire [0:0] v_6732;
  wire [0:0] v_6733;
  wire [0:0] v_6734;
  reg [0:0] v_6735 = 1'h0;
  wire [0:0] v_6736;
  wire [0:0] v_6737;
  wire [0:0] act_6738;
  wire [0:0] v_6739;
  wire [0:0] v_6740;
  wire [0:0] v_6741;
  wire [0:0] vin0_consume_en_6742;
  wire [0:0] vout_canPeek_6742;
  wire [7:0] vout_peek_6742;
  wire [0:0] v_6743;
  wire [0:0] v_6744;
  function [0:0] mux_6744(input [0:0] sel);
    case (sel) 0: mux_6744 = 1'h0; 1: mux_6744 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6745;
  wire [0:0] v_6746;
  wire [0:0] v_6747;
  wire [0:0] v_6748;
  wire [0:0] v_6749;
  function [0:0] mux_6749(input [0:0] sel);
    case (sel) 0: mux_6749 = 1'h0; 1: mux_6749 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6750;
  wire [0:0] vin0_consume_en_6751;
  wire [0:0] vout_canPeek_6751;
  wire [7:0] vout_peek_6751;
  wire [0:0] v_6752;
  wire [0:0] v_6753;
  function [0:0] mux_6753(input [0:0] sel);
    case (sel) 0: mux_6753 = 1'h0; 1: mux_6753 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6754;
  function [0:0] mux_6754(input [0:0] sel);
    case (sel) 0: mux_6754 = 1'h0; 1: mux_6754 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6755;
  wire [0:0] v_6756;
  wire [0:0] v_6757;
  wire [0:0] v_6758;
  wire [0:0] v_6759;
  wire [0:0] v_6760;
  wire [0:0] v_6761;
  function [0:0] mux_6761(input [0:0] sel);
    case (sel) 0: mux_6761 = 1'h0; 1: mux_6761 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6762;
  wire [0:0] v_6763;
  wire [0:0] v_6764;
  wire [0:0] v_6765;
  wire [0:0] v_6766;
  function [0:0] mux_6766(input [0:0] sel);
    case (sel) 0: mux_6766 = 1'h0; 1: mux_6766 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6767;
  wire [0:0] v_6768;
  wire [0:0] v_6769;
  wire [0:0] v_6770;
  function [0:0] mux_6770(input [0:0] sel);
    case (sel) 0: mux_6770 = 1'h0; 1: mux_6770 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6771;
  function [0:0] mux_6771(input [0:0] sel);
    case (sel) 0: mux_6771 = 1'h0; 1: mux_6771 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6772 = 1'h0;
  wire [0:0] v_6773;
  wire [0:0] v_6774;
  wire [0:0] act_6775;
  wire [0:0] v_6776;
  wire [0:0] v_6777;
  wire [0:0] v_6778;
  wire [0:0] vin0_consume_en_6779;
  wire [0:0] vout_canPeek_6779;
  wire [7:0] vout_peek_6779;
  wire [0:0] v_6780;
  wire [0:0] v_6781;
  function [0:0] mux_6781(input [0:0] sel);
    case (sel) 0: mux_6781 = 1'h0; 1: mux_6781 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6782;
  wire [0:0] v_6783;
  wire [0:0] v_6784;
  wire [0:0] v_6785;
  wire [0:0] v_6786;
  function [0:0] mux_6786(input [0:0] sel);
    case (sel) 0: mux_6786 = 1'h0; 1: mux_6786 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6787;
  wire [0:0] vin0_consume_en_6788;
  wire [0:0] vout_canPeek_6788;
  wire [7:0] vout_peek_6788;
  wire [0:0] v_6789;
  wire [0:0] v_6790;
  function [0:0] mux_6790(input [0:0] sel);
    case (sel) 0: mux_6790 = 1'h0; 1: mux_6790 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6791;
  function [0:0] mux_6791(input [0:0] sel);
    case (sel) 0: mux_6791 = 1'h0; 1: mux_6791 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6792;
  wire [0:0] v_6793;
  wire [0:0] v_6794;
  wire [0:0] v_6795;
  wire [0:0] v_6796;
  wire [0:0] v_6797;
  wire [0:0] v_6798;
  function [0:0] mux_6798(input [0:0] sel);
    case (sel) 0: mux_6798 = 1'h0; 1: mux_6798 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6799;
  function [0:0] mux_6799(input [0:0] sel);
    case (sel) 0: mux_6799 = 1'h0; 1: mux_6799 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6800;
  wire [0:0] v_6801;
  wire [0:0] v_6802;
  wire [0:0] v_6803;
  function [0:0] mux_6803(input [0:0] sel);
    case (sel) 0: mux_6803 = 1'h0; 1: mux_6803 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6804;
  function [0:0] mux_6804(input [0:0] sel);
    case (sel) 0: mux_6804 = 1'h0; 1: mux_6804 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6805;
  wire [0:0] v_6806;
  wire [0:0] v_6807;
  wire [0:0] v_6808;
  wire [0:0] v_6809;
  wire [0:0] v_6810;
  function [0:0] mux_6810(input [0:0] sel);
    case (sel) 0: mux_6810 = 1'h0; 1: mux_6810 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6811;
  function [0:0] mux_6811(input [0:0] sel);
    case (sel) 0: mux_6811 = 1'h0; 1: mux_6811 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6812;
  wire [0:0] v_6813;
  wire [0:0] v_6814;
  wire [0:0] v_6815;
  function [0:0] mux_6815(input [0:0] sel);
    case (sel) 0: mux_6815 = 1'h0; 1: mux_6815 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6816;
  function [0:0] mux_6816(input [0:0] sel);
    case (sel) 0: mux_6816 = 1'h0; 1: mux_6816 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6817;
  wire [0:0] v_6818;
  wire [0:0] v_6819;
  wire [0:0] v_6820;
  wire [0:0] v_6821;
  wire [0:0] v_6822;
  function [0:0] mux_6822(input [0:0] sel);
    case (sel) 0: mux_6822 = 1'h0; 1: mux_6822 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6823;
  wire [0:0] v_6824;
  wire [0:0] v_6825;
  wire [0:0] v_6826;
  wire [0:0] v_6827;
  function [0:0] mux_6827(input [0:0] sel);
    case (sel) 0: mux_6827 = 1'h0; 1: mux_6827 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6828;
  wire [0:0] v_6829;
  wire [0:0] v_6830;
  wire [0:0] v_6831;
  function [0:0] mux_6831(input [0:0] sel);
    case (sel) 0: mux_6831 = 1'h0; 1: mux_6831 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6832;
  function [0:0] mux_6832(input [0:0] sel);
    case (sel) 0: mux_6832 = 1'h0; 1: mux_6832 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6833 = 1'h0;
  wire [0:0] v_6834;
  wire [0:0] v_6835;
  wire [0:0] act_6836;
  wire [0:0] v_6837;
  wire [0:0] v_6838;
  wire [0:0] v_6839;
  reg [0:0] v_6840 = 1'h0;
  wire [0:0] v_6841;
  wire [0:0] v_6842;
  wire [0:0] act_6843;
  wire [0:0] v_6844;
  wire [0:0] v_6845;
  wire [0:0] v_6846;
  reg [0:0] v_6847 = 1'h0;
  wire [0:0] v_6848;
  wire [0:0] v_6849;
  wire [0:0] act_6850;
  wire [0:0] v_6851;
  wire [0:0] v_6852;
  wire [0:0] v_6853;
  wire [0:0] vin0_consume_en_6854;
  wire [0:0] vout_canPeek_6854;
  wire [7:0] vout_peek_6854;
  wire [0:0] v_6855;
  wire [0:0] v_6856;
  function [0:0] mux_6856(input [0:0] sel);
    case (sel) 0: mux_6856 = 1'h0; 1: mux_6856 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6857;
  wire [0:0] v_6858;
  wire [0:0] v_6859;
  wire [0:0] v_6860;
  wire [0:0] v_6861;
  function [0:0] mux_6861(input [0:0] sel);
    case (sel) 0: mux_6861 = 1'h0; 1: mux_6861 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6862;
  wire [0:0] vin0_consume_en_6863;
  wire [0:0] vout_canPeek_6863;
  wire [7:0] vout_peek_6863;
  wire [0:0] v_6864;
  wire [0:0] v_6865;
  function [0:0] mux_6865(input [0:0] sel);
    case (sel) 0: mux_6865 = 1'h0; 1: mux_6865 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6866;
  function [0:0] mux_6866(input [0:0] sel);
    case (sel) 0: mux_6866 = 1'h0; 1: mux_6866 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6867;
  wire [0:0] v_6868;
  wire [0:0] v_6869;
  wire [0:0] v_6870;
  wire [0:0] v_6871;
  wire [0:0] v_6872;
  wire [0:0] v_6873;
  function [0:0] mux_6873(input [0:0] sel);
    case (sel) 0: mux_6873 = 1'h0; 1: mux_6873 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6874;
  wire [0:0] v_6875;
  wire [0:0] v_6876;
  wire [0:0] v_6877;
  wire [0:0] v_6878;
  function [0:0] mux_6878(input [0:0] sel);
    case (sel) 0: mux_6878 = 1'h0; 1: mux_6878 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6879;
  wire [0:0] v_6880;
  wire [0:0] v_6881;
  wire [0:0] v_6882;
  function [0:0] mux_6882(input [0:0] sel);
    case (sel) 0: mux_6882 = 1'h0; 1: mux_6882 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6883;
  function [0:0] mux_6883(input [0:0] sel);
    case (sel) 0: mux_6883 = 1'h0; 1: mux_6883 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6884 = 1'h0;
  wire [0:0] v_6885;
  wire [0:0] v_6886;
  wire [0:0] act_6887;
  wire [0:0] v_6888;
  wire [0:0] v_6889;
  wire [0:0] v_6890;
  wire [0:0] vin0_consume_en_6891;
  wire [0:0] vout_canPeek_6891;
  wire [7:0] vout_peek_6891;
  wire [0:0] v_6892;
  wire [0:0] v_6893;
  function [0:0] mux_6893(input [0:0] sel);
    case (sel) 0: mux_6893 = 1'h0; 1: mux_6893 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6894;
  wire [0:0] v_6895;
  wire [0:0] v_6896;
  wire [0:0] v_6897;
  wire [0:0] v_6898;
  function [0:0] mux_6898(input [0:0] sel);
    case (sel) 0: mux_6898 = 1'h0; 1: mux_6898 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6899;
  wire [0:0] vin0_consume_en_6900;
  wire [0:0] vout_canPeek_6900;
  wire [7:0] vout_peek_6900;
  wire [0:0] v_6901;
  wire [0:0] v_6902;
  function [0:0] mux_6902(input [0:0] sel);
    case (sel) 0: mux_6902 = 1'h0; 1: mux_6902 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6903;
  function [0:0] mux_6903(input [0:0] sel);
    case (sel) 0: mux_6903 = 1'h0; 1: mux_6903 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6904;
  wire [0:0] v_6905;
  wire [0:0] v_6906;
  wire [0:0] v_6907;
  wire [0:0] v_6908;
  wire [0:0] v_6909;
  wire [0:0] v_6910;
  function [0:0] mux_6910(input [0:0] sel);
    case (sel) 0: mux_6910 = 1'h0; 1: mux_6910 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6911;
  function [0:0] mux_6911(input [0:0] sel);
    case (sel) 0: mux_6911 = 1'h0; 1: mux_6911 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6912;
  wire [0:0] v_6913;
  wire [0:0] v_6914;
  wire [0:0] v_6915;
  function [0:0] mux_6915(input [0:0] sel);
    case (sel) 0: mux_6915 = 1'h0; 1: mux_6915 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6916;
  function [0:0] mux_6916(input [0:0] sel);
    case (sel) 0: mux_6916 = 1'h0; 1: mux_6916 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6917;
  wire [0:0] v_6918;
  wire [0:0] v_6919;
  wire [0:0] v_6920;
  wire [0:0] v_6921;
  wire [0:0] v_6922;
  function [0:0] mux_6922(input [0:0] sel);
    case (sel) 0: mux_6922 = 1'h0; 1: mux_6922 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6923;
  wire [0:0] v_6924;
  wire [0:0] v_6925;
  wire [0:0] v_6926;
  wire [0:0] v_6927;
  function [0:0] mux_6927(input [0:0] sel);
    case (sel) 0: mux_6927 = 1'h0; 1: mux_6927 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6928;
  wire [0:0] v_6929;
  wire [0:0] v_6930;
  wire [0:0] v_6931;
  function [0:0] mux_6931(input [0:0] sel);
    case (sel) 0: mux_6931 = 1'h0; 1: mux_6931 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6932;
  function [0:0] mux_6932(input [0:0] sel);
    case (sel) 0: mux_6932 = 1'h0; 1: mux_6932 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6933 = 1'h0;
  wire [0:0] v_6934;
  wire [0:0] v_6935;
  wire [0:0] act_6936;
  wire [0:0] v_6937;
  wire [0:0] v_6938;
  wire [0:0] v_6939;
  reg [0:0] v_6940 = 1'h0;
  wire [0:0] v_6941;
  wire [0:0] v_6942;
  wire [0:0] act_6943;
  wire [0:0] v_6944;
  wire [0:0] v_6945;
  wire [0:0] v_6946;
  wire [0:0] vin0_consume_en_6947;
  wire [0:0] vout_canPeek_6947;
  wire [7:0] vout_peek_6947;
  wire [0:0] v_6948;
  wire [0:0] v_6949;
  function [0:0] mux_6949(input [0:0] sel);
    case (sel) 0: mux_6949 = 1'h0; 1: mux_6949 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6950;
  wire [0:0] v_6951;
  wire [0:0] v_6952;
  wire [0:0] v_6953;
  wire [0:0] v_6954;
  function [0:0] mux_6954(input [0:0] sel);
    case (sel) 0: mux_6954 = 1'h0; 1: mux_6954 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6955;
  wire [0:0] vin0_consume_en_6956;
  wire [0:0] vout_canPeek_6956;
  wire [7:0] vout_peek_6956;
  wire [0:0] v_6957;
  wire [0:0] v_6958;
  function [0:0] mux_6958(input [0:0] sel);
    case (sel) 0: mux_6958 = 1'h0; 1: mux_6958 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6959;
  function [0:0] mux_6959(input [0:0] sel);
    case (sel) 0: mux_6959 = 1'h0; 1: mux_6959 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6960;
  wire [0:0] v_6961;
  wire [0:0] v_6962;
  wire [0:0] v_6963;
  wire [0:0] v_6964;
  wire [0:0] v_6965;
  wire [0:0] v_6966;
  function [0:0] mux_6966(input [0:0] sel);
    case (sel) 0: mux_6966 = 1'h0; 1: mux_6966 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6967;
  wire [0:0] v_6968;
  wire [0:0] v_6969;
  wire [0:0] v_6970;
  wire [0:0] v_6971;
  function [0:0] mux_6971(input [0:0] sel);
    case (sel) 0: mux_6971 = 1'h0; 1: mux_6971 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6972;
  wire [0:0] v_6973;
  wire [0:0] v_6974;
  wire [0:0] v_6975;
  function [0:0] mux_6975(input [0:0] sel);
    case (sel) 0: mux_6975 = 1'h0; 1: mux_6975 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6976;
  function [0:0] mux_6976(input [0:0] sel);
    case (sel) 0: mux_6976 = 1'h0; 1: mux_6976 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6977 = 1'h0;
  wire [0:0] v_6978;
  wire [0:0] v_6979;
  wire [0:0] act_6980;
  wire [0:0] v_6981;
  wire [0:0] v_6982;
  wire [0:0] v_6983;
  wire [0:0] vin0_consume_en_6984;
  wire [0:0] vout_canPeek_6984;
  wire [7:0] vout_peek_6984;
  wire [0:0] v_6985;
  wire [0:0] v_6986;
  function [0:0] mux_6986(input [0:0] sel);
    case (sel) 0: mux_6986 = 1'h0; 1: mux_6986 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6987;
  wire [0:0] v_6988;
  wire [0:0] v_6989;
  wire [0:0] v_6990;
  wire [0:0] v_6991;
  function [0:0] mux_6991(input [0:0] sel);
    case (sel) 0: mux_6991 = 1'h0; 1: mux_6991 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6992;
  wire [0:0] vin0_consume_en_6993;
  wire [0:0] vout_canPeek_6993;
  wire [7:0] vout_peek_6993;
  wire [0:0] v_6994;
  wire [0:0] v_6995;
  function [0:0] mux_6995(input [0:0] sel);
    case (sel) 0: mux_6995 = 1'h0; 1: mux_6995 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6996;
  function [0:0] mux_6996(input [0:0] sel);
    case (sel) 0: mux_6996 = 1'h0; 1: mux_6996 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6997;
  wire [0:0] v_6998;
  wire [0:0] v_6999;
  wire [0:0] v_7000;
  wire [0:0] v_7001;
  wire [0:0] v_7002;
  wire [0:0] v_7003;
  function [0:0] mux_7003(input [0:0] sel);
    case (sel) 0: mux_7003 = 1'h0; 1: mux_7003 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7004;
  function [0:0] mux_7004(input [0:0] sel);
    case (sel) 0: mux_7004 = 1'h0; 1: mux_7004 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7005;
  wire [0:0] v_7006;
  wire [0:0] v_7007;
  wire [0:0] v_7008;
  function [0:0] mux_7008(input [0:0] sel);
    case (sel) 0: mux_7008 = 1'h0; 1: mux_7008 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7009;
  function [0:0] mux_7009(input [0:0] sel);
    case (sel) 0: mux_7009 = 1'h0; 1: mux_7009 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7010;
  wire [0:0] v_7011;
  wire [0:0] v_7012;
  wire [0:0] v_7013;
  wire [0:0] v_7014;
  wire [0:0] v_7015;
  function [0:0] mux_7015(input [0:0] sel);
    case (sel) 0: mux_7015 = 1'h0; 1: mux_7015 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7016;
  function [0:0] mux_7016(input [0:0] sel);
    case (sel) 0: mux_7016 = 1'h0; 1: mux_7016 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7017;
  wire [0:0] v_7018;
  wire [0:0] v_7019;
  wire [0:0] v_7020;
  function [0:0] mux_7020(input [0:0] sel);
    case (sel) 0: mux_7020 = 1'h0; 1: mux_7020 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7021;
  function [0:0] mux_7021(input [0:0] sel);
    case (sel) 0: mux_7021 = 1'h0; 1: mux_7021 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7022;
  wire [0:0] v_7023;
  wire [0:0] v_7024;
  wire [0:0] v_7025;
  wire [0:0] v_7026;
  wire [0:0] v_7027;
  function [0:0] mux_7027(input [0:0] sel);
    case (sel) 0: mux_7027 = 1'h0; 1: mux_7027 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7028;
  function [0:0] mux_7028(input [0:0] sel);
    case (sel) 0: mux_7028 = 1'h0; 1: mux_7028 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7029;
  wire [0:0] v_7030;
  wire [0:0] v_7031;
  wire [0:0] v_7032;
  function [0:0] mux_7032(input [0:0] sel);
    case (sel) 0: mux_7032 = 1'h0; 1: mux_7032 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7033;
  function [0:0] mux_7033(input [0:0] sel);
    case (sel) 0: mux_7033 = 1'h0; 1: mux_7033 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7034;
  wire [0:0] v_7035;
  wire [0:0] v_7036;
  wire [0:0] v_7037;
  wire [0:0] v_7038;
  wire [0:0] v_7039;
  function [0:0] mux_7039(input [0:0] sel);
    case (sel) 0: mux_7039 = 1'h0; 1: mux_7039 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7040;
  function [0:0] mux_7040(input [0:0] sel);
    case (sel) 0: mux_7040 = 1'h0; 1: mux_7040 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7041;
  wire [0:0] v_7042;
  wire [0:0] v_7043;
  wire [0:0] v_7044;
  function [0:0] mux_7044(input [0:0] sel);
    case (sel) 0: mux_7044 = 1'h0; 1: mux_7044 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7045;
  function [0:0] mux_7045(input [0:0] sel);
    case (sel) 0: mux_7045 = 1'h0; 1: mux_7045 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7046;
  wire [0:0] v_7047;
  wire [0:0] v_7048;
  wire [0:0] v_7049;
  wire [0:0] v_7050;
  wire [0:0] v_7051;
  function [0:0] mux_7051(input [0:0] sel);
    case (sel) 0: mux_7051 = 1'h0; 1: mux_7051 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7052;
  wire [0:0] v_7053;
  wire [0:0] v_7054;
  wire [0:0] v_7055;
  wire [0:0] v_7056;
  function [0:0] mux_7056(input [0:0] sel);
    case (sel) 0: mux_7056 = 1'h0; 1: mux_7056 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7057;
  wire [0:0] v_7058;
  wire [0:0] v_7059;
  wire [0:0] v_7060;
  function [0:0] mux_7060(input [0:0] sel);
    case (sel) 0: mux_7060 = 1'h0; 1: mux_7060 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7061;
  function [0:0] mux_7061(input [0:0] sel);
    case (sel) 0: mux_7061 = 1'h0; 1: mux_7061 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7062 = 1'h0;
  wire [0:0] v_7063;
  wire [0:0] v_7064;
  wire [0:0] act_7065;
  wire [0:0] v_7066;
  wire [0:0] v_7067;
  wire [0:0] v_7068;
  reg [0:0] v_7069 = 1'h0;
  wire [0:0] v_7070;
  wire [0:0] v_7071;
  wire [0:0] act_7072;
  wire [0:0] v_7073;
  wire [0:0] v_7074;
  wire [0:0] v_7075;
  reg [0:0] v_7076 = 1'h0;
  wire [0:0] v_7077;
  wire [0:0] v_7078;
  wire [0:0] act_7079;
  wire [0:0] v_7080;
  wire [0:0] v_7081;
  wire [0:0] v_7082;
  reg [0:0] v_7083 = 1'h0;
  wire [0:0] v_7084;
  wire [0:0] v_7085;
  wire [0:0] act_7086;
  wire [0:0] v_7087;
  wire [0:0] v_7088;
  wire [0:0] v_7089;
  reg [0:0] v_7090 = 1'h0;
  wire [0:0] v_7091;
  wire [0:0] v_7092;
  wire [0:0] act_7093;
  wire [0:0] v_7094;
  wire [0:0] v_7095;
  wire [0:0] v_7096;
  wire [0:0] vin0_consume_en_7097;
  wire [0:0] vout_canPeek_7097;
  wire [7:0] vout_peek_7097;
  wire [0:0] v_7098;
  wire [0:0] v_7099;
  function [0:0] mux_7099(input [0:0] sel);
    case (sel) 0: mux_7099 = 1'h0; 1: mux_7099 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7100;
  wire [0:0] v_7101;
  wire [0:0] v_7102;
  wire [0:0] v_7103;
  wire [0:0] v_7104;
  function [0:0] mux_7104(input [0:0] sel);
    case (sel) 0: mux_7104 = 1'h0; 1: mux_7104 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7105;
  wire [0:0] vin0_consume_en_7106;
  wire [0:0] vout_canPeek_7106;
  wire [7:0] vout_peek_7106;
  wire [0:0] v_7107;
  wire [0:0] v_7108;
  function [0:0] mux_7108(input [0:0] sel);
    case (sel) 0: mux_7108 = 1'h0; 1: mux_7108 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7109;
  function [0:0] mux_7109(input [0:0] sel);
    case (sel) 0: mux_7109 = 1'h0; 1: mux_7109 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7110;
  wire [0:0] v_7111;
  wire [0:0] v_7112;
  wire [0:0] v_7113;
  wire [0:0] v_7114;
  wire [0:0] v_7115;
  wire [0:0] v_7116;
  function [0:0] mux_7116(input [0:0] sel);
    case (sel) 0: mux_7116 = 1'h0; 1: mux_7116 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7117;
  wire [0:0] v_7118;
  wire [0:0] v_7119;
  wire [0:0] v_7120;
  wire [0:0] v_7121;
  function [0:0] mux_7121(input [0:0] sel);
    case (sel) 0: mux_7121 = 1'h0; 1: mux_7121 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7122;
  wire [0:0] v_7123;
  wire [0:0] v_7124;
  wire [0:0] v_7125;
  function [0:0] mux_7125(input [0:0] sel);
    case (sel) 0: mux_7125 = 1'h0; 1: mux_7125 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7126;
  function [0:0] mux_7126(input [0:0] sel);
    case (sel) 0: mux_7126 = 1'h0; 1: mux_7126 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7127 = 1'h0;
  wire [0:0] v_7128;
  wire [0:0] v_7129;
  wire [0:0] act_7130;
  wire [0:0] v_7131;
  wire [0:0] v_7132;
  wire [0:0] v_7133;
  wire [0:0] vin0_consume_en_7134;
  wire [0:0] vout_canPeek_7134;
  wire [7:0] vout_peek_7134;
  wire [0:0] v_7135;
  wire [0:0] v_7136;
  function [0:0] mux_7136(input [0:0] sel);
    case (sel) 0: mux_7136 = 1'h0; 1: mux_7136 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7137;
  wire [0:0] v_7138;
  wire [0:0] v_7139;
  wire [0:0] v_7140;
  wire [0:0] v_7141;
  function [0:0] mux_7141(input [0:0] sel);
    case (sel) 0: mux_7141 = 1'h0; 1: mux_7141 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7142;
  wire [0:0] vin0_consume_en_7143;
  wire [0:0] vout_canPeek_7143;
  wire [7:0] vout_peek_7143;
  wire [0:0] v_7144;
  wire [0:0] v_7145;
  function [0:0] mux_7145(input [0:0] sel);
    case (sel) 0: mux_7145 = 1'h0; 1: mux_7145 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7146;
  function [0:0] mux_7146(input [0:0] sel);
    case (sel) 0: mux_7146 = 1'h0; 1: mux_7146 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7147;
  wire [0:0] v_7148;
  wire [0:0] v_7149;
  wire [0:0] v_7150;
  wire [0:0] v_7151;
  wire [0:0] v_7152;
  wire [0:0] v_7153;
  function [0:0] mux_7153(input [0:0] sel);
    case (sel) 0: mux_7153 = 1'h0; 1: mux_7153 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7154;
  function [0:0] mux_7154(input [0:0] sel);
    case (sel) 0: mux_7154 = 1'h0; 1: mux_7154 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7155;
  wire [0:0] v_7156;
  wire [0:0] v_7157;
  wire [0:0] v_7158;
  function [0:0] mux_7158(input [0:0] sel);
    case (sel) 0: mux_7158 = 1'h0; 1: mux_7158 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7159;
  function [0:0] mux_7159(input [0:0] sel);
    case (sel) 0: mux_7159 = 1'h0; 1: mux_7159 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7160;
  wire [0:0] v_7161;
  wire [0:0] v_7162;
  wire [0:0] v_7163;
  wire [0:0] v_7164;
  wire [0:0] v_7165;
  function [0:0] mux_7165(input [0:0] sel);
    case (sel) 0: mux_7165 = 1'h0; 1: mux_7165 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7166;
  wire [0:0] v_7167;
  wire [0:0] v_7168;
  wire [0:0] v_7169;
  wire [0:0] v_7170;
  function [0:0] mux_7170(input [0:0] sel);
    case (sel) 0: mux_7170 = 1'h0; 1: mux_7170 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7171;
  wire [0:0] v_7172;
  wire [0:0] v_7173;
  wire [0:0] v_7174;
  function [0:0] mux_7174(input [0:0] sel);
    case (sel) 0: mux_7174 = 1'h0; 1: mux_7174 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7175;
  function [0:0] mux_7175(input [0:0] sel);
    case (sel) 0: mux_7175 = 1'h0; 1: mux_7175 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7176 = 1'h0;
  wire [0:0] v_7177;
  wire [0:0] v_7178;
  wire [0:0] act_7179;
  wire [0:0] v_7180;
  wire [0:0] v_7181;
  wire [0:0] v_7182;
  reg [0:0] v_7183 = 1'h0;
  wire [0:0] v_7184;
  wire [0:0] v_7185;
  wire [0:0] act_7186;
  wire [0:0] v_7187;
  wire [0:0] v_7188;
  wire [0:0] v_7189;
  wire [0:0] vin0_consume_en_7190;
  wire [0:0] vout_canPeek_7190;
  wire [7:0] vout_peek_7190;
  wire [0:0] v_7191;
  wire [0:0] v_7192;
  function [0:0] mux_7192(input [0:0] sel);
    case (sel) 0: mux_7192 = 1'h0; 1: mux_7192 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7193;
  wire [0:0] v_7194;
  wire [0:0] v_7195;
  wire [0:0] v_7196;
  wire [0:0] v_7197;
  function [0:0] mux_7197(input [0:0] sel);
    case (sel) 0: mux_7197 = 1'h0; 1: mux_7197 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7198;
  wire [0:0] vin0_consume_en_7199;
  wire [0:0] vout_canPeek_7199;
  wire [7:0] vout_peek_7199;
  wire [0:0] v_7200;
  wire [0:0] v_7201;
  function [0:0] mux_7201(input [0:0] sel);
    case (sel) 0: mux_7201 = 1'h0; 1: mux_7201 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7202;
  function [0:0] mux_7202(input [0:0] sel);
    case (sel) 0: mux_7202 = 1'h0; 1: mux_7202 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7203;
  wire [0:0] v_7204;
  wire [0:0] v_7205;
  wire [0:0] v_7206;
  wire [0:0] v_7207;
  wire [0:0] v_7208;
  wire [0:0] v_7209;
  function [0:0] mux_7209(input [0:0] sel);
    case (sel) 0: mux_7209 = 1'h0; 1: mux_7209 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7210;
  wire [0:0] v_7211;
  wire [0:0] v_7212;
  wire [0:0] v_7213;
  wire [0:0] v_7214;
  function [0:0] mux_7214(input [0:0] sel);
    case (sel) 0: mux_7214 = 1'h0; 1: mux_7214 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7215;
  wire [0:0] v_7216;
  wire [0:0] v_7217;
  wire [0:0] v_7218;
  function [0:0] mux_7218(input [0:0] sel);
    case (sel) 0: mux_7218 = 1'h0; 1: mux_7218 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7219;
  function [0:0] mux_7219(input [0:0] sel);
    case (sel) 0: mux_7219 = 1'h0; 1: mux_7219 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7220 = 1'h0;
  wire [0:0] v_7221;
  wire [0:0] v_7222;
  wire [0:0] act_7223;
  wire [0:0] v_7224;
  wire [0:0] v_7225;
  wire [0:0] v_7226;
  wire [0:0] vin0_consume_en_7227;
  wire [0:0] vout_canPeek_7227;
  wire [7:0] vout_peek_7227;
  wire [0:0] v_7228;
  wire [0:0] v_7229;
  function [0:0] mux_7229(input [0:0] sel);
    case (sel) 0: mux_7229 = 1'h0; 1: mux_7229 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7230;
  wire [0:0] v_7231;
  wire [0:0] v_7232;
  wire [0:0] v_7233;
  wire [0:0] v_7234;
  function [0:0] mux_7234(input [0:0] sel);
    case (sel) 0: mux_7234 = 1'h0; 1: mux_7234 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7235;
  wire [0:0] vin0_consume_en_7236;
  wire [0:0] vout_canPeek_7236;
  wire [7:0] vout_peek_7236;
  wire [0:0] v_7237;
  wire [0:0] v_7238;
  function [0:0] mux_7238(input [0:0] sel);
    case (sel) 0: mux_7238 = 1'h0; 1: mux_7238 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7239;
  function [0:0] mux_7239(input [0:0] sel);
    case (sel) 0: mux_7239 = 1'h0; 1: mux_7239 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7240;
  wire [0:0] v_7241;
  wire [0:0] v_7242;
  wire [0:0] v_7243;
  wire [0:0] v_7244;
  wire [0:0] v_7245;
  wire [0:0] v_7246;
  function [0:0] mux_7246(input [0:0] sel);
    case (sel) 0: mux_7246 = 1'h0; 1: mux_7246 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7247;
  function [0:0] mux_7247(input [0:0] sel);
    case (sel) 0: mux_7247 = 1'h0; 1: mux_7247 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7248;
  wire [0:0] v_7249;
  wire [0:0] v_7250;
  wire [0:0] v_7251;
  function [0:0] mux_7251(input [0:0] sel);
    case (sel) 0: mux_7251 = 1'h0; 1: mux_7251 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7252;
  function [0:0] mux_7252(input [0:0] sel);
    case (sel) 0: mux_7252 = 1'h0; 1: mux_7252 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7253;
  wire [0:0] v_7254;
  wire [0:0] v_7255;
  wire [0:0] v_7256;
  wire [0:0] v_7257;
  wire [0:0] v_7258;
  function [0:0] mux_7258(input [0:0] sel);
    case (sel) 0: mux_7258 = 1'h0; 1: mux_7258 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7259;
  function [0:0] mux_7259(input [0:0] sel);
    case (sel) 0: mux_7259 = 1'h0; 1: mux_7259 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7260;
  wire [0:0] v_7261;
  wire [0:0] v_7262;
  wire [0:0] v_7263;
  function [0:0] mux_7263(input [0:0] sel);
    case (sel) 0: mux_7263 = 1'h0; 1: mux_7263 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7264;
  function [0:0] mux_7264(input [0:0] sel);
    case (sel) 0: mux_7264 = 1'h0; 1: mux_7264 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7265;
  wire [0:0] v_7266;
  wire [0:0] v_7267;
  wire [0:0] v_7268;
  wire [0:0] v_7269;
  wire [0:0] v_7270;
  function [0:0] mux_7270(input [0:0] sel);
    case (sel) 0: mux_7270 = 1'h0; 1: mux_7270 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7271;
  wire [0:0] v_7272;
  wire [0:0] v_7273;
  wire [0:0] v_7274;
  wire [0:0] v_7275;
  function [0:0] mux_7275(input [0:0] sel);
    case (sel) 0: mux_7275 = 1'h0; 1: mux_7275 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7276;
  wire [0:0] v_7277;
  wire [0:0] v_7278;
  wire [0:0] v_7279;
  function [0:0] mux_7279(input [0:0] sel);
    case (sel) 0: mux_7279 = 1'h0; 1: mux_7279 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7280;
  function [0:0] mux_7280(input [0:0] sel);
    case (sel) 0: mux_7280 = 1'h0; 1: mux_7280 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7281 = 1'h0;
  wire [0:0] v_7282;
  wire [0:0] v_7283;
  wire [0:0] act_7284;
  wire [0:0] v_7285;
  wire [0:0] v_7286;
  wire [0:0] v_7287;
  reg [0:0] v_7288 = 1'h0;
  wire [0:0] v_7289;
  wire [0:0] v_7290;
  wire [0:0] act_7291;
  wire [0:0] v_7292;
  wire [0:0] v_7293;
  wire [0:0] v_7294;
  reg [0:0] v_7295 = 1'h0;
  wire [0:0] v_7296;
  wire [0:0] v_7297;
  wire [0:0] act_7298;
  wire [0:0] v_7299;
  wire [0:0] v_7300;
  wire [0:0] v_7301;
  wire [0:0] vin0_consume_en_7302;
  wire [0:0] vout_canPeek_7302;
  wire [7:0] vout_peek_7302;
  wire [0:0] v_7303;
  wire [0:0] v_7304;
  function [0:0] mux_7304(input [0:0] sel);
    case (sel) 0: mux_7304 = 1'h0; 1: mux_7304 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7305;
  wire [0:0] v_7306;
  wire [0:0] v_7307;
  wire [0:0] v_7308;
  wire [0:0] v_7309;
  function [0:0] mux_7309(input [0:0] sel);
    case (sel) 0: mux_7309 = 1'h0; 1: mux_7309 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7310;
  wire [0:0] vin0_consume_en_7311;
  wire [0:0] vout_canPeek_7311;
  wire [7:0] vout_peek_7311;
  wire [0:0] v_7312;
  wire [0:0] v_7313;
  function [0:0] mux_7313(input [0:0] sel);
    case (sel) 0: mux_7313 = 1'h0; 1: mux_7313 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7314;
  function [0:0] mux_7314(input [0:0] sel);
    case (sel) 0: mux_7314 = 1'h0; 1: mux_7314 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7315;
  wire [0:0] v_7316;
  wire [0:0] v_7317;
  wire [0:0] v_7318;
  wire [0:0] v_7319;
  wire [0:0] v_7320;
  wire [0:0] v_7321;
  function [0:0] mux_7321(input [0:0] sel);
    case (sel) 0: mux_7321 = 1'h0; 1: mux_7321 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7322;
  wire [0:0] v_7323;
  wire [0:0] v_7324;
  wire [0:0] v_7325;
  wire [0:0] v_7326;
  function [0:0] mux_7326(input [0:0] sel);
    case (sel) 0: mux_7326 = 1'h0; 1: mux_7326 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7327;
  wire [0:0] v_7328;
  wire [0:0] v_7329;
  wire [0:0] v_7330;
  function [0:0] mux_7330(input [0:0] sel);
    case (sel) 0: mux_7330 = 1'h0; 1: mux_7330 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7331;
  function [0:0] mux_7331(input [0:0] sel);
    case (sel) 0: mux_7331 = 1'h0; 1: mux_7331 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7332 = 1'h0;
  wire [0:0] v_7333;
  wire [0:0] v_7334;
  wire [0:0] act_7335;
  wire [0:0] v_7336;
  wire [0:0] v_7337;
  wire [0:0] v_7338;
  wire [0:0] vin0_consume_en_7339;
  wire [0:0] vout_canPeek_7339;
  wire [7:0] vout_peek_7339;
  wire [0:0] v_7340;
  wire [0:0] v_7341;
  function [0:0] mux_7341(input [0:0] sel);
    case (sel) 0: mux_7341 = 1'h0; 1: mux_7341 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7342;
  wire [0:0] v_7343;
  wire [0:0] v_7344;
  wire [0:0] v_7345;
  wire [0:0] v_7346;
  function [0:0] mux_7346(input [0:0] sel);
    case (sel) 0: mux_7346 = 1'h0; 1: mux_7346 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7347;
  wire [0:0] vin0_consume_en_7348;
  wire [0:0] vout_canPeek_7348;
  wire [7:0] vout_peek_7348;
  wire [0:0] v_7349;
  wire [0:0] v_7350;
  function [0:0] mux_7350(input [0:0] sel);
    case (sel) 0: mux_7350 = 1'h0; 1: mux_7350 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7351;
  function [0:0] mux_7351(input [0:0] sel);
    case (sel) 0: mux_7351 = 1'h0; 1: mux_7351 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7352;
  wire [0:0] v_7353;
  wire [0:0] v_7354;
  wire [0:0] v_7355;
  wire [0:0] v_7356;
  wire [0:0] v_7357;
  wire [0:0] v_7358;
  function [0:0] mux_7358(input [0:0] sel);
    case (sel) 0: mux_7358 = 1'h0; 1: mux_7358 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7359;
  function [0:0] mux_7359(input [0:0] sel);
    case (sel) 0: mux_7359 = 1'h0; 1: mux_7359 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7360;
  wire [0:0] v_7361;
  wire [0:0] v_7362;
  wire [0:0] v_7363;
  function [0:0] mux_7363(input [0:0] sel);
    case (sel) 0: mux_7363 = 1'h0; 1: mux_7363 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7364;
  function [0:0] mux_7364(input [0:0] sel);
    case (sel) 0: mux_7364 = 1'h0; 1: mux_7364 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7365;
  wire [0:0] v_7366;
  wire [0:0] v_7367;
  wire [0:0] v_7368;
  wire [0:0] v_7369;
  wire [0:0] v_7370;
  function [0:0] mux_7370(input [0:0] sel);
    case (sel) 0: mux_7370 = 1'h0; 1: mux_7370 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7371;
  wire [0:0] v_7372;
  wire [0:0] v_7373;
  wire [0:0] v_7374;
  wire [0:0] v_7375;
  function [0:0] mux_7375(input [0:0] sel);
    case (sel) 0: mux_7375 = 1'h0; 1: mux_7375 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7376;
  wire [0:0] v_7377;
  wire [0:0] v_7378;
  wire [0:0] v_7379;
  function [0:0] mux_7379(input [0:0] sel);
    case (sel) 0: mux_7379 = 1'h0; 1: mux_7379 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7380;
  function [0:0] mux_7380(input [0:0] sel);
    case (sel) 0: mux_7380 = 1'h0; 1: mux_7380 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7381 = 1'h0;
  wire [0:0] v_7382;
  wire [0:0] v_7383;
  wire [0:0] act_7384;
  wire [0:0] v_7385;
  wire [0:0] v_7386;
  wire [0:0] v_7387;
  reg [0:0] v_7388 = 1'h0;
  wire [0:0] v_7389;
  wire [0:0] v_7390;
  wire [0:0] act_7391;
  wire [0:0] v_7392;
  wire [0:0] v_7393;
  wire [0:0] v_7394;
  wire [0:0] vin0_consume_en_7395;
  wire [0:0] vout_canPeek_7395;
  wire [7:0] vout_peek_7395;
  wire [0:0] v_7396;
  wire [0:0] v_7397;
  function [0:0] mux_7397(input [0:0] sel);
    case (sel) 0: mux_7397 = 1'h0; 1: mux_7397 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7398;
  wire [0:0] v_7399;
  wire [0:0] v_7400;
  wire [0:0] v_7401;
  wire [0:0] v_7402;
  function [0:0] mux_7402(input [0:0] sel);
    case (sel) 0: mux_7402 = 1'h0; 1: mux_7402 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7403;
  wire [0:0] vin0_consume_en_7404;
  wire [0:0] vout_canPeek_7404;
  wire [7:0] vout_peek_7404;
  wire [0:0] v_7405;
  wire [0:0] v_7406;
  function [0:0] mux_7406(input [0:0] sel);
    case (sel) 0: mux_7406 = 1'h0; 1: mux_7406 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7407;
  function [0:0] mux_7407(input [0:0] sel);
    case (sel) 0: mux_7407 = 1'h0; 1: mux_7407 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7408;
  wire [0:0] v_7409;
  wire [0:0] v_7410;
  wire [0:0] v_7411;
  wire [0:0] v_7412;
  wire [0:0] v_7413;
  wire [0:0] v_7414;
  function [0:0] mux_7414(input [0:0] sel);
    case (sel) 0: mux_7414 = 1'h0; 1: mux_7414 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7415;
  wire [0:0] v_7416;
  wire [0:0] v_7417;
  wire [0:0] v_7418;
  wire [0:0] v_7419;
  function [0:0] mux_7419(input [0:0] sel);
    case (sel) 0: mux_7419 = 1'h0; 1: mux_7419 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7420;
  wire [0:0] v_7421;
  wire [0:0] v_7422;
  wire [0:0] v_7423;
  function [0:0] mux_7423(input [0:0] sel);
    case (sel) 0: mux_7423 = 1'h0; 1: mux_7423 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7424;
  function [0:0] mux_7424(input [0:0] sel);
    case (sel) 0: mux_7424 = 1'h0; 1: mux_7424 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7425 = 1'h0;
  wire [0:0] v_7426;
  wire [0:0] v_7427;
  wire [0:0] act_7428;
  wire [0:0] v_7429;
  wire [0:0] v_7430;
  wire [0:0] v_7431;
  wire [0:0] vin0_consume_en_7432;
  wire [0:0] vout_canPeek_7432;
  wire [7:0] vout_peek_7432;
  wire [0:0] v_7433;
  wire [0:0] v_7434;
  function [0:0] mux_7434(input [0:0] sel);
    case (sel) 0: mux_7434 = 1'h0; 1: mux_7434 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7435;
  wire [0:0] v_7436;
  wire [0:0] v_7437;
  wire [0:0] v_7438;
  wire [0:0] v_7439;
  function [0:0] mux_7439(input [0:0] sel);
    case (sel) 0: mux_7439 = 1'h0; 1: mux_7439 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7440;
  wire [0:0] vin0_consume_en_7441;
  wire [0:0] vout_canPeek_7441;
  wire [7:0] vout_peek_7441;
  wire [0:0] v_7442;
  wire [0:0] v_7443;
  function [0:0] mux_7443(input [0:0] sel);
    case (sel) 0: mux_7443 = 1'h0; 1: mux_7443 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7444;
  function [0:0] mux_7444(input [0:0] sel);
    case (sel) 0: mux_7444 = 1'h0; 1: mux_7444 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7445;
  wire [0:0] v_7446;
  wire [0:0] v_7447;
  wire [0:0] v_7448;
  wire [0:0] v_7449;
  wire [0:0] v_7450;
  wire [0:0] v_7451;
  function [0:0] mux_7451(input [0:0] sel);
    case (sel) 0: mux_7451 = 1'h0; 1: mux_7451 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7452;
  function [0:0] mux_7452(input [0:0] sel);
    case (sel) 0: mux_7452 = 1'h0; 1: mux_7452 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7453;
  wire [0:0] v_7454;
  wire [0:0] v_7455;
  wire [0:0] v_7456;
  function [0:0] mux_7456(input [0:0] sel);
    case (sel) 0: mux_7456 = 1'h0; 1: mux_7456 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7457;
  function [0:0] mux_7457(input [0:0] sel);
    case (sel) 0: mux_7457 = 1'h0; 1: mux_7457 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7458;
  wire [0:0] v_7459;
  wire [0:0] v_7460;
  wire [0:0] v_7461;
  wire [0:0] v_7462;
  wire [0:0] v_7463;
  function [0:0] mux_7463(input [0:0] sel);
    case (sel) 0: mux_7463 = 1'h0; 1: mux_7463 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7464;
  function [0:0] mux_7464(input [0:0] sel);
    case (sel) 0: mux_7464 = 1'h0; 1: mux_7464 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7465;
  wire [0:0] v_7466;
  wire [0:0] v_7467;
  wire [0:0] v_7468;
  function [0:0] mux_7468(input [0:0] sel);
    case (sel) 0: mux_7468 = 1'h0; 1: mux_7468 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7469;
  function [0:0] mux_7469(input [0:0] sel);
    case (sel) 0: mux_7469 = 1'h0; 1: mux_7469 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7470;
  wire [0:0] v_7471;
  wire [0:0] v_7472;
  wire [0:0] v_7473;
  wire [0:0] v_7474;
  wire [0:0] v_7475;
  function [0:0] mux_7475(input [0:0] sel);
    case (sel) 0: mux_7475 = 1'h0; 1: mux_7475 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7476;
  function [0:0] mux_7476(input [0:0] sel);
    case (sel) 0: mux_7476 = 1'h0; 1: mux_7476 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7477;
  wire [0:0] v_7478;
  wire [0:0] v_7479;
  wire [0:0] v_7480;
  function [0:0] mux_7480(input [0:0] sel);
    case (sel) 0: mux_7480 = 1'h0; 1: mux_7480 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7481;
  function [0:0] mux_7481(input [0:0] sel);
    case (sel) 0: mux_7481 = 1'h0; 1: mux_7481 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7482;
  wire [0:0] v_7483;
  wire [0:0] v_7484;
  wire [0:0] v_7485;
  wire [0:0] v_7486;
  wire [0:0] v_7487;
  function [0:0] mux_7487(input [0:0] sel);
    case (sel) 0: mux_7487 = 1'h0; 1: mux_7487 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7488;
  wire [0:0] v_7489;
  wire [0:0] v_7490;
  wire [0:0] v_7491;
  wire [0:0] v_7492;
  function [0:0] mux_7492(input [0:0] sel);
    case (sel) 0: mux_7492 = 1'h0; 1: mux_7492 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7493;
  wire [0:0] v_7494;
  wire [0:0] v_7495;
  wire [0:0] v_7496;
  function [0:0] mux_7496(input [0:0] sel);
    case (sel) 0: mux_7496 = 1'h0; 1: mux_7496 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7497;
  function [0:0] mux_7497(input [0:0] sel);
    case (sel) 0: mux_7497 = 1'h0; 1: mux_7497 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7498 = 1'h0;
  wire [0:0] v_7499;
  wire [0:0] v_7500;
  wire [0:0] act_7501;
  wire [0:0] v_7502;
  wire [0:0] v_7503;
  wire [0:0] v_7504;
  reg [0:0] v_7505 = 1'h0;
  wire [0:0] v_7506;
  wire [0:0] v_7507;
  wire [0:0] act_7508;
  wire [0:0] v_7509;
  wire [0:0] v_7510;
  wire [0:0] v_7511;
  reg [0:0] v_7512 = 1'h0;
  wire [0:0] v_7513;
  wire [0:0] v_7514;
  wire [0:0] act_7515;
  wire [0:0] v_7516;
  wire [0:0] v_7517;
  wire [0:0] v_7518;
  reg [0:0] v_7519 = 1'h0;
  wire [0:0] v_7520;
  wire [0:0] v_7521;
  wire [0:0] act_7522;
  wire [0:0] v_7523;
  wire [0:0] v_7524;
  wire [0:0] v_7525;
  wire [0:0] vin0_consume_en_7526;
  wire [0:0] vout_canPeek_7526;
  wire [7:0] vout_peek_7526;
  wire [0:0] v_7527;
  wire [0:0] v_7528;
  function [0:0] mux_7528(input [0:0] sel);
    case (sel) 0: mux_7528 = 1'h0; 1: mux_7528 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7529;
  wire [0:0] v_7530;
  wire [0:0] v_7531;
  wire [0:0] v_7532;
  wire [0:0] v_7533;
  function [0:0] mux_7533(input [0:0] sel);
    case (sel) 0: mux_7533 = 1'h0; 1: mux_7533 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7534;
  wire [0:0] vin0_consume_en_7535;
  wire [0:0] vout_canPeek_7535;
  wire [7:0] vout_peek_7535;
  wire [0:0] v_7536;
  wire [0:0] v_7537;
  function [0:0] mux_7537(input [0:0] sel);
    case (sel) 0: mux_7537 = 1'h0; 1: mux_7537 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7538;
  function [0:0] mux_7538(input [0:0] sel);
    case (sel) 0: mux_7538 = 1'h0; 1: mux_7538 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7539;
  wire [0:0] v_7540;
  wire [0:0] v_7541;
  wire [0:0] v_7542;
  wire [0:0] v_7543;
  wire [0:0] v_7544;
  wire [0:0] v_7545;
  function [0:0] mux_7545(input [0:0] sel);
    case (sel) 0: mux_7545 = 1'h0; 1: mux_7545 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7546;
  wire [0:0] v_7547;
  wire [0:0] v_7548;
  wire [0:0] v_7549;
  wire [0:0] v_7550;
  function [0:0] mux_7550(input [0:0] sel);
    case (sel) 0: mux_7550 = 1'h0; 1: mux_7550 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7551;
  wire [0:0] v_7552;
  wire [0:0] v_7553;
  wire [0:0] v_7554;
  function [0:0] mux_7554(input [0:0] sel);
    case (sel) 0: mux_7554 = 1'h0; 1: mux_7554 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7555;
  function [0:0] mux_7555(input [0:0] sel);
    case (sel) 0: mux_7555 = 1'h0; 1: mux_7555 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7556 = 1'h0;
  wire [0:0] v_7557;
  wire [0:0] v_7558;
  wire [0:0] act_7559;
  wire [0:0] v_7560;
  wire [0:0] v_7561;
  wire [0:0] v_7562;
  wire [0:0] vin0_consume_en_7563;
  wire [0:0] vout_canPeek_7563;
  wire [7:0] vout_peek_7563;
  wire [0:0] v_7564;
  wire [0:0] v_7565;
  function [0:0] mux_7565(input [0:0] sel);
    case (sel) 0: mux_7565 = 1'h0; 1: mux_7565 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7566;
  wire [0:0] v_7567;
  wire [0:0] v_7568;
  wire [0:0] v_7569;
  wire [0:0] v_7570;
  function [0:0] mux_7570(input [0:0] sel);
    case (sel) 0: mux_7570 = 1'h0; 1: mux_7570 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7571;
  wire [0:0] vin0_consume_en_7572;
  wire [0:0] vout_canPeek_7572;
  wire [7:0] vout_peek_7572;
  wire [0:0] v_7573;
  wire [0:0] v_7574;
  function [0:0] mux_7574(input [0:0] sel);
    case (sel) 0: mux_7574 = 1'h0; 1: mux_7574 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7575;
  function [0:0] mux_7575(input [0:0] sel);
    case (sel) 0: mux_7575 = 1'h0; 1: mux_7575 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7576;
  wire [0:0] v_7577;
  wire [0:0] v_7578;
  wire [0:0] v_7579;
  wire [0:0] v_7580;
  wire [0:0] v_7581;
  wire [0:0] v_7582;
  function [0:0] mux_7582(input [0:0] sel);
    case (sel) 0: mux_7582 = 1'h0; 1: mux_7582 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7583;
  function [0:0] mux_7583(input [0:0] sel);
    case (sel) 0: mux_7583 = 1'h0; 1: mux_7583 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7584;
  wire [0:0] v_7585;
  wire [0:0] v_7586;
  wire [0:0] v_7587;
  function [0:0] mux_7587(input [0:0] sel);
    case (sel) 0: mux_7587 = 1'h0; 1: mux_7587 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7588;
  function [0:0] mux_7588(input [0:0] sel);
    case (sel) 0: mux_7588 = 1'h0; 1: mux_7588 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7589;
  wire [0:0] v_7590;
  wire [0:0] v_7591;
  wire [0:0] v_7592;
  wire [0:0] v_7593;
  wire [0:0] v_7594;
  function [0:0] mux_7594(input [0:0] sel);
    case (sel) 0: mux_7594 = 1'h0; 1: mux_7594 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7595;
  wire [0:0] v_7596;
  wire [0:0] v_7597;
  wire [0:0] v_7598;
  wire [0:0] v_7599;
  function [0:0] mux_7599(input [0:0] sel);
    case (sel) 0: mux_7599 = 1'h0; 1: mux_7599 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7600;
  wire [0:0] v_7601;
  wire [0:0] v_7602;
  wire [0:0] v_7603;
  function [0:0] mux_7603(input [0:0] sel);
    case (sel) 0: mux_7603 = 1'h0; 1: mux_7603 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7604;
  function [0:0] mux_7604(input [0:0] sel);
    case (sel) 0: mux_7604 = 1'h0; 1: mux_7604 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7605 = 1'h0;
  wire [0:0] v_7606;
  wire [0:0] v_7607;
  wire [0:0] act_7608;
  wire [0:0] v_7609;
  wire [0:0] v_7610;
  wire [0:0] v_7611;
  reg [0:0] v_7612 = 1'h0;
  wire [0:0] v_7613;
  wire [0:0] v_7614;
  wire [0:0] act_7615;
  wire [0:0] v_7616;
  wire [0:0] v_7617;
  wire [0:0] v_7618;
  wire [0:0] vin0_consume_en_7619;
  wire [0:0] vout_canPeek_7619;
  wire [7:0] vout_peek_7619;
  wire [0:0] v_7620;
  wire [0:0] v_7621;
  function [0:0] mux_7621(input [0:0] sel);
    case (sel) 0: mux_7621 = 1'h0; 1: mux_7621 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7622;
  wire [0:0] v_7623;
  wire [0:0] v_7624;
  wire [0:0] v_7625;
  wire [0:0] v_7626;
  function [0:0] mux_7626(input [0:0] sel);
    case (sel) 0: mux_7626 = 1'h0; 1: mux_7626 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7627;
  wire [0:0] vin0_consume_en_7628;
  wire [0:0] vout_canPeek_7628;
  wire [7:0] vout_peek_7628;
  wire [0:0] v_7629;
  wire [0:0] v_7630;
  function [0:0] mux_7630(input [0:0] sel);
    case (sel) 0: mux_7630 = 1'h0; 1: mux_7630 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7631;
  function [0:0] mux_7631(input [0:0] sel);
    case (sel) 0: mux_7631 = 1'h0; 1: mux_7631 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7632;
  wire [0:0] v_7633;
  wire [0:0] v_7634;
  wire [0:0] v_7635;
  wire [0:0] v_7636;
  wire [0:0] v_7637;
  wire [0:0] v_7638;
  function [0:0] mux_7638(input [0:0] sel);
    case (sel) 0: mux_7638 = 1'h0; 1: mux_7638 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7639;
  wire [0:0] v_7640;
  wire [0:0] v_7641;
  wire [0:0] v_7642;
  wire [0:0] v_7643;
  function [0:0] mux_7643(input [0:0] sel);
    case (sel) 0: mux_7643 = 1'h0; 1: mux_7643 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7644;
  wire [0:0] v_7645;
  wire [0:0] v_7646;
  wire [0:0] v_7647;
  function [0:0] mux_7647(input [0:0] sel);
    case (sel) 0: mux_7647 = 1'h0; 1: mux_7647 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7648;
  function [0:0] mux_7648(input [0:0] sel);
    case (sel) 0: mux_7648 = 1'h0; 1: mux_7648 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7649 = 1'h0;
  wire [0:0] v_7650;
  wire [0:0] v_7651;
  wire [0:0] act_7652;
  wire [0:0] v_7653;
  wire [0:0] v_7654;
  wire [0:0] v_7655;
  wire [0:0] vin0_consume_en_7656;
  wire [0:0] vout_canPeek_7656;
  wire [7:0] vout_peek_7656;
  wire [0:0] v_7657;
  wire [0:0] v_7658;
  function [0:0] mux_7658(input [0:0] sel);
    case (sel) 0: mux_7658 = 1'h0; 1: mux_7658 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7659;
  wire [0:0] v_7660;
  wire [0:0] v_7661;
  wire [0:0] v_7662;
  wire [0:0] v_7663;
  function [0:0] mux_7663(input [0:0] sel);
    case (sel) 0: mux_7663 = 1'h0; 1: mux_7663 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7664;
  wire [0:0] vin0_consume_en_7665;
  wire [0:0] vout_canPeek_7665;
  wire [7:0] vout_peek_7665;
  wire [0:0] v_7666;
  wire [0:0] v_7667;
  function [0:0] mux_7667(input [0:0] sel);
    case (sel) 0: mux_7667 = 1'h0; 1: mux_7667 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7668;
  function [0:0] mux_7668(input [0:0] sel);
    case (sel) 0: mux_7668 = 1'h0; 1: mux_7668 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7669;
  wire [0:0] v_7670;
  wire [0:0] v_7671;
  wire [0:0] v_7672;
  wire [0:0] v_7673;
  wire [0:0] v_7674;
  wire [0:0] v_7675;
  function [0:0] mux_7675(input [0:0] sel);
    case (sel) 0: mux_7675 = 1'h0; 1: mux_7675 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7676;
  function [0:0] mux_7676(input [0:0] sel);
    case (sel) 0: mux_7676 = 1'h0; 1: mux_7676 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7677;
  wire [0:0] v_7678;
  wire [0:0] v_7679;
  wire [0:0] v_7680;
  function [0:0] mux_7680(input [0:0] sel);
    case (sel) 0: mux_7680 = 1'h0; 1: mux_7680 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7681;
  function [0:0] mux_7681(input [0:0] sel);
    case (sel) 0: mux_7681 = 1'h0; 1: mux_7681 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7682;
  wire [0:0] v_7683;
  wire [0:0] v_7684;
  wire [0:0] v_7685;
  wire [0:0] v_7686;
  wire [0:0] v_7687;
  function [0:0] mux_7687(input [0:0] sel);
    case (sel) 0: mux_7687 = 1'h0; 1: mux_7687 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7688;
  function [0:0] mux_7688(input [0:0] sel);
    case (sel) 0: mux_7688 = 1'h0; 1: mux_7688 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7689;
  wire [0:0] v_7690;
  wire [0:0] v_7691;
  wire [0:0] v_7692;
  function [0:0] mux_7692(input [0:0] sel);
    case (sel) 0: mux_7692 = 1'h0; 1: mux_7692 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7693;
  function [0:0] mux_7693(input [0:0] sel);
    case (sel) 0: mux_7693 = 1'h0; 1: mux_7693 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7694;
  wire [0:0] v_7695;
  wire [0:0] v_7696;
  wire [0:0] v_7697;
  wire [0:0] v_7698;
  wire [0:0] v_7699;
  function [0:0] mux_7699(input [0:0] sel);
    case (sel) 0: mux_7699 = 1'h0; 1: mux_7699 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7700;
  wire [0:0] v_7701;
  wire [0:0] v_7702;
  wire [0:0] v_7703;
  wire [0:0] v_7704;
  function [0:0] mux_7704(input [0:0] sel);
    case (sel) 0: mux_7704 = 1'h0; 1: mux_7704 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7705;
  wire [0:0] v_7706;
  wire [0:0] v_7707;
  wire [0:0] v_7708;
  function [0:0] mux_7708(input [0:0] sel);
    case (sel) 0: mux_7708 = 1'h0; 1: mux_7708 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7709;
  function [0:0] mux_7709(input [0:0] sel);
    case (sel) 0: mux_7709 = 1'h0; 1: mux_7709 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7710 = 1'h0;
  wire [0:0] v_7711;
  wire [0:0] v_7712;
  wire [0:0] act_7713;
  wire [0:0] v_7714;
  wire [0:0] v_7715;
  wire [0:0] v_7716;
  reg [0:0] v_7717 = 1'h0;
  wire [0:0] v_7718;
  wire [0:0] v_7719;
  wire [0:0] act_7720;
  wire [0:0] v_7721;
  wire [0:0] v_7722;
  wire [0:0] v_7723;
  reg [0:0] v_7724 = 1'h0;
  wire [0:0] v_7725;
  wire [0:0] v_7726;
  wire [0:0] act_7727;
  wire [0:0] v_7728;
  wire [0:0] v_7729;
  wire [0:0] v_7730;
  wire [0:0] vin0_consume_en_7731;
  wire [0:0] vout_canPeek_7731;
  wire [7:0] vout_peek_7731;
  wire [0:0] v_7732;
  wire [0:0] v_7733;
  function [0:0] mux_7733(input [0:0] sel);
    case (sel) 0: mux_7733 = 1'h0; 1: mux_7733 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7734;
  wire [0:0] v_7735;
  wire [0:0] v_7736;
  wire [0:0] v_7737;
  wire [0:0] v_7738;
  function [0:0] mux_7738(input [0:0] sel);
    case (sel) 0: mux_7738 = 1'h0; 1: mux_7738 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7739;
  wire [0:0] vin0_consume_en_7740;
  wire [0:0] vout_canPeek_7740;
  wire [7:0] vout_peek_7740;
  wire [0:0] v_7741;
  wire [0:0] v_7742;
  function [0:0] mux_7742(input [0:0] sel);
    case (sel) 0: mux_7742 = 1'h0; 1: mux_7742 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7743;
  function [0:0] mux_7743(input [0:0] sel);
    case (sel) 0: mux_7743 = 1'h0; 1: mux_7743 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7744;
  wire [0:0] v_7745;
  wire [0:0] v_7746;
  wire [0:0] v_7747;
  wire [0:0] v_7748;
  wire [0:0] v_7749;
  wire [0:0] v_7750;
  function [0:0] mux_7750(input [0:0] sel);
    case (sel) 0: mux_7750 = 1'h0; 1: mux_7750 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7751;
  wire [0:0] v_7752;
  wire [0:0] v_7753;
  wire [0:0] v_7754;
  wire [0:0] v_7755;
  function [0:0] mux_7755(input [0:0] sel);
    case (sel) 0: mux_7755 = 1'h0; 1: mux_7755 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7756;
  wire [0:0] v_7757;
  wire [0:0] v_7758;
  wire [0:0] v_7759;
  function [0:0] mux_7759(input [0:0] sel);
    case (sel) 0: mux_7759 = 1'h0; 1: mux_7759 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7760;
  function [0:0] mux_7760(input [0:0] sel);
    case (sel) 0: mux_7760 = 1'h0; 1: mux_7760 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7761 = 1'h0;
  wire [0:0] v_7762;
  wire [0:0] v_7763;
  wire [0:0] act_7764;
  wire [0:0] v_7765;
  wire [0:0] v_7766;
  wire [0:0] v_7767;
  wire [0:0] vin0_consume_en_7768;
  wire [0:0] vout_canPeek_7768;
  wire [7:0] vout_peek_7768;
  wire [0:0] v_7769;
  wire [0:0] v_7770;
  function [0:0] mux_7770(input [0:0] sel);
    case (sel) 0: mux_7770 = 1'h0; 1: mux_7770 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7771;
  wire [0:0] v_7772;
  wire [0:0] v_7773;
  wire [0:0] v_7774;
  wire [0:0] v_7775;
  function [0:0] mux_7775(input [0:0] sel);
    case (sel) 0: mux_7775 = 1'h0; 1: mux_7775 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7776;
  wire [0:0] vin0_consume_en_7777;
  wire [0:0] vout_canPeek_7777;
  wire [7:0] vout_peek_7777;
  wire [0:0] v_7778;
  wire [0:0] v_7779;
  function [0:0] mux_7779(input [0:0] sel);
    case (sel) 0: mux_7779 = 1'h0; 1: mux_7779 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7780;
  function [0:0] mux_7780(input [0:0] sel);
    case (sel) 0: mux_7780 = 1'h0; 1: mux_7780 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7781;
  wire [0:0] v_7782;
  wire [0:0] v_7783;
  wire [0:0] v_7784;
  wire [0:0] v_7785;
  wire [0:0] v_7786;
  wire [0:0] v_7787;
  function [0:0] mux_7787(input [0:0] sel);
    case (sel) 0: mux_7787 = 1'h0; 1: mux_7787 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7788;
  function [0:0] mux_7788(input [0:0] sel);
    case (sel) 0: mux_7788 = 1'h0; 1: mux_7788 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7789;
  wire [0:0] v_7790;
  wire [0:0] v_7791;
  wire [0:0] v_7792;
  function [0:0] mux_7792(input [0:0] sel);
    case (sel) 0: mux_7792 = 1'h0; 1: mux_7792 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7793;
  function [0:0] mux_7793(input [0:0] sel);
    case (sel) 0: mux_7793 = 1'h0; 1: mux_7793 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7794;
  wire [0:0] v_7795;
  wire [0:0] v_7796;
  wire [0:0] v_7797;
  wire [0:0] v_7798;
  wire [0:0] v_7799;
  function [0:0] mux_7799(input [0:0] sel);
    case (sel) 0: mux_7799 = 1'h0; 1: mux_7799 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7800;
  wire [0:0] v_7801;
  wire [0:0] v_7802;
  wire [0:0] v_7803;
  wire [0:0] v_7804;
  function [0:0] mux_7804(input [0:0] sel);
    case (sel) 0: mux_7804 = 1'h0; 1: mux_7804 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7805;
  wire [0:0] v_7806;
  wire [0:0] v_7807;
  wire [0:0] v_7808;
  function [0:0] mux_7808(input [0:0] sel);
    case (sel) 0: mux_7808 = 1'h0; 1: mux_7808 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7809;
  function [0:0] mux_7809(input [0:0] sel);
    case (sel) 0: mux_7809 = 1'h0; 1: mux_7809 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7810 = 1'h0;
  wire [0:0] v_7811;
  wire [0:0] v_7812;
  wire [0:0] act_7813;
  wire [0:0] v_7814;
  wire [0:0] v_7815;
  wire [0:0] v_7816;
  reg [0:0] v_7817 = 1'h0;
  wire [0:0] v_7818;
  wire [0:0] v_7819;
  wire [0:0] act_7820;
  wire [0:0] v_7821;
  wire [0:0] v_7822;
  wire [0:0] v_7823;
  wire [0:0] vin0_consume_en_7824;
  wire [0:0] vout_canPeek_7824;
  wire [7:0] vout_peek_7824;
  wire [0:0] v_7825;
  wire [0:0] v_7826;
  function [0:0] mux_7826(input [0:0] sel);
    case (sel) 0: mux_7826 = 1'h0; 1: mux_7826 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7827;
  wire [0:0] v_7828;
  wire [0:0] v_7829;
  wire [0:0] v_7830;
  wire [0:0] v_7831;
  function [0:0] mux_7831(input [0:0] sel);
    case (sel) 0: mux_7831 = 1'h0; 1: mux_7831 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7832;
  wire [0:0] vin0_consume_en_7833;
  wire [0:0] vout_canPeek_7833;
  wire [7:0] vout_peek_7833;
  wire [0:0] v_7834;
  wire [0:0] v_7835;
  function [0:0] mux_7835(input [0:0] sel);
    case (sel) 0: mux_7835 = 1'h0; 1: mux_7835 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7836;
  function [0:0] mux_7836(input [0:0] sel);
    case (sel) 0: mux_7836 = 1'h0; 1: mux_7836 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7837;
  wire [0:0] v_7838;
  wire [0:0] v_7839;
  wire [0:0] v_7840;
  wire [0:0] v_7841;
  wire [0:0] v_7842;
  wire [0:0] v_7843;
  function [0:0] mux_7843(input [0:0] sel);
    case (sel) 0: mux_7843 = 1'h0; 1: mux_7843 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7844;
  wire [0:0] v_7845;
  wire [0:0] v_7846;
  wire [0:0] v_7847;
  wire [0:0] v_7848;
  function [0:0] mux_7848(input [0:0] sel);
    case (sel) 0: mux_7848 = 1'h0; 1: mux_7848 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7849;
  wire [0:0] v_7850;
  wire [0:0] v_7851;
  wire [0:0] v_7852;
  function [0:0] mux_7852(input [0:0] sel);
    case (sel) 0: mux_7852 = 1'h0; 1: mux_7852 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7853;
  function [0:0] mux_7853(input [0:0] sel);
    case (sel) 0: mux_7853 = 1'h0; 1: mux_7853 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7854 = 1'h0;
  wire [0:0] v_7855;
  wire [0:0] v_7856;
  wire [0:0] act_7857;
  wire [0:0] v_7858;
  wire [0:0] v_7859;
  wire [0:0] v_7860;
  wire [0:0] vin0_consume_en_7861;
  wire [0:0] vout_canPeek_7861;
  wire [7:0] vout_peek_7861;
  wire [0:0] v_7862;
  wire [0:0] v_7863;
  function [0:0] mux_7863(input [0:0] sel);
    case (sel) 0: mux_7863 = 1'h0; 1: mux_7863 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7864;
  wire [0:0] v_7865;
  wire [0:0] v_7866;
  wire [0:0] v_7867;
  wire [0:0] v_7868;
  function [0:0] mux_7868(input [0:0] sel);
    case (sel) 0: mux_7868 = 1'h0; 1: mux_7868 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7869;
  wire [0:0] vin0_consume_en_7870;
  wire [0:0] vout_canPeek_7870;
  wire [7:0] vout_peek_7870;
  wire [0:0] v_7871;
  wire [0:0] v_7872;
  function [0:0] mux_7872(input [0:0] sel);
    case (sel) 0: mux_7872 = 1'h0; 1: mux_7872 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7873;
  function [0:0] mux_7873(input [0:0] sel);
    case (sel) 0: mux_7873 = 1'h0; 1: mux_7873 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7874;
  wire [0:0] v_7875;
  wire [0:0] v_7876;
  wire [0:0] v_7877;
  wire [0:0] v_7878;
  wire [0:0] v_7879;
  wire [0:0] v_7880;
  function [0:0] mux_7880(input [0:0] sel);
    case (sel) 0: mux_7880 = 1'h0; 1: mux_7880 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7881;
  function [0:0] mux_7881(input [0:0] sel);
    case (sel) 0: mux_7881 = 1'h0; 1: mux_7881 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7882;
  wire [0:0] v_7883;
  wire [0:0] v_7884;
  wire [0:0] v_7885;
  function [0:0] mux_7885(input [0:0] sel);
    case (sel) 0: mux_7885 = 1'h0; 1: mux_7885 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7886;
  function [0:0] mux_7886(input [0:0] sel);
    case (sel) 0: mux_7886 = 1'h0; 1: mux_7886 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7887;
  wire [0:0] v_7888;
  wire [0:0] v_7889;
  wire [0:0] v_7890;
  wire [0:0] v_7891;
  wire [0:0] v_7892;
  function [0:0] mux_7892(input [0:0] sel);
    case (sel) 0: mux_7892 = 1'h0; 1: mux_7892 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7893;
  function [0:0] mux_7893(input [0:0] sel);
    case (sel) 0: mux_7893 = 1'h0; 1: mux_7893 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7894;
  wire [0:0] v_7895;
  wire [0:0] v_7896;
  wire [0:0] v_7897;
  function [0:0] mux_7897(input [0:0] sel);
    case (sel) 0: mux_7897 = 1'h0; 1: mux_7897 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7898;
  function [0:0] mux_7898(input [0:0] sel);
    case (sel) 0: mux_7898 = 1'h0; 1: mux_7898 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7899;
  wire [0:0] v_7900;
  wire [0:0] v_7901;
  wire [0:0] v_7902;
  wire [0:0] v_7903;
  wire [0:0] v_7904;
  function [0:0] mux_7904(input [0:0] sel);
    case (sel) 0: mux_7904 = 1'h0; 1: mux_7904 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7905;
  function [0:0] mux_7905(input [0:0] sel);
    case (sel) 0: mux_7905 = 1'h0; 1: mux_7905 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7906;
  wire [0:0] v_7907;
  wire [0:0] v_7908;
  wire [0:0] v_7909;
  function [0:0] mux_7909(input [0:0] sel);
    case (sel) 0: mux_7909 = 1'h0; 1: mux_7909 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7910;
  function [0:0] mux_7910(input [0:0] sel);
    case (sel) 0: mux_7910 = 1'h0; 1: mux_7910 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7911;
  wire [0:0] v_7912;
  wire [0:0] v_7913;
  wire [0:0] v_7914;
  wire [0:0] v_7915;
  wire [0:0] v_7916;
  function [0:0] mux_7916(input [0:0] sel);
    case (sel) 0: mux_7916 = 1'h0; 1: mux_7916 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7917;
  function [0:0] mux_7917(input [0:0] sel);
    case (sel) 0: mux_7917 = 1'h0; 1: mux_7917 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7918;
  wire [0:0] v_7919;
  wire [0:0] v_7920;
  wire [0:0] v_7921;
  function [0:0] mux_7921(input [0:0] sel);
    case (sel) 0: mux_7921 = 1'h0; 1: mux_7921 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7922;
  function [0:0] mux_7922(input [0:0] sel);
    case (sel) 0: mux_7922 = 1'h0; 1: mux_7922 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7923;
  wire [0:0] v_7924;
  wire [0:0] v_7925;
  wire [0:0] v_7926;
  wire [0:0] v_7927;
  wire [0:0] v_7928;
  function [0:0] mux_7928(input [0:0] sel);
    case (sel) 0: mux_7928 = 1'h0; 1: mux_7928 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7929;
  function [0:0] mux_7929(input [0:0] sel);
    case (sel) 0: mux_7929 = 1'h0; 1: mux_7929 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7930;
  wire [0:0] v_7931;
  wire [0:0] v_7932;
  wire [0:0] v_7933;
  function [0:0] mux_7933(input [0:0] sel);
    case (sel) 0: mux_7933 = 1'h0; 1: mux_7933 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7934;
  function [0:0] mux_7934(input [0:0] sel);
    case (sel) 0: mux_7934 = 1'h0; 1: mux_7934 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7935;
  wire [0:0] v_7936;
  wire [0:0] v_7937;
  wire [0:0] v_7938;
  wire [0:0] v_7939;
  wire [0:0] v_7940;
  function [0:0] mux_7940(input [0:0] sel);
    case (sel) 0: mux_7940 = 1'h0; 1: mux_7940 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7941;
  function [0:0] mux_7941(input [0:0] sel);
    case (sel) 0: mux_7941 = 1'h0; 1: mux_7941 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7942;
  wire [0:0] v_7943;
  wire [0:0] v_7944;
  wire [0:0] v_7945;
  function [0:0] mux_7945(input [0:0] sel);
    case (sel) 0: mux_7945 = 1'h0; 1: mux_7945 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7946;
  function [0:0] mux_7946(input [0:0] sel);
    case (sel) 0: mux_7946 = 1'h0; 1: mux_7946 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7947;
  wire [0:0] v_7948;
  wire [0:0] v_7949;
  wire [0:0] v_7950;
  wire [0:0] v_7951;
  wire [0:0] v_7952;
  function [0:0] mux_7952(input [0:0] sel);
    case (sel) 0: mux_7952 = 1'h0; 1: mux_7952 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7953;
  wire [0:0] v_7954;
  wire [0:0] v_7955;
  wire [0:0] v_7956;
  reg [0:0] v_7957 = 1'h0;
  wire [0:0] v_7958;
  wire [0:0] v_7959;
  wire [0:0] act_7960;
  wire [0:0] v_7961;
  wire [0:0] v_7962;
  wire [0:0] v_7963;
  wire [0:0] v_7964;
  wire [0:0] v_7965;
  wire [0:0] v_7966;
  function [0:0] mux_7966(input [0:0] sel);
    case (sel) 0: mux_7966 = 1'h0; 1: mux_7966 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7967;
  wire [0:0] v_7968;
  wire [0:0] v_7969;
  wire [0:0] v_7970;
  reg [0:0] v_7971 = 1'h0;
  wire [0:0] v_7972;
  wire [0:0] v_7973;
  wire [0:0] act_7974;
  wire [0:0] v_7975;
  wire [0:0] v_7976;
  wire [0:0] v_7977;
  reg [0:0] v_7978 = 1'h0;
  wire [0:0] v_7979;
  wire [0:0] v_7980;
  wire [0:0] act_7981;
  wire [0:0] v_7982;
  wire [0:0] v_7983;
  wire [0:0] v_7984;
  reg [0:0] v_7985 = 1'h0;
  wire [0:0] v_7986;
  wire [0:0] v_7987;
  wire [0:0] act_7988;
  wire [0:0] v_7989;
  wire [0:0] v_7990;
  wire [0:0] v_7991;
  reg [0:0] v_7992 = 1'h0;
  wire [0:0] v_7993;
  wire [0:0] v_7994;
  wire [0:0] act_7995;
  wire [0:0] v_7996;
  wire [0:0] v_7997;
  wire [0:0] v_7998;
  reg [0:0] v_7999 = 1'h0;
  wire [0:0] v_8000;
  wire [0:0] v_8001;
  wire [0:0] act_8002;
  wire [0:0] v_8003;
  wire [0:0] v_8004;
  wire [0:0] v_8005;
  reg [0:0] v_8006 = 1'h0;
  wire [0:0] v_8007;
  wire [0:0] v_8008;
  wire [0:0] act_8009;
  wire [0:0] v_8010;
  wire [0:0] v_8011;
  wire [0:0] v_8012;
  reg [0:0] v_8013 = 1'h0;
  wire [0:0] v_8014;
  wire [0:0] v_8015;
  wire [0:0] act_8016;
  wire [0:0] v_8017;
  wire [0:0] v_8018;
  wire [0:0] v_8019;
  reg [0:0] v_8020 = 1'h0;
  wire [0:0] v_8021;
  wire [0:0] v_8022;
  wire [0:0] act_8023;
  wire [0:0] v_8024;
  wire [0:0] v_8025;
  wire [0:0] v_8026;
  reg [0:0] v_8027 = 1'h0;
  wire [0:0] v_8028;
  wire [0:0] v_8029;
  wire [0:0] act_8030;
  wire [0:0] v_8031;
  wire [0:0] v_8032;
  wire [0:0] v_8033;
  reg [0:0] v_8034 = 1'h0;
  wire [0:0] v_8035;
  wire [0:0] v_8036;
  wire [0:0] act_8037;
  wire [0:0] v_8038;
  wire [0:0] v_8039;
  wire [0:0] v_8040;
  wire [0:0] vin0_consume_en_8041;
  wire [0:0] vout_canPeek_8041;
  wire [7:0] vout_peek_8041;
  wire [0:0] v_8042;
  wire [0:0] v_8043;
  function [0:0] mux_8043(input [0:0] sel);
    case (sel) 0: mux_8043 = 1'h0; 1: mux_8043 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8044;
  wire [0:0] v_8045;
  wire [0:0] v_8046;
  wire [0:0] v_8047;
  wire [0:0] v_8048;
  function [0:0] mux_8048(input [0:0] sel);
    case (sel) 0: mux_8048 = 1'h0; 1: mux_8048 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8049;
  wire [0:0] vin0_consume_en_8050;
  wire [0:0] vout_canPeek_8050;
  wire [7:0] vout_peek_8050;
  wire [0:0] v_8051;
  wire [0:0] v_8052;
  function [0:0] mux_8052(input [0:0] sel);
    case (sel) 0: mux_8052 = 1'h0; 1: mux_8052 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8053;
  function [0:0] mux_8053(input [0:0] sel);
    case (sel) 0: mux_8053 = 1'h0; 1: mux_8053 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8054;
  wire [0:0] v_8055;
  wire [0:0] v_8056;
  wire [0:0] v_8057;
  wire [0:0] v_8058;
  wire [0:0] v_8059;
  wire [0:0] v_8060;
  function [0:0] mux_8060(input [0:0] sel);
    case (sel) 0: mux_8060 = 1'h0; 1: mux_8060 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8061;
  wire [0:0] v_8062;
  wire [0:0] v_8063;
  wire [0:0] v_8064;
  wire [0:0] v_8065;
  function [0:0] mux_8065(input [0:0] sel);
    case (sel) 0: mux_8065 = 1'h0; 1: mux_8065 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8066;
  wire [0:0] v_8067;
  wire [0:0] v_8068;
  wire [0:0] v_8069;
  function [0:0] mux_8069(input [0:0] sel);
    case (sel) 0: mux_8069 = 1'h0; 1: mux_8069 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8070;
  function [0:0] mux_8070(input [0:0] sel);
    case (sel) 0: mux_8070 = 1'h0; 1: mux_8070 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8071 = 1'h0;
  wire [0:0] v_8072;
  wire [0:0] v_8073;
  wire [0:0] act_8074;
  wire [0:0] v_8075;
  wire [0:0] v_8076;
  wire [0:0] v_8077;
  wire [0:0] vin0_consume_en_8078;
  wire [0:0] vout_canPeek_8078;
  wire [7:0] vout_peek_8078;
  wire [0:0] v_8079;
  wire [0:0] v_8080;
  function [0:0] mux_8080(input [0:0] sel);
    case (sel) 0: mux_8080 = 1'h0; 1: mux_8080 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8081;
  wire [0:0] v_8082;
  wire [0:0] v_8083;
  wire [0:0] v_8084;
  wire [0:0] v_8085;
  function [0:0] mux_8085(input [0:0] sel);
    case (sel) 0: mux_8085 = 1'h0; 1: mux_8085 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8086;
  wire [0:0] vin0_consume_en_8087;
  wire [0:0] vout_canPeek_8087;
  wire [7:0] vout_peek_8087;
  wire [0:0] v_8088;
  wire [0:0] v_8089;
  function [0:0] mux_8089(input [0:0] sel);
    case (sel) 0: mux_8089 = 1'h0; 1: mux_8089 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8090;
  function [0:0] mux_8090(input [0:0] sel);
    case (sel) 0: mux_8090 = 1'h0; 1: mux_8090 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8091;
  wire [0:0] v_8092;
  wire [0:0] v_8093;
  wire [0:0] v_8094;
  wire [0:0] v_8095;
  wire [0:0] v_8096;
  wire [0:0] v_8097;
  function [0:0] mux_8097(input [0:0] sel);
    case (sel) 0: mux_8097 = 1'h0; 1: mux_8097 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8098;
  function [0:0] mux_8098(input [0:0] sel);
    case (sel) 0: mux_8098 = 1'h0; 1: mux_8098 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8099;
  wire [0:0] v_8100;
  wire [0:0] v_8101;
  wire [0:0] v_8102;
  function [0:0] mux_8102(input [0:0] sel);
    case (sel) 0: mux_8102 = 1'h0; 1: mux_8102 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8103;
  function [0:0] mux_8103(input [0:0] sel);
    case (sel) 0: mux_8103 = 1'h0; 1: mux_8103 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8104;
  wire [0:0] v_8105;
  wire [0:0] v_8106;
  wire [0:0] v_8107;
  wire [0:0] v_8108;
  wire [0:0] v_8109;
  function [0:0] mux_8109(input [0:0] sel);
    case (sel) 0: mux_8109 = 1'h0; 1: mux_8109 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8110;
  wire [0:0] v_8111;
  wire [0:0] v_8112;
  wire [0:0] v_8113;
  wire [0:0] v_8114;
  function [0:0] mux_8114(input [0:0] sel);
    case (sel) 0: mux_8114 = 1'h0; 1: mux_8114 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8115;
  wire [0:0] v_8116;
  wire [0:0] v_8117;
  wire [0:0] v_8118;
  function [0:0] mux_8118(input [0:0] sel);
    case (sel) 0: mux_8118 = 1'h0; 1: mux_8118 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8119;
  function [0:0] mux_8119(input [0:0] sel);
    case (sel) 0: mux_8119 = 1'h0; 1: mux_8119 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8120 = 1'h0;
  wire [0:0] v_8121;
  wire [0:0] v_8122;
  wire [0:0] act_8123;
  wire [0:0] v_8124;
  wire [0:0] v_8125;
  wire [0:0] v_8126;
  reg [0:0] v_8127 = 1'h0;
  wire [0:0] v_8128;
  wire [0:0] v_8129;
  wire [0:0] act_8130;
  wire [0:0] v_8131;
  wire [0:0] v_8132;
  wire [0:0] v_8133;
  wire [0:0] vin0_consume_en_8134;
  wire [0:0] vout_canPeek_8134;
  wire [7:0] vout_peek_8134;
  wire [0:0] v_8135;
  wire [0:0] v_8136;
  function [0:0] mux_8136(input [0:0] sel);
    case (sel) 0: mux_8136 = 1'h0; 1: mux_8136 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8137;
  wire [0:0] v_8138;
  wire [0:0] v_8139;
  wire [0:0] v_8140;
  wire [0:0] v_8141;
  function [0:0] mux_8141(input [0:0] sel);
    case (sel) 0: mux_8141 = 1'h0; 1: mux_8141 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8142;
  wire [0:0] vin0_consume_en_8143;
  wire [0:0] vout_canPeek_8143;
  wire [7:0] vout_peek_8143;
  wire [0:0] v_8144;
  wire [0:0] v_8145;
  function [0:0] mux_8145(input [0:0] sel);
    case (sel) 0: mux_8145 = 1'h0; 1: mux_8145 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8146;
  function [0:0] mux_8146(input [0:0] sel);
    case (sel) 0: mux_8146 = 1'h0; 1: mux_8146 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8147;
  wire [0:0] v_8148;
  wire [0:0] v_8149;
  wire [0:0] v_8150;
  wire [0:0] v_8151;
  wire [0:0] v_8152;
  wire [0:0] v_8153;
  function [0:0] mux_8153(input [0:0] sel);
    case (sel) 0: mux_8153 = 1'h0; 1: mux_8153 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8154;
  wire [0:0] v_8155;
  wire [0:0] v_8156;
  wire [0:0] v_8157;
  wire [0:0] v_8158;
  function [0:0] mux_8158(input [0:0] sel);
    case (sel) 0: mux_8158 = 1'h0; 1: mux_8158 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8159;
  wire [0:0] v_8160;
  wire [0:0] v_8161;
  wire [0:0] v_8162;
  function [0:0] mux_8162(input [0:0] sel);
    case (sel) 0: mux_8162 = 1'h0; 1: mux_8162 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8163;
  function [0:0] mux_8163(input [0:0] sel);
    case (sel) 0: mux_8163 = 1'h0; 1: mux_8163 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8164 = 1'h0;
  wire [0:0] v_8165;
  wire [0:0] v_8166;
  wire [0:0] act_8167;
  wire [0:0] v_8168;
  wire [0:0] v_8169;
  wire [0:0] v_8170;
  wire [0:0] vin0_consume_en_8171;
  wire [0:0] vout_canPeek_8171;
  wire [7:0] vout_peek_8171;
  wire [0:0] v_8172;
  wire [0:0] v_8173;
  function [0:0] mux_8173(input [0:0] sel);
    case (sel) 0: mux_8173 = 1'h0; 1: mux_8173 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8174;
  wire [0:0] v_8175;
  wire [0:0] v_8176;
  wire [0:0] v_8177;
  wire [0:0] v_8178;
  function [0:0] mux_8178(input [0:0] sel);
    case (sel) 0: mux_8178 = 1'h0; 1: mux_8178 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8179;
  wire [0:0] vin0_consume_en_8180;
  wire [0:0] vout_canPeek_8180;
  wire [7:0] vout_peek_8180;
  wire [0:0] v_8181;
  wire [0:0] v_8182;
  function [0:0] mux_8182(input [0:0] sel);
    case (sel) 0: mux_8182 = 1'h0; 1: mux_8182 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8183;
  function [0:0] mux_8183(input [0:0] sel);
    case (sel) 0: mux_8183 = 1'h0; 1: mux_8183 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8184;
  wire [0:0] v_8185;
  wire [0:0] v_8186;
  wire [0:0] v_8187;
  wire [0:0] v_8188;
  wire [0:0] v_8189;
  wire [0:0] v_8190;
  function [0:0] mux_8190(input [0:0] sel);
    case (sel) 0: mux_8190 = 1'h0; 1: mux_8190 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8191;
  function [0:0] mux_8191(input [0:0] sel);
    case (sel) 0: mux_8191 = 1'h0; 1: mux_8191 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8192;
  wire [0:0] v_8193;
  wire [0:0] v_8194;
  wire [0:0] v_8195;
  function [0:0] mux_8195(input [0:0] sel);
    case (sel) 0: mux_8195 = 1'h0; 1: mux_8195 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8196;
  function [0:0] mux_8196(input [0:0] sel);
    case (sel) 0: mux_8196 = 1'h0; 1: mux_8196 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8197;
  wire [0:0] v_8198;
  wire [0:0] v_8199;
  wire [0:0] v_8200;
  wire [0:0] v_8201;
  wire [0:0] v_8202;
  function [0:0] mux_8202(input [0:0] sel);
    case (sel) 0: mux_8202 = 1'h0; 1: mux_8202 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8203;
  function [0:0] mux_8203(input [0:0] sel);
    case (sel) 0: mux_8203 = 1'h0; 1: mux_8203 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8204;
  wire [0:0] v_8205;
  wire [0:0] v_8206;
  wire [0:0] v_8207;
  function [0:0] mux_8207(input [0:0] sel);
    case (sel) 0: mux_8207 = 1'h0; 1: mux_8207 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8208;
  function [0:0] mux_8208(input [0:0] sel);
    case (sel) 0: mux_8208 = 1'h0; 1: mux_8208 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8209;
  wire [0:0] v_8210;
  wire [0:0] v_8211;
  wire [0:0] v_8212;
  wire [0:0] v_8213;
  wire [0:0] v_8214;
  function [0:0] mux_8214(input [0:0] sel);
    case (sel) 0: mux_8214 = 1'h0; 1: mux_8214 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8215;
  wire [0:0] v_8216;
  wire [0:0] v_8217;
  wire [0:0] v_8218;
  wire [0:0] v_8219;
  function [0:0] mux_8219(input [0:0] sel);
    case (sel) 0: mux_8219 = 1'h0; 1: mux_8219 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8220;
  wire [0:0] v_8221;
  wire [0:0] v_8222;
  wire [0:0] v_8223;
  function [0:0] mux_8223(input [0:0] sel);
    case (sel) 0: mux_8223 = 1'h0; 1: mux_8223 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8224;
  function [0:0] mux_8224(input [0:0] sel);
    case (sel) 0: mux_8224 = 1'h0; 1: mux_8224 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8225 = 1'h0;
  wire [0:0] v_8226;
  wire [0:0] v_8227;
  wire [0:0] act_8228;
  wire [0:0] v_8229;
  wire [0:0] v_8230;
  wire [0:0] v_8231;
  reg [0:0] v_8232 = 1'h0;
  wire [0:0] v_8233;
  wire [0:0] v_8234;
  wire [0:0] act_8235;
  wire [0:0] v_8236;
  wire [0:0] v_8237;
  wire [0:0] v_8238;
  reg [0:0] v_8239 = 1'h0;
  wire [0:0] v_8240;
  wire [0:0] v_8241;
  wire [0:0] act_8242;
  wire [0:0] v_8243;
  wire [0:0] v_8244;
  wire [0:0] v_8245;
  wire [0:0] vin0_consume_en_8246;
  wire [0:0] vout_canPeek_8246;
  wire [7:0] vout_peek_8246;
  wire [0:0] v_8247;
  wire [0:0] v_8248;
  function [0:0] mux_8248(input [0:0] sel);
    case (sel) 0: mux_8248 = 1'h0; 1: mux_8248 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8249;
  wire [0:0] v_8250;
  wire [0:0] v_8251;
  wire [0:0] v_8252;
  wire [0:0] v_8253;
  function [0:0] mux_8253(input [0:0] sel);
    case (sel) 0: mux_8253 = 1'h0; 1: mux_8253 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8254;
  wire [0:0] vin0_consume_en_8255;
  wire [0:0] vout_canPeek_8255;
  wire [7:0] vout_peek_8255;
  wire [0:0] v_8256;
  wire [0:0] v_8257;
  function [0:0] mux_8257(input [0:0] sel);
    case (sel) 0: mux_8257 = 1'h0; 1: mux_8257 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8258;
  function [0:0] mux_8258(input [0:0] sel);
    case (sel) 0: mux_8258 = 1'h0; 1: mux_8258 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8259;
  wire [0:0] v_8260;
  wire [0:0] v_8261;
  wire [0:0] v_8262;
  wire [0:0] v_8263;
  wire [0:0] v_8264;
  wire [0:0] v_8265;
  function [0:0] mux_8265(input [0:0] sel);
    case (sel) 0: mux_8265 = 1'h0; 1: mux_8265 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8266;
  wire [0:0] v_8267;
  wire [0:0] v_8268;
  wire [0:0] v_8269;
  wire [0:0] v_8270;
  function [0:0] mux_8270(input [0:0] sel);
    case (sel) 0: mux_8270 = 1'h0; 1: mux_8270 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8271;
  wire [0:0] v_8272;
  wire [0:0] v_8273;
  wire [0:0] v_8274;
  function [0:0] mux_8274(input [0:0] sel);
    case (sel) 0: mux_8274 = 1'h0; 1: mux_8274 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8275;
  function [0:0] mux_8275(input [0:0] sel);
    case (sel) 0: mux_8275 = 1'h0; 1: mux_8275 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8276 = 1'h0;
  wire [0:0] v_8277;
  wire [0:0] v_8278;
  wire [0:0] act_8279;
  wire [0:0] v_8280;
  wire [0:0] v_8281;
  wire [0:0] v_8282;
  wire [0:0] vin0_consume_en_8283;
  wire [0:0] vout_canPeek_8283;
  wire [7:0] vout_peek_8283;
  wire [0:0] v_8284;
  wire [0:0] v_8285;
  function [0:0] mux_8285(input [0:0] sel);
    case (sel) 0: mux_8285 = 1'h0; 1: mux_8285 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8286;
  wire [0:0] v_8287;
  wire [0:0] v_8288;
  wire [0:0] v_8289;
  wire [0:0] v_8290;
  function [0:0] mux_8290(input [0:0] sel);
    case (sel) 0: mux_8290 = 1'h0; 1: mux_8290 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8291;
  wire [0:0] vin0_consume_en_8292;
  wire [0:0] vout_canPeek_8292;
  wire [7:0] vout_peek_8292;
  wire [0:0] v_8293;
  wire [0:0] v_8294;
  function [0:0] mux_8294(input [0:0] sel);
    case (sel) 0: mux_8294 = 1'h0; 1: mux_8294 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8295;
  function [0:0] mux_8295(input [0:0] sel);
    case (sel) 0: mux_8295 = 1'h0; 1: mux_8295 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8296;
  wire [0:0] v_8297;
  wire [0:0] v_8298;
  wire [0:0] v_8299;
  wire [0:0] v_8300;
  wire [0:0] v_8301;
  wire [0:0] v_8302;
  function [0:0] mux_8302(input [0:0] sel);
    case (sel) 0: mux_8302 = 1'h0; 1: mux_8302 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8303;
  function [0:0] mux_8303(input [0:0] sel);
    case (sel) 0: mux_8303 = 1'h0; 1: mux_8303 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8304;
  wire [0:0] v_8305;
  wire [0:0] v_8306;
  wire [0:0] v_8307;
  function [0:0] mux_8307(input [0:0] sel);
    case (sel) 0: mux_8307 = 1'h0; 1: mux_8307 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8308;
  function [0:0] mux_8308(input [0:0] sel);
    case (sel) 0: mux_8308 = 1'h0; 1: mux_8308 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8309;
  wire [0:0] v_8310;
  wire [0:0] v_8311;
  wire [0:0] v_8312;
  wire [0:0] v_8313;
  wire [0:0] v_8314;
  function [0:0] mux_8314(input [0:0] sel);
    case (sel) 0: mux_8314 = 1'h0; 1: mux_8314 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8315;
  wire [0:0] v_8316;
  wire [0:0] v_8317;
  wire [0:0] v_8318;
  wire [0:0] v_8319;
  function [0:0] mux_8319(input [0:0] sel);
    case (sel) 0: mux_8319 = 1'h0; 1: mux_8319 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8320;
  wire [0:0] v_8321;
  wire [0:0] v_8322;
  wire [0:0] v_8323;
  function [0:0] mux_8323(input [0:0] sel);
    case (sel) 0: mux_8323 = 1'h0; 1: mux_8323 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8324;
  function [0:0] mux_8324(input [0:0] sel);
    case (sel) 0: mux_8324 = 1'h0; 1: mux_8324 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8325 = 1'h0;
  wire [0:0] v_8326;
  wire [0:0] v_8327;
  wire [0:0] act_8328;
  wire [0:0] v_8329;
  wire [0:0] v_8330;
  wire [0:0] v_8331;
  reg [0:0] v_8332 = 1'h0;
  wire [0:0] v_8333;
  wire [0:0] v_8334;
  wire [0:0] act_8335;
  wire [0:0] v_8336;
  wire [0:0] v_8337;
  wire [0:0] v_8338;
  wire [0:0] vin0_consume_en_8339;
  wire [0:0] vout_canPeek_8339;
  wire [7:0] vout_peek_8339;
  wire [0:0] v_8340;
  wire [0:0] v_8341;
  function [0:0] mux_8341(input [0:0] sel);
    case (sel) 0: mux_8341 = 1'h0; 1: mux_8341 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8342;
  wire [0:0] v_8343;
  wire [0:0] v_8344;
  wire [0:0] v_8345;
  wire [0:0] v_8346;
  function [0:0] mux_8346(input [0:0] sel);
    case (sel) 0: mux_8346 = 1'h0; 1: mux_8346 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8347;
  wire [0:0] vin0_consume_en_8348;
  wire [0:0] vout_canPeek_8348;
  wire [7:0] vout_peek_8348;
  wire [0:0] v_8349;
  wire [0:0] v_8350;
  function [0:0] mux_8350(input [0:0] sel);
    case (sel) 0: mux_8350 = 1'h0; 1: mux_8350 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8351;
  function [0:0] mux_8351(input [0:0] sel);
    case (sel) 0: mux_8351 = 1'h0; 1: mux_8351 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8352;
  wire [0:0] v_8353;
  wire [0:0] v_8354;
  wire [0:0] v_8355;
  wire [0:0] v_8356;
  wire [0:0] v_8357;
  wire [0:0] v_8358;
  function [0:0] mux_8358(input [0:0] sel);
    case (sel) 0: mux_8358 = 1'h0; 1: mux_8358 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8359;
  wire [0:0] v_8360;
  wire [0:0] v_8361;
  wire [0:0] v_8362;
  wire [0:0] v_8363;
  function [0:0] mux_8363(input [0:0] sel);
    case (sel) 0: mux_8363 = 1'h0; 1: mux_8363 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8364;
  wire [0:0] v_8365;
  wire [0:0] v_8366;
  wire [0:0] v_8367;
  function [0:0] mux_8367(input [0:0] sel);
    case (sel) 0: mux_8367 = 1'h0; 1: mux_8367 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8368;
  function [0:0] mux_8368(input [0:0] sel);
    case (sel) 0: mux_8368 = 1'h0; 1: mux_8368 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8369 = 1'h0;
  wire [0:0] v_8370;
  wire [0:0] v_8371;
  wire [0:0] act_8372;
  wire [0:0] v_8373;
  wire [0:0] v_8374;
  wire [0:0] v_8375;
  wire [0:0] vin0_consume_en_8376;
  wire [0:0] vout_canPeek_8376;
  wire [7:0] vout_peek_8376;
  wire [0:0] v_8377;
  wire [0:0] v_8378;
  function [0:0] mux_8378(input [0:0] sel);
    case (sel) 0: mux_8378 = 1'h0; 1: mux_8378 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8379;
  wire [0:0] v_8380;
  wire [0:0] v_8381;
  wire [0:0] v_8382;
  wire [0:0] v_8383;
  function [0:0] mux_8383(input [0:0] sel);
    case (sel) 0: mux_8383 = 1'h0; 1: mux_8383 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8384;
  wire [0:0] vin0_consume_en_8385;
  wire [0:0] vout_canPeek_8385;
  wire [7:0] vout_peek_8385;
  wire [0:0] v_8386;
  wire [0:0] v_8387;
  function [0:0] mux_8387(input [0:0] sel);
    case (sel) 0: mux_8387 = 1'h0; 1: mux_8387 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8388;
  function [0:0] mux_8388(input [0:0] sel);
    case (sel) 0: mux_8388 = 1'h0; 1: mux_8388 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8389;
  wire [0:0] v_8390;
  wire [0:0] v_8391;
  wire [0:0] v_8392;
  wire [0:0] v_8393;
  wire [0:0] v_8394;
  wire [0:0] v_8395;
  function [0:0] mux_8395(input [0:0] sel);
    case (sel) 0: mux_8395 = 1'h0; 1: mux_8395 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8396;
  function [0:0] mux_8396(input [0:0] sel);
    case (sel) 0: mux_8396 = 1'h0; 1: mux_8396 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8397;
  wire [0:0] v_8398;
  wire [0:0] v_8399;
  wire [0:0] v_8400;
  function [0:0] mux_8400(input [0:0] sel);
    case (sel) 0: mux_8400 = 1'h0; 1: mux_8400 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8401;
  function [0:0] mux_8401(input [0:0] sel);
    case (sel) 0: mux_8401 = 1'h0; 1: mux_8401 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8402;
  wire [0:0] v_8403;
  wire [0:0] v_8404;
  wire [0:0] v_8405;
  wire [0:0] v_8406;
  wire [0:0] v_8407;
  function [0:0] mux_8407(input [0:0] sel);
    case (sel) 0: mux_8407 = 1'h0; 1: mux_8407 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8408;
  function [0:0] mux_8408(input [0:0] sel);
    case (sel) 0: mux_8408 = 1'h0; 1: mux_8408 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8409;
  wire [0:0] v_8410;
  wire [0:0] v_8411;
  wire [0:0] v_8412;
  function [0:0] mux_8412(input [0:0] sel);
    case (sel) 0: mux_8412 = 1'h0; 1: mux_8412 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8413;
  function [0:0] mux_8413(input [0:0] sel);
    case (sel) 0: mux_8413 = 1'h0; 1: mux_8413 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8414;
  wire [0:0] v_8415;
  wire [0:0] v_8416;
  wire [0:0] v_8417;
  wire [0:0] v_8418;
  wire [0:0] v_8419;
  function [0:0] mux_8419(input [0:0] sel);
    case (sel) 0: mux_8419 = 1'h0; 1: mux_8419 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8420;
  function [0:0] mux_8420(input [0:0] sel);
    case (sel) 0: mux_8420 = 1'h0; 1: mux_8420 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8421;
  wire [0:0] v_8422;
  wire [0:0] v_8423;
  wire [0:0] v_8424;
  function [0:0] mux_8424(input [0:0] sel);
    case (sel) 0: mux_8424 = 1'h0; 1: mux_8424 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8425;
  function [0:0] mux_8425(input [0:0] sel);
    case (sel) 0: mux_8425 = 1'h0; 1: mux_8425 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8426;
  wire [0:0] v_8427;
  wire [0:0] v_8428;
  wire [0:0] v_8429;
  wire [0:0] v_8430;
  wire [0:0] v_8431;
  function [0:0] mux_8431(input [0:0] sel);
    case (sel) 0: mux_8431 = 1'h0; 1: mux_8431 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8432;
  wire [0:0] v_8433;
  wire [0:0] v_8434;
  wire [0:0] v_8435;
  wire [0:0] v_8436;
  function [0:0] mux_8436(input [0:0] sel);
    case (sel) 0: mux_8436 = 1'h0; 1: mux_8436 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8437;
  wire [0:0] v_8438;
  wire [0:0] v_8439;
  wire [0:0] v_8440;
  function [0:0] mux_8440(input [0:0] sel);
    case (sel) 0: mux_8440 = 1'h0; 1: mux_8440 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8441;
  function [0:0] mux_8441(input [0:0] sel);
    case (sel) 0: mux_8441 = 1'h0; 1: mux_8441 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8442 = 1'h0;
  wire [0:0] v_8443;
  wire [0:0] v_8444;
  wire [0:0] act_8445;
  wire [0:0] v_8446;
  wire [0:0] v_8447;
  wire [0:0] v_8448;
  reg [0:0] v_8449 = 1'h0;
  wire [0:0] v_8450;
  wire [0:0] v_8451;
  wire [0:0] act_8452;
  wire [0:0] v_8453;
  wire [0:0] v_8454;
  wire [0:0] v_8455;
  reg [0:0] v_8456 = 1'h0;
  wire [0:0] v_8457;
  wire [0:0] v_8458;
  wire [0:0] act_8459;
  wire [0:0] v_8460;
  wire [0:0] v_8461;
  wire [0:0] v_8462;
  reg [0:0] v_8463 = 1'h0;
  wire [0:0] v_8464;
  wire [0:0] v_8465;
  wire [0:0] act_8466;
  wire [0:0] v_8467;
  wire [0:0] v_8468;
  wire [0:0] v_8469;
  wire [0:0] vin0_consume_en_8470;
  wire [0:0] vout_canPeek_8470;
  wire [7:0] vout_peek_8470;
  wire [0:0] v_8471;
  wire [0:0] v_8472;
  function [0:0] mux_8472(input [0:0] sel);
    case (sel) 0: mux_8472 = 1'h0; 1: mux_8472 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8473;
  wire [0:0] v_8474;
  wire [0:0] v_8475;
  wire [0:0] v_8476;
  wire [0:0] v_8477;
  function [0:0] mux_8477(input [0:0] sel);
    case (sel) 0: mux_8477 = 1'h0; 1: mux_8477 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8478;
  wire [0:0] vin0_consume_en_8479;
  wire [0:0] vout_canPeek_8479;
  wire [7:0] vout_peek_8479;
  wire [0:0] v_8480;
  wire [0:0] v_8481;
  function [0:0] mux_8481(input [0:0] sel);
    case (sel) 0: mux_8481 = 1'h0; 1: mux_8481 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8482;
  function [0:0] mux_8482(input [0:0] sel);
    case (sel) 0: mux_8482 = 1'h0; 1: mux_8482 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8483;
  wire [0:0] v_8484;
  wire [0:0] v_8485;
  wire [0:0] v_8486;
  wire [0:0] v_8487;
  wire [0:0] v_8488;
  wire [0:0] v_8489;
  function [0:0] mux_8489(input [0:0] sel);
    case (sel) 0: mux_8489 = 1'h0; 1: mux_8489 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8490;
  wire [0:0] v_8491;
  wire [0:0] v_8492;
  wire [0:0] v_8493;
  wire [0:0] v_8494;
  function [0:0] mux_8494(input [0:0] sel);
    case (sel) 0: mux_8494 = 1'h0; 1: mux_8494 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8495;
  wire [0:0] v_8496;
  wire [0:0] v_8497;
  wire [0:0] v_8498;
  function [0:0] mux_8498(input [0:0] sel);
    case (sel) 0: mux_8498 = 1'h0; 1: mux_8498 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8499;
  function [0:0] mux_8499(input [0:0] sel);
    case (sel) 0: mux_8499 = 1'h0; 1: mux_8499 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8500 = 1'h0;
  wire [0:0] v_8501;
  wire [0:0] v_8502;
  wire [0:0] act_8503;
  wire [0:0] v_8504;
  wire [0:0] v_8505;
  wire [0:0] v_8506;
  wire [0:0] vin0_consume_en_8507;
  wire [0:0] vout_canPeek_8507;
  wire [7:0] vout_peek_8507;
  wire [0:0] v_8508;
  wire [0:0] v_8509;
  function [0:0] mux_8509(input [0:0] sel);
    case (sel) 0: mux_8509 = 1'h0; 1: mux_8509 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8510;
  wire [0:0] v_8511;
  wire [0:0] v_8512;
  wire [0:0] v_8513;
  wire [0:0] v_8514;
  function [0:0] mux_8514(input [0:0] sel);
    case (sel) 0: mux_8514 = 1'h0; 1: mux_8514 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8515;
  wire [0:0] vin0_consume_en_8516;
  wire [0:0] vout_canPeek_8516;
  wire [7:0] vout_peek_8516;
  wire [0:0] v_8517;
  wire [0:0] v_8518;
  function [0:0] mux_8518(input [0:0] sel);
    case (sel) 0: mux_8518 = 1'h0; 1: mux_8518 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8519;
  function [0:0] mux_8519(input [0:0] sel);
    case (sel) 0: mux_8519 = 1'h0; 1: mux_8519 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8520;
  wire [0:0] v_8521;
  wire [0:0] v_8522;
  wire [0:0] v_8523;
  wire [0:0] v_8524;
  wire [0:0] v_8525;
  wire [0:0] v_8526;
  function [0:0] mux_8526(input [0:0] sel);
    case (sel) 0: mux_8526 = 1'h0; 1: mux_8526 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8527;
  function [0:0] mux_8527(input [0:0] sel);
    case (sel) 0: mux_8527 = 1'h0; 1: mux_8527 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8528;
  wire [0:0] v_8529;
  wire [0:0] v_8530;
  wire [0:0] v_8531;
  function [0:0] mux_8531(input [0:0] sel);
    case (sel) 0: mux_8531 = 1'h0; 1: mux_8531 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8532;
  function [0:0] mux_8532(input [0:0] sel);
    case (sel) 0: mux_8532 = 1'h0; 1: mux_8532 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8533;
  wire [0:0] v_8534;
  wire [0:0] v_8535;
  wire [0:0] v_8536;
  wire [0:0] v_8537;
  wire [0:0] v_8538;
  function [0:0] mux_8538(input [0:0] sel);
    case (sel) 0: mux_8538 = 1'h0; 1: mux_8538 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8539;
  wire [0:0] v_8540;
  wire [0:0] v_8541;
  wire [0:0] v_8542;
  wire [0:0] v_8543;
  function [0:0] mux_8543(input [0:0] sel);
    case (sel) 0: mux_8543 = 1'h0; 1: mux_8543 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8544;
  wire [0:0] v_8545;
  wire [0:0] v_8546;
  wire [0:0] v_8547;
  function [0:0] mux_8547(input [0:0] sel);
    case (sel) 0: mux_8547 = 1'h0; 1: mux_8547 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8548;
  function [0:0] mux_8548(input [0:0] sel);
    case (sel) 0: mux_8548 = 1'h0; 1: mux_8548 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8549 = 1'h0;
  wire [0:0] v_8550;
  wire [0:0] v_8551;
  wire [0:0] act_8552;
  wire [0:0] v_8553;
  wire [0:0] v_8554;
  wire [0:0] v_8555;
  reg [0:0] v_8556 = 1'h0;
  wire [0:0] v_8557;
  wire [0:0] v_8558;
  wire [0:0] act_8559;
  wire [0:0] v_8560;
  wire [0:0] v_8561;
  wire [0:0] v_8562;
  wire [0:0] vin0_consume_en_8563;
  wire [0:0] vout_canPeek_8563;
  wire [7:0] vout_peek_8563;
  wire [0:0] v_8564;
  wire [0:0] v_8565;
  function [0:0] mux_8565(input [0:0] sel);
    case (sel) 0: mux_8565 = 1'h0; 1: mux_8565 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8566;
  wire [0:0] v_8567;
  wire [0:0] v_8568;
  wire [0:0] v_8569;
  wire [0:0] v_8570;
  function [0:0] mux_8570(input [0:0] sel);
    case (sel) 0: mux_8570 = 1'h0; 1: mux_8570 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8571;
  wire [0:0] vin0_consume_en_8572;
  wire [0:0] vout_canPeek_8572;
  wire [7:0] vout_peek_8572;
  wire [0:0] v_8573;
  wire [0:0] v_8574;
  function [0:0] mux_8574(input [0:0] sel);
    case (sel) 0: mux_8574 = 1'h0; 1: mux_8574 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8575;
  function [0:0] mux_8575(input [0:0] sel);
    case (sel) 0: mux_8575 = 1'h0; 1: mux_8575 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8576;
  wire [0:0] v_8577;
  wire [0:0] v_8578;
  wire [0:0] v_8579;
  wire [0:0] v_8580;
  wire [0:0] v_8581;
  wire [0:0] v_8582;
  function [0:0] mux_8582(input [0:0] sel);
    case (sel) 0: mux_8582 = 1'h0; 1: mux_8582 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8583;
  wire [0:0] v_8584;
  wire [0:0] v_8585;
  wire [0:0] v_8586;
  wire [0:0] v_8587;
  function [0:0] mux_8587(input [0:0] sel);
    case (sel) 0: mux_8587 = 1'h0; 1: mux_8587 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8588;
  wire [0:0] v_8589;
  wire [0:0] v_8590;
  wire [0:0] v_8591;
  function [0:0] mux_8591(input [0:0] sel);
    case (sel) 0: mux_8591 = 1'h0; 1: mux_8591 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8592;
  function [0:0] mux_8592(input [0:0] sel);
    case (sel) 0: mux_8592 = 1'h0; 1: mux_8592 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8593 = 1'h0;
  wire [0:0] v_8594;
  wire [0:0] v_8595;
  wire [0:0] act_8596;
  wire [0:0] v_8597;
  wire [0:0] v_8598;
  wire [0:0] v_8599;
  wire [0:0] vin0_consume_en_8600;
  wire [0:0] vout_canPeek_8600;
  wire [7:0] vout_peek_8600;
  wire [0:0] v_8601;
  wire [0:0] v_8602;
  function [0:0] mux_8602(input [0:0] sel);
    case (sel) 0: mux_8602 = 1'h0; 1: mux_8602 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8603;
  wire [0:0] v_8604;
  wire [0:0] v_8605;
  wire [0:0] v_8606;
  wire [0:0] v_8607;
  function [0:0] mux_8607(input [0:0] sel);
    case (sel) 0: mux_8607 = 1'h0; 1: mux_8607 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8608;
  wire [0:0] vin0_consume_en_8609;
  wire [0:0] vout_canPeek_8609;
  wire [7:0] vout_peek_8609;
  wire [0:0] v_8610;
  wire [0:0] v_8611;
  function [0:0] mux_8611(input [0:0] sel);
    case (sel) 0: mux_8611 = 1'h0; 1: mux_8611 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8612;
  function [0:0] mux_8612(input [0:0] sel);
    case (sel) 0: mux_8612 = 1'h0; 1: mux_8612 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8613;
  wire [0:0] v_8614;
  wire [0:0] v_8615;
  wire [0:0] v_8616;
  wire [0:0] v_8617;
  wire [0:0] v_8618;
  wire [0:0] v_8619;
  function [0:0] mux_8619(input [0:0] sel);
    case (sel) 0: mux_8619 = 1'h0; 1: mux_8619 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8620;
  function [0:0] mux_8620(input [0:0] sel);
    case (sel) 0: mux_8620 = 1'h0; 1: mux_8620 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8621;
  wire [0:0] v_8622;
  wire [0:0] v_8623;
  wire [0:0] v_8624;
  function [0:0] mux_8624(input [0:0] sel);
    case (sel) 0: mux_8624 = 1'h0; 1: mux_8624 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8625;
  function [0:0] mux_8625(input [0:0] sel);
    case (sel) 0: mux_8625 = 1'h0; 1: mux_8625 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8626;
  wire [0:0] v_8627;
  wire [0:0] v_8628;
  wire [0:0] v_8629;
  wire [0:0] v_8630;
  wire [0:0] v_8631;
  function [0:0] mux_8631(input [0:0] sel);
    case (sel) 0: mux_8631 = 1'h0; 1: mux_8631 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8632;
  function [0:0] mux_8632(input [0:0] sel);
    case (sel) 0: mux_8632 = 1'h0; 1: mux_8632 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8633;
  wire [0:0] v_8634;
  wire [0:0] v_8635;
  wire [0:0] v_8636;
  function [0:0] mux_8636(input [0:0] sel);
    case (sel) 0: mux_8636 = 1'h0; 1: mux_8636 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8637;
  function [0:0] mux_8637(input [0:0] sel);
    case (sel) 0: mux_8637 = 1'h0; 1: mux_8637 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8638;
  wire [0:0] v_8639;
  wire [0:0] v_8640;
  wire [0:0] v_8641;
  wire [0:0] v_8642;
  wire [0:0] v_8643;
  function [0:0] mux_8643(input [0:0] sel);
    case (sel) 0: mux_8643 = 1'h0; 1: mux_8643 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8644;
  wire [0:0] v_8645;
  wire [0:0] v_8646;
  wire [0:0] v_8647;
  wire [0:0] v_8648;
  function [0:0] mux_8648(input [0:0] sel);
    case (sel) 0: mux_8648 = 1'h0; 1: mux_8648 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8649;
  wire [0:0] v_8650;
  wire [0:0] v_8651;
  wire [0:0] v_8652;
  function [0:0] mux_8652(input [0:0] sel);
    case (sel) 0: mux_8652 = 1'h0; 1: mux_8652 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8653;
  function [0:0] mux_8653(input [0:0] sel);
    case (sel) 0: mux_8653 = 1'h0; 1: mux_8653 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8654 = 1'h0;
  wire [0:0] v_8655;
  wire [0:0] v_8656;
  wire [0:0] act_8657;
  wire [0:0] v_8658;
  wire [0:0] v_8659;
  wire [0:0] v_8660;
  reg [0:0] v_8661 = 1'h0;
  wire [0:0] v_8662;
  wire [0:0] v_8663;
  wire [0:0] act_8664;
  wire [0:0] v_8665;
  wire [0:0] v_8666;
  wire [0:0] v_8667;
  reg [0:0] v_8668 = 1'h0;
  wire [0:0] v_8669;
  wire [0:0] v_8670;
  wire [0:0] act_8671;
  wire [0:0] v_8672;
  wire [0:0] v_8673;
  wire [0:0] v_8674;
  wire [0:0] vin0_consume_en_8675;
  wire [0:0] vout_canPeek_8675;
  wire [7:0] vout_peek_8675;
  wire [0:0] v_8676;
  wire [0:0] v_8677;
  function [0:0] mux_8677(input [0:0] sel);
    case (sel) 0: mux_8677 = 1'h0; 1: mux_8677 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8678;
  wire [0:0] v_8679;
  wire [0:0] v_8680;
  wire [0:0] v_8681;
  wire [0:0] v_8682;
  function [0:0] mux_8682(input [0:0] sel);
    case (sel) 0: mux_8682 = 1'h0; 1: mux_8682 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8683;
  wire [0:0] vin0_consume_en_8684;
  wire [0:0] vout_canPeek_8684;
  wire [7:0] vout_peek_8684;
  wire [0:0] v_8685;
  wire [0:0] v_8686;
  function [0:0] mux_8686(input [0:0] sel);
    case (sel) 0: mux_8686 = 1'h0; 1: mux_8686 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8687;
  function [0:0] mux_8687(input [0:0] sel);
    case (sel) 0: mux_8687 = 1'h0; 1: mux_8687 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8688;
  wire [0:0] v_8689;
  wire [0:0] v_8690;
  wire [0:0] v_8691;
  wire [0:0] v_8692;
  wire [0:0] v_8693;
  wire [0:0] v_8694;
  function [0:0] mux_8694(input [0:0] sel);
    case (sel) 0: mux_8694 = 1'h0; 1: mux_8694 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8695;
  wire [0:0] v_8696;
  wire [0:0] v_8697;
  wire [0:0] v_8698;
  wire [0:0] v_8699;
  function [0:0] mux_8699(input [0:0] sel);
    case (sel) 0: mux_8699 = 1'h0; 1: mux_8699 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8700;
  wire [0:0] v_8701;
  wire [0:0] v_8702;
  wire [0:0] v_8703;
  function [0:0] mux_8703(input [0:0] sel);
    case (sel) 0: mux_8703 = 1'h0; 1: mux_8703 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8704;
  function [0:0] mux_8704(input [0:0] sel);
    case (sel) 0: mux_8704 = 1'h0; 1: mux_8704 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8705 = 1'h0;
  wire [0:0] v_8706;
  wire [0:0] v_8707;
  wire [0:0] act_8708;
  wire [0:0] v_8709;
  wire [0:0] v_8710;
  wire [0:0] v_8711;
  wire [0:0] vin0_consume_en_8712;
  wire [0:0] vout_canPeek_8712;
  wire [7:0] vout_peek_8712;
  wire [0:0] v_8713;
  wire [0:0] v_8714;
  function [0:0] mux_8714(input [0:0] sel);
    case (sel) 0: mux_8714 = 1'h0; 1: mux_8714 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8715;
  wire [0:0] v_8716;
  wire [0:0] v_8717;
  wire [0:0] v_8718;
  wire [0:0] v_8719;
  function [0:0] mux_8719(input [0:0] sel);
    case (sel) 0: mux_8719 = 1'h0; 1: mux_8719 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8720;
  wire [0:0] vin0_consume_en_8721;
  wire [0:0] vout_canPeek_8721;
  wire [7:0] vout_peek_8721;
  wire [0:0] v_8722;
  wire [0:0] v_8723;
  function [0:0] mux_8723(input [0:0] sel);
    case (sel) 0: mux_8723 = 1'h0; 1: mux_8723 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8724;
  function [0:0] mux_8724(input [0:0] sel);
    case (sel) 0: mux_8724 = 1'h0; 1: mux_8724 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8725;
  wire [0:0] v_8726;
  wire [0:0] v_8727;
  wire [0:0] v_8728;
  wire [0:0] v_8729;
  wire [0:0] v_8730;
  wire [0:0] v_8731;
  function [0:0] mux_8731(input [0:0] sel);
    case (sel) 0: mux_8731 = 1'h0; 1: mux_8731 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8732;
  function [0:0] mux_8732(input [0:0] sel);
    case (sel) 0: mux_8732 = 1'h0; 1: mux_8732 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8733;
  wire [0:0] v_8734;
  wire [0:0] v_8735;
  wire [0:0] v_8736;
  function [0:0] mux_8736(input [0:0] sel);
    case (sel) 0: mux_8736 = 1'h0; 1: mux_8736 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8737;
  function [0:0] mux_8737(input [0:0] sel);
    case (sel) 0: mux_8737 = 1'h0; 1: mux_8737 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8738;
  wire [0:0] v_8739;
  wire [0:0] v_8740;
  wire [0:0] v_8741;
  wire [0:0] v_8742;
  wire [0:0] v_8743;
  function [0:0] mux_8743(input [0:0] sel);
    case (sel) 0: mux_8743 = 1'h0; 1: mux_8743 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8744;
  wire [0:0] v_8745;
  wire [0:0] v_8746;
  wire [0:0] v_8747;
  wire [0:0] v_8748;
  function [0:0] mux_8748(input [0:0] sel);
    case (sel) 0: mux_8748 = 1'h0; 1: mux_8748 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8749;
  wire [0:0] v_8750;
  wire [0:0] v_8751;
  wire [0:0] v_8752;
  function [0:0] mux_8752(input [0:0] sel);
    case (sel) 0: mux_8752 = 1'h0; 1: mux_8752 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8753;
  function [0:0] mux_8753(input [0:0] sel);
    case (sel) 0: mux_8753 = 1'h0; 1: mux_8753 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8754 = 1'h0;
  wire [0:0] v_8755;
  wire [0:0] v_8756;
  wire [0:0] act_8757;
  wire [0:0] v_8758;
  wire [0:0] v_8759;
  wire [0:0] v_8760;
  reg [0:0] v_8761 = 1'h0;
  wire [0:0] v_8762;
  wire [0:0] v_8763;
  wire [0:0] act_8764;
  wire [0:0] v_8765;
  wire [0:0] v_8766;
  wire [0:0] v_8767;
  wire [0:0] vin0_consume_en_8768;
  wire [0:0] vout_canPeek_8768;
  wire [7:0] vout_peek_8768;
  wire [0:0] v_8769;
  wire [0:0] v_8770;
  function [0:0] mux_8770(input [0:0] sel);
    case (sel) 0: mux_8770 = 1'h0; 1: mux_8770 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8771;
  wire [0:0] v_8772;
  wire [0:0] v_8773;
  wire [0:0] v_8774;
  wire [0:0] v_8775;
  function [0:0] mux_8775(input [0:0] sel);
    case (sel) 0: mux_8775 = 1'h0; 1: mux_8775 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8776;
  wire [0:0] vin0_consume_en_8777;
  wire [0:0] vout_canPeek_8777;
  wire [7:0] vout_peek_8777;
  wire [0:0] v_8778;
  wire [0:0] v_8779;
  function [0:0] mux_8779(input [0:0] sel);
    case (sel) 0: mux_8779 = 1'h0; 1: mux_8779 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8780;
  function [0:0] mux_8780(input [0:0] sel);
    case (sel) 0: mux_8780 = 1'h0; 1: mux_8780 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8781;
  wire [0:0] v_8782;
  wire [0:0] v_8783;
  wire [0:0] v_8784;
  wire [0:0] v_8785;
  wire [0:0] v_8786;
  wire [0:0] v_8787;
  function [0:0] mux_8787(input [0:0] sel);
    case (sel) 0: mux_8787 = 1'h0; 1: mux_8787 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8788;
  wire [0:0] v_8789;
  wire [0:0] v_8790;
  wire [0:0] v_8791;
  wire [0:0] v_8792;
  function [0:0] mux_8792(input [0:0] sel);
    case (sel) 0: mux_8792 = 1'h0; 1: mux_8792 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8793;
  wire [0:0] v_8794;
  wire [0:0] v_8795;
  wire [0:0] v_8796;
  function [0:0] mux_8796(input [0:0] sel);
    case (sel) 0: mux_8796 = 1'h0; 1: mux_8796 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8797;
  function [0:0] mux_8797(input [0:0] sel);
    case (sel) 0: mux_8797 = 1'h0; 1: mux_8797 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8798 = 1'h0;
  wire [0:0] v_8799;
  wire [0:0] v_8800;
  wire [0:0] act_8801;
  wire [0:0] v_8802;
  wire [0:0] v_8803;
  wire [0:0] v_8804;
  wire [0:0] vin0_consume_en_8805;
  wire [0:0] vout_canPeek_8805;
  wire [7:0] vout_peek_8805;
  wire [0:0] v_8806;
  wire [0:0] v_8807;
  function [0:0] mux_8807(input [0:0] sel);
    case (sel) 0: mux_8807 = 1'h0; 1: mux_8807 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8808;
  wire [0:0] v_8809;
  wire [0:0] v_8810;
  wire [0:0] v_8811;
  wire [0:0] v_8812;
  function [0:0] mux_8812(input [0:0] sel);
    case (sel) 0: mux_8812 = 1'h0; 1: mux_8812 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8813;
  wire [0:0] vin0_consume_en_8814;
  wire [0:0] vout_canPeek_8814;
  wire [7:0] vout_peek_8814;
  wire [0:0] v_8815;
  wire [0:0] v_8816;
  function [0:0] mux_8816(input [0:0] sel);
    case (sel) 0: mux_8816 = 1'h0; 1: mux_8816 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8817;
  function [0:0] mux_8817(input [0:0] sel);
    case (sel) 0: mux_8817 = 1'h0; 1: mux_8817 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8818;
  wire [0:0] v_8819;
  wire [0:0] v_8820;
  wire [0:0] v_8821;
  wire [0:0] v_8822;
  wire [0:0] v_8823;
  wire [0:0] v_8824;
  function [0:0] mux_8824(input [0:0] sel);
    case (sel) 0: mux_8824 = 1'h0; 1: mux_8824 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8825;
  function [0:0] mux_8825(input [0:0] sel);
    case (sel) 0: mux_8825 = 1'h0; 1: mux_8825 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8826;
  wire [0:0] v_8827;
  wire [0:0] v_8828;
  wire [0:0] v_8829;
  function [0:0] mux_8829(input [0:0] sel);
    case (sel) 0: mux_8829 = 1'h0; 1: mux_8829 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8830;
  function [0:0] mux_8830(input [0:0] sel);
    case (sel) 0: mux_8830 = 1'h0; 1: mux_8830 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8831;
  wire [0:0] v_8832;
  wire [0:0] v_8833;
  wire [0:0] v_8834;
  wire [0:0] v_8835;
  wire [0:0] v_8836;
  function [0:0] mux_8836(input [0:0] sel);
    case (sel) 0: mux_8836 = 1'h0; 1: mux_8836 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8837;
  function [0:0] mux_8837(input [0:0] sel);
    case (sel) 0: mux_8837 = 1'h0; 1: mux_8837 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8838;
  wire [0:0] v_8839;
  wire [0:0] v_8840;
  wire [0:0] v_8841;
  function [0:0] mux_8841(input [0:0] sel);
    case (sel) 0: mux_8841 = 1'h0; 1: mux_8841 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8842;
  function [0:0] mux_8842(input [0:0] sel);
    case (sel) 0: mux_8842 = 1'h0; 1: mux_8842 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8843;
  wire [0:0] v_8844;
  wire [0:0] v_8845;
  wire [0:0] v_8846;
  wire [0:0] v_8847;
  wire [0:0] v_8848;
  function [0:0] mux_8848(input [0:0] sel);
    case (sel) 0: mux_8848 = 1'h0; 1: mux_8848 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8849;
  function [0:0] mux_8849(input [0:0] sel);
    case (sel) 0: mux_8849 = 1'h0; 1: mux_8849 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8850;
  wire [0:0] v_8851;
  wire [0:0] v_8852;
  wire [0:0] v_8853;
  function [0:0] mux_8853(input [0:0] sel);
    case (sel) 0: mux_8853 = 1'h0; 1: mux_8853 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8854;
  function [0:0] mux_8854(input [0:0] sel);
    case (sel) 0: mux_8854 = 1'h0; 1: mux_8854 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8855;
  wire [0:0] v_8856;
  wire [0:0] v_8857;
  wire [0:0] v_8858;
  wire [0:0] v_8859;
  wire [0:0] v_8860;
  function [0:0] mux_8860(input [0:0] sel);
    case (sel) 0: mux_8860 = 1'h0; 1: mux_8860 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8861;
  function [0:0] mux_8861(input [0:0] sel);
    case (sel) 0: mux_8861 = 1'h0; 1: mux_8861 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8862;
  wire [0:0] v_8863;
  wire [0:0] v_8864;
  wire [0:0] v_8865;
  function [0:0] mux_8865(input [0:0] sel);
    case (sel) 0: mux_8865 = 1'h0; 1: mux_8865 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8866;
  function [0:0] mux_8866(input [0:0] sel);
    case (sel) 0: mux_8866 = 1'h0; 1: mux_8866 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8867;
  wire [0:0] v_8868;
  wire [0:0] v_8869;
  wire [0:0] v_8870;
  wire [0:0] v_8871;
  wire [0:0] v_8872;
  function [0:0] mux_8872(input [0:0] sel);
    case (sel) 0: mux_8872 = 1'h0; 1: mux_8872 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8873;
  wire [0:0] v_8874;
  wire [0:0] v_8875;
  wire [0:0] v_8876;
  wire [0:0] v_8877;
  function [0:0] mux_8877(input [0:0] sel);
    case (sel) 0: mux_8877 = 1'h0; 1: mux_8877 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8878;
  wire [0:0] v_8879;
  wire [0:0] v_8880;
  wire [0:0] v_8881;
  function [0:0] mux_8881(input [0:0] sel);
    case (sel) 0: mux_8881 = 1'h0; 1: mux_8881 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8882;
  function [0:0] mux_8882(input [0:0] sel);
    case (sel) 0: mux_8882 = 1'h0; 1: mux_8882 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8883 = 1'h0;
  wire [0:0] v_8884;
  wire [0:0] v_8885;
  wire [0:0] act_8886;
  wire [0:0] v_8887;
  wire [0:0] v_8888;
  wire [0:0] v_8889;
  reg [0:0] v_8890 = 1'h0;
  wire [0:0] v_8891;
  wire [0:0] v_8892;
  wire [0:0] act_8893;
  wire [0:0] v_8894;
  wire [0:0] v_8895;
  wire [0:0] v_8896;
  reg [0:0] v_8897 = 1'h0;
  wire [0:0] v_8898;
  wire [0:0] v_8899;
  wire [0:0] act_8900;
  wire [0:0] v_8901;
  wire [0:0] v_8902;
  wire [0:0] v_8903;
  reg [0:0] v_8904 = 1'h0;
  wire [0:0] v_8905;
  wire [0:0] v_8906;
  wire [0:0] act_8907;
  wire [0:0] v_8908;
  wire [0:0] v_8909;
  wire [0:0] v_8910;
  reg [0:0] v_8911 = 1'h0;
  wire [0:0] v_8912;
  wire [0:0] v_8913;
  wire [0:0] act_8914;
  wire [0:0] v_8915;
  wire [0:0] v_8916;
  wire [0:0] v_8917;
  wire [0:0] vin0_consume_en_8918;
  wire [0:0] vout_canPeek_8918;
  wire [7:0] vout_peek_8918;
  wire [0:0] v_8919;
  wire [0:0] v_8920;
  function [0:0] mux_8920(input [0:0] sel);
    case (sel) 0: mux_8920 = 1'h0; 1: mux_8920 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8921;
  wire [0:0] v_8922;
  wire [0:0] v_8923;
  wire [0:0] v_8924;
  wire [0:0] v_8925;
  function [0:0] mux_8925(input [0:0] sel);
    case (sel) 0: mux_8925 = 1'h0; 1: mux_8925 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8926;
  wire [0:0] vin0_consume_en_8927;
  wire [0:0] vout_canPeek_8927;
  wire [7:0] vout_peek_8927;
  wire [0:0] v_8928;
  wire [0:0] v_8929;
  function [0:0] mux_8929(input [0:0] sel);
    case (sel) 0: mux_8929 = 1'h0; 1: mux_8929 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8930;
  function [0:0] mux_8930(input [0:0] sel);
    case (sel) 0: mux_8930 = 1'h0; 1: mux_8930 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8931;
  wire [0:0] v_8932;
  wire [0:0] v_8933;
  wire [0:0] v_8934;
  wire [0:0] v_8935;
  wire [0:0] v_8936;
  wire [0:0] v_8937;
  function [0:0] mux_8937(input [0:0] sel);
    case (sel) 0: mux_8937 = 1'h0; 1: mux_8937 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8938;
  wire [0:0] v_8939;
  wire [0:0] v_8940;
  wire [0:0] v_8941;
  wire [0:0] v_8942;
  function [0:0] mux_8942(input [0:0] sel);
    case (sel) 0: mux_8942 = 1'h0; 1: mux_8942 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8943;
  wire [0:0] v_8944;
  wire [0:0] v_8945;
  wire [0:0] v_8946;
  function [0:0] mux_8946(input [0:0] sel);
    case (sel) 0: mux_8946 = 1'h0; 1: mux_8946 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8947;
  function [0:0] mux_8947(input [0:0] sel);
    case (sel) 0: mux_8947 = 1'h0; 1: mux_8947 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8948 = 1'h0;
  wire [0:0] v_8949;
  wire [0:0] v_8950;
  wire [0:0] act_8951;
  wire [0:0] v_8952;
  wire [0:0] v_8953;
  wire [0:0] v_8954;
  wire [0:0] vin0_consume_en_8955;
  wire [0:0] vout_canPeek_8955;
  wire [7:0] vout_peek_8955;
  wire [0:0] v_8956;
  wire [0:0] v_8957;
  function [0:0] mux_8957(input [0:0] sel);
    case (sel) 0: mux_8957 = 1'h0; 1: mux_8957 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8958;
  wire [0:0] v_8959;
  wire [0:0] v_8960;
  wire [0:0] v_8961;
  wire [0:0] v_8962;
  function [0:0] mux_8962(input [0:0] sel);
    case (sel) 0: mux_8962 = 1'h0; 1: mux_8962 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8963;
  wire [0:0] vin0_consume_en_8964;
  wire [0:0] vout_canPeek_8964;
  wire [7:0] vout_peek_8964;
  wire [0:0] v_8965;
  wire [0:0] v_8966;
  function [0:0] mux_8966(input [0:0] sel);
    case (sel) 0: mux_8966 = 1'h0; 1: mux_8966 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8967;
  function [0:0] mux_8967(input [0:0] sel);
    case (sel) 0: mux_8967 = 1'h0; 1: mux_8967 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8968;
  wire [0:0] v_8969;
  wire [0:0] v_8970;
  wire [0:0] v_8971;
  wire [0:0] v_8972;
  wire [0:0] v_8973;
  wire [0:0] v_8974;
  function [0:0] mux_8974(input [0:0] sel);
    case (sel) 0: mux_8974 = 1'h0; 1: mux_8974 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8975;
  function [0:0] mux_8975(input [0:0] sel);
    case (sel) 0: mux_8975 = 1'h0; 1: mux_8975 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8976;
  wire [0:0] v_8977;
  wire [0:0] v_8978;
  wire [0:0] v_8979;
  function [0:0] mux_8979(input [0:0] sel);
    case (sel) 0: mux_8979 = 1'h0; 1: mux_8979 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8980;
  function [0:0] mux_8980(input [0:0] sel);
    case (sel) 0: mux_8980 = 1'h0; 1: mux_8980 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8981;
  wire [0:0] v_8982;
  wire [0:0] v_8983;
  wire [0:0] v_8984;
  wire [0:0] v_8985;
  wire [0:0] v_8986;
  function [0:0] mux_8986(input [0:0] sel);
    case (sel) 0: mux_8986 = 1'h0; 1: mux_8986 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8987;
  wire [0:0] v_8988;
  wire [0:0] v_8989;
  wire [0:0] v_8990;
  wire [0:0] v_8991;
  function [0:0] mux_8991(input [0:0] sel);
    case (sel) 0: mux_8991 = 1'h0; 1: mux_8991 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8992;
  wire [0:0] v_8993;
  wire [0:0] v_8994;
  wire [0:0] v_8995;
  function [0:0] mux_8995(input [0:0] sel);
    case (sel) 0: mux_8995 = 1'h0; 1: mux_8995 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8996;
  function [0:0] mux_8996(input [0:0] sel);
    case (sel) 0: mux_8996 = 1'h0; 1: mux_8996 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8997 = 1'h0;
  wire [0:0] v_8998;
  wire [0:0] v_8999;
  wire [0:0] act_9000;
  wire [0:0] v_9001;
  wire [0:0] v_9002;
  wire [0:0] v_9003;
  reg [0:0] v_9004 = 1'h0;
  wire [0:0] v_9005;
  wire [0:0] v_9006;
  wire [0:0] act_9007;
  wire [0:0] v_9008;
  wire [0:0] v_9009;
  wire [0:0] v_9010;
  wire [0:0] vin0_consume_en_9011;
  wire [0:0] vout_canPeek_9011;
  wire [7:0] vout_peek_9011;
  wire [0:0] v_9012;
  wire [0:0] v_9013;
  function [0:0] mux_9013(input [0:0] sel);
    case (sel) 0: mux_9013 = 1'h0; 1: mux_9013 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9014;
  wire [0:0] v_9015;
  wire [0:0] v_9016;
  wire [0:0] v_9017;
  wire [0:0] v_9018;
  function [0:0] mux_9018(input [0:0] sel);
    case (sel) 0: mux_9018 = 1'h0; 1: mux_9018 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9019;
  wire [0:0] vin0_consume_en_9020;
  wire [0:0] vout_canPeek_9020;
  wire [7:0] vout_peek_9020;
  wire [0:0] v_9021;
  wire [0:0] v_9022;
  function [0:0] mux_9022(input [0:0] sel);
    case (sel) 0: mux_9022 = 1'h0; 1: mux_9022 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9023;
  function [0:0] mux_9023(input [0:0] sel);
    case (sel) 0: mux_9023 = 1'h0; 1: mux_9023 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9024;
  wire [0:0] v_9025;
  wire [0:0] v_9026;
  wire [0:0] v_9027;
  wire [0:0] v_9028;
  wire [0:0] v_9029;
  wire [0:0] v_9030;
  function [0:0] mux_9030(input [0:0] sel);
    case (sel) 0: mux_9030 = 1'h0; 1: mux_9030 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9031;
  wire [0:0] v_9032;
  wire [0:0] v_9033;
  wire [0:0] v_9034;
  wire [0:0] v_9035;
  function [0:0] mux_9035(input [0:0] sel);
    case (sel) 0: mux_9035 = 1'h0; 1: mux_9035 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9036;
  wire [0:0] v_9037;
  wire [0:0] v_9038;
  wire [0:0] v_9039;
  function [0:0] mux_9039(input [0:0] sel);
    case (sel) 0: mux_9039 = 1'h0; 1: mux_9039 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9040;
  function [0:0] mux_9040(input [0:0] sel);
    case (sel) 0: mux_9040 = 1'h0; 1: mux_9040 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9041 = 1'h0;
  wire [0:0] v_9042;
  wire [0:0] v_9043;
  wire [0:0] act_9044;
  wire [0:0] v_9045;
  wire [0:0] v_9046;
  wire [0:0] v_9047;
  wire [0:0] vin0_consume_en_9048;
  wire [0:0] vout_canPeek_9048;
  wire [7:0] vout_peek_9048;
  wire [0:0] v_9049;
  wire [0:0] v_9050;
  function [0:0] mux_9050(input [0:0] sel);
    case (sel) 0: mux_9050 = 1'h0; 1: mux_9050 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9051;
  wire [0:0] v_9052;
  wire [0:0] v_9053;
  wire [0:0] v_9054;
  wire [0:0] v_9055;
  function [0:0] mux_9055(input [0:0] sel);
    case (sel) 0: mux_9055 = 1'h0; 1: mux_9055 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9056;
  wire [0:0] vin0_consume_en_9057;
  wire [0:0] vout_canPeek_9057;
  wire [7:0] vout_peek_9057;
  wire [0:0] v_9058;
  wire [0:0] v_9059;
  function [0:0] mux_9059(input [0:0] sel);
    case (sel) 0: mux_9059 = 1'h0; 1: mux_9059 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9060;
  function [0:0] mux_9060(input [0:0] sel);
    case (sel) 0: mux_9060 = 1'h0; 1: mux_9060 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9061;
  wire [0:0] v_9062;
  wire [0:0] v_9063;
  wire [0:0] v_9064;
  wire [0:0] v_9065;
  wire [0:0] v_9066;
  wire [0:0] v_9067;
  function [0:0] mux_9067(input [0:0] sel);
    case (sel) 0: mux_9067 = 1'h0; 1: mux_9067 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9068;
  function [0:0] mux_9068(input [0:0] sel);
    case (sel) 0: mux_9068 = 1'h0; 1: mux_9068 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9069;
  wire [0:0] v_9070;
  wire [0:0] v_9071;
  wire [0:0] v_9072;
  function [0:0] mux_9072(input [0:0] sel);
    case (sel) 0: mux_9072 = 1'h0; 1: mux_9072 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9073;
  function [0:0] mux_9073(input [0:0] sel);
    case (sel) 0: mux_9073 = 1'h0; 1: mux_9073 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9074;
  wire [0:0] v_9075;
  wire [0:0] v_9076;
  wire [0:0] v_9077;
  wire [0:0] v_9078;
  wire [0:0] v_9079;
  function [0:0] mux_9079(input [0:0] sel);
    case (sel) 0: mux_9079 = 1'h0; 1: mux_9079 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9080;
  function [0:0] mux_9080(input [0:0] sel);
    case (sel) 0: mux_9080 = 1'h0; 1: mux_9080 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9081;
  wire [0:0] v_9082;
  wire [0:0] v_9083;
  wire [0:0] v_9084;
  function [0:0] mux_9084(input [0:0] sel);
    case (sel) 0: mux_9084 = 1'h0; 1: mux_9084 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9085;
  function [0:0] mux_9085(input [0:0] sel);
    case (sel) 0: mux_9085 = 1'h0; 1: mux_9085 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9086;
  wire [0:0] v_9087;
  wire [0:0] v_9088;
  wire [0:0] v_9089;
  wire [0:0] v_9090;
  wire [0:0] v_9091;
  function [0:0] mux_9091(input [0:0] sel);
    case (sel) 0: mux_9091 = 1'h0; 1: mux_9091 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9092;
  wire [0:0] v_9093;
  wire [0:0] v_9094;
  wire [0:0] v_9095;
  wire [0:0] v_9096;
  function [0:0] mux_9096(input [0:0] sel);
    case (sel) 0: mux_9096 = 1'h0; 1: mux_9096 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9097;
  wire [0:0] v_9098;
  wire [0:0] v_9099;
  wire [0:0] v_9100;
  function [0:0] mux_9100(input [0:0] sel);
    case (sel) 0: mux_9100 = 1'h0; 1: mux_9100 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9101;
  function [0:0] mux_9101(input [0:0] sel);
    case (sel) 0: mux_9101 = 1'h0; 1: mux_9101 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9102 = 1'h0;
  wire [0:0] v_9103;
  wire [0:0] v_9104;
  wire [0:0] act_9105;
  wire [0:0] v_9106;
  wire [0:0] v_9107;
  wire [0:0] v_9108;
  reg [0:0] v_9109 = 1'h0;
  wire [0:0] v_9110;
  wire [0:0] v_9111;
  wire [0:0] act_9112;
  wire [0:0] v_9113;
  wire [0:0] v_9114;
  wire [0:0] v_9115;
  reg [0:0] v_9116 = 1'h0;
  wire [0:0] v_9117;
  wire [0:0] v_9118;
  wire [0:0] act_9119;
  wire [0:0] v_9120;
  wire [0:0] v_9121;
  wire [0:0] v_9122;
  wire [0:0] vin0_consume_en_9123;
  wire [0:0] vout_canPeek_9123;
  wire [7:0] vout_peek_9123;
  wire [0:0] v_9124;
  wire [0:0] v_9125;
  function [0:0] mux_9125(input [0:0] sel);
    case (sel) 0: mux_9125 = 1'h0; 1: mux_9125 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9126;
  wire [0:0] v_9127;
  wire [0:0] v_9128;
  wire [0:0] v_9129;
  wire [0:0] v_9130;
  function [0:0] mux_9130(input [0:0] sel);
    case (sel) 0: mux_9130 = 1'h0; 1: mux_9130 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9131;
  wire [0:0] vin0_consume_en_9132;
  wire [0:0] vout_canPeek_9132;
  wire [7:0] vout_peek_9132;
  wire [0:0] v_9133;
  wire [0:0] v_9134;
  function [0:0] mux_9134(input [0:0] sel);
    case (sel) 0: mux_9134 = 1'h0; 1: mux_9134 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9135;
  function [0:0] mux_9135(input [0:0] sel);
    case (sel) 0: mux_9135 = 1'h0; 1: mux_9135 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9136;
  wire [0:0] v_9137;
  wire [0:0] v_9138;
  wire [0:0] v_9139;
  wire [0:0] v_9140;
  wire [0:0] v_9141;
  wire [0:0] v_9142;
  function [0:0] mux_9142(input [0:0] sel);
    case (sel) 0: mux_9142 = 1'h0; 1: mux_9142 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9143;
  wire [0:0] v_9144;
  wire [0:0] v_9145;
  wire [0:0] v_9146;
  wire [0:0] v_9147;
  function [0:0] mux_9147(input [0:0] sel);
    case (sel) 0: mux_9147 = 1'h0; 1: mux_9147 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9148;
  wire [0:0] v_9149;
  wire [0:0] v_9150;
  wire [0:0] v_9151;
  function [0:0] mux_9151(input [0:0] sel);
    case (sel) 0: mux_9151 = 1'h0; 1: mux_9151 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9152;
  function [0:0] mux_9152(input [0:0] sel);
    case (sel) 0: mux_9152 = 1'h0; 1: mux_9152 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9153 = 1'h0;
  wire [0:0] v_9154;
  wire [0:0] v_9155;
  wire [0:0] act_9156;
  wire [0:0] v_9157;
  wire [0:0] v_9158;
  wire [0:0] v_9159;
  wire [0:0] vin0_consume_en_9160;
  wire [0:0] vout_canPeek_9160;
  wire [7:0] vout_peek_9160;
  wire [0:0] v_9161;
  wire [0:0] v_9162;
  function [0:0] mux_9162(input [0:0] sel);
    case (sel) 0: mux_9162 = 1'h0; 1: mux_9162 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9163;
  wire [0:0] v_9164;
  wire [0:0] v_9165;
  wire [0:0] v_9166;
  wire [0:0] v_9167;
  function [0:0] mux_9167(input [0:0] sel);
    case (sel) 0: mux_9167 = 1'h0; 1: mux_9167 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9168;
  wire [0:0] vin0_consume_en_9169;
  wire [0:0] vout_canPeek_9169;
  wire [7:0] vout_peek_9169;
  wire [0:0] v_9170;
  wire [0:0] v_9171;
  function [0:0] mux_9171(input [0:0] sel);
    case (sel) 0: mux_9171 = 1'h0; 1: mux_9171 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9172;
  function [0:0] mux_9172(input [0:0] sel);
    case (sel) 0: mux_9172 = 1'h0; 1: mux_9172 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9173;
  wire [0:0] v_9174;
  wire [0:0] v_9175;
  wire [0:0] v_9176;
  wire [0:0] v_9177;
  wire [0:0] v_9178;
  wire [0:0] v_9179;
  function [0:0] mux_9179(input [0:0] sel);
    case (sel) 0: mux_9179 = 1'h0; 1: mux_9179 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9180;
  function [0:0] mux_9180(input [0:0] sel);
    case (sel) 0: mux_9180 = 1'h0; 1: mux_9180 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9181;
  wire [0:0] v_9182;
  wire [0:0] v_9183;
  wire [0:0] v_9184;
  function [0:0] mux_9184(input [0:0] sel);
    case (sel) 0: mux_9184 = 1'h0; 1: mux_9184 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9185;
  function [0:0] mux_9185(input [0:0] sel);
    case (sel) 0: mux_9185 = 1'h0; 1: mux_9185 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9186;
  wire [0:0] v_9187;
  wire [0:0] v_9188;
  wire [0:0] v_9189;
  wire [0:0] v_9190;
  wire [0:0] v_9191;
  function [0:0] mux_9191(input [0:0] sel);
    case (sel) 0: mux_9191 = 1'h0; 1: mux_9191 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9192;
  wire [0:0] v_9193;
  wire [0:0] v_9194;
  wire [0:0] v_9195;
  wire [0:0] v_9196;
  function [0:0] mux_9196(input [0:0] sel);
    case (sel) 0: mux_9196 = 1'h0; 1: mux_9196 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9197;
  wire [0:0] v_9198;
  wire [0:0] v_9199;
  wire [0:0] v_9200;
  function [0:0] mux_9200(input [0:0] sel);
    case (sel) 0: mux_9200 = 1'h0; 1: mux_9200 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9201;
  function [0:0] mux_9201(input [0:0] sel);
    case (sel) 0: mux_9201 = 1'h0; 1: mux_9201 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9202 = 1'h0;
  wire [0:0] v_9203;
  wire [0:0] v_9204;
  wire [0:0] act_9205;
  wire [0:0] v_9206;
  wire [0:0] v_9207;
  wire [0:0] v_9208;
  reg [0:0] v_9209 = 1'h0;
  wire [0:0] v_9210;
  wire [0:0] v_9211;
  wire [0:0] act_9212;
  wire [0:0] v_9213;
  wire [0:0] v_9214;
  wire [0:0] v_9215;
  wire [0:0] vin0_consume_en_9216;
  wire [0:0] vout_canPeek_9216;
  wire [7:0] vout_peek_9216;
  wire [0:0] v_9217;
  wire [0:0] v_9218;
  function [0:0] mux_9218(input [0:0] sel);
    case (sel) 0: mux_9218 = 1'h0; 1: mux_9218 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9219;
  wire [0:0] v_9220;
  wire [0:0] v_9221;
  wire [0:0] v_9222;
  wire [0:0] v_9223;
  function [0:0] mux_9223(input [0:0] sel);
    case (sel) 0: mux_9223 = 1'h0; 1: mux_9223 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9224;
  wire [0:0] vin0_consume_en_9225;
  wire [0:0] vout_canPeek_9225;
  wire [7:0] vout_peek_9225;
  wire [0:0] v_9226;
  wire [0:0] v_9227;
  function [0:0] mux_9227(input [0:0] sel);
    case (sel) 0: mux_9227 = 1'h0; 1: mux_9227 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9228;
  function [0:0] mux_9228(input [0:0] sel);
    case (sel) 0: mux_9228 = 1'h0; 1: mux_9228 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9229;
  wire [0:0] v_9230;
  wire [0:0] v_9231;
  wire [0:0] v_9232;
  wire [0:0] v_9233;
  wire [0:0] v_9234;
  wire [0:0] v_9235;
  function [0:0] mux_9235(input [0:0] sel);
    case (sel) 0: mux_9235 = 1'h0; 1: mux_9235 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9236;
  wire [0:0] v_9237;
  wire [0:0] v_9238;
  wire [0:0] v_9239;
  wire [0:0] v_9240;
  function [0:0] mux_9240(input [0:0] sel);
    case (sel) 0: mux_9240 = 1'h0; 1: mux_9240 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9241;
  wire [0:0] v_9242;
  wire [0:0] v_9243;
  wire [0:0] v_9244;
  function [0:0] mux_9244(input [0:0] sel);
    case (sel) 0: mux_9244 = 1'h0; 1: mux_9244 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9245;
  function [0:0] mux_9245(input [0:0] sel);
    case (sel) 0: mux_9245 = 1'h0; 1: mux_9245 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9246 = 1'h0;
  wire [0:0] v_9247;
  wire [0:0] v_9248;
  wire [0:0] act_9249;
  wire [0:0] v_9250;
  wire [0:0] v_9251;
  wire [0:0] v_9252;
  wire [0:0] vin0_consume_en_9253;
  wire [0:0] vout_canPeek_9253;
  wire [7:0] vout_peek_9253;
  wire [0:0] v_9254;
  wire [0:0] v_9255;
  function [0:0] mux_9255(input [0:0] sel);
    case (sel) 0: mux_9255 = 1'h0; 1: mux_9255 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9256;
  wire [0:0] v_9257;
  wire [0:0] v_9258;
  wire [0:0] v_9259;
  wire [0:0] v_9260;
  function [0:0] mux_9260(input [0:0] sel);
    case (sel) 0: mux_9260 = 1'h0; 1: mux_9260 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9261;
  wire [0:0] vin0_consume_en_9262;
  wire [0:0] vout_canPeek_9262;
  wire [7:0] vout_peek_9262;
  wire [0:0] v_9263;
  wire [0:0] v_9264;
  function [0:0] mux_9264(input [0:0] sel);
    case (sel) 0: mux_9264 = 1'h0; 1: mux_9264 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9265;
  function [0:0] mux_9265(input [0:0] sel);
    case (sel) 0: mux_9265 = 1'h0; 1: mux_9265 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9266;
  wire [0:0] v_9267;
  wire [0:0] v_9268;
  wire [0:0] v_9269;
  wire [0:0] v_9270;
  wire [0:0] v_9271;
  wire [0:0] v_9272;
  function [0:0] mux_9272(input [0:0] sel);
    case (sel) 0: mux_9272 = 1'h0; 1: mux_9272 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9273;
  function [0:0] mux_9273(input [0:0] sel);
    case (sel) 0: mux_9273 = 1'h0; 1: mux_9273 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9274;
  wire [0:0] v_9275;
  wire [0:0] v_9276;
  wire [0:0] v_9277;
  function [0:0] mux_9277(input [0:0] sel);
    case (sel) 0: mux_9277 = 1'h0; 1: mux_9277 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9278;
  function [0:0] mux_9278(input [0:0] sel);
    case (sel) 0: mux_9278 = 1'h0; 1: mux_9278 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9279;
  wire [0:0] v_9280;
  wire [0:0] v_9281;
  wire [0:0] v_9282;
  wire [0:0] v_9283;
  wire [0:0] v_9284;
  function [0:0] mux_9284(input [0:0] sel);
    case (sel) 0: mux_9284 = 1'h0; 1: mux_9284 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9285;
  function [0:0] mux_9285(input [0:0] sel);
    case (sel) 0: mux_9285 = 1'h0; 1: mux_9285 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9286;
  wire [0:0] v_9287;
  wire [0:0] v_9288;
  wire [0:0] v_9289;
  function [0:0] mux_9289(input [0:0] sel);
    case (sel) 0: mux_9289 = 1'h0; 1: mux_9289 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9290;
  function [0:0] mux_9290(input [0:0] sel);
    case (sel) 0: mux_9290 = 1'h0; 1: mux_9290 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9291;
  wire [0:0] v_9292;
  wire [0:0] v_9293;
  wire [0:0] v_9294;
  wire [0:0] v_9295;
  wire [0:0] v_9296;
  function [0:0] mux_9296(input [0:0] sel);
    case (sel) 0: mux_9296 = 1'h0; 1: mux_9296 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9297;
  function [0:0] mux_9297(input [0:0] sel);
    case (sel) 0: mux_9297 = 1'h0; 1: mux_9297 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9298;
  wire [0:0] v_9299;
  wire [0:0] v_9300;
  wire [0:0] v_9301;
  function [0:0] mux_9301(input [0:0] sel);
    case (sel) 0: mux_9301 = 1'h0; 1: mux_9301 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9302;
  function [0:0] mux_9302(input [0:0] sel);
    case (sel) 0: mux_9302 = 1'h0; 1: mux_9302 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9303;
  wire [0:0] v_9304;
  wire [0:0] v_9305;
  wire [0:0] v_9306;
  wire [0:0] v_9307;
  wire [0:0] v_9308;
  function [0:0] mux_9308(input [0:0] sel);
    case (sel) 0: mux_9308 = 1'h0; 1: mux_9308 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9309;
  wire [0:0] v_9310;
  wire [0:0] v_9311;
  wire [0:0] v_9312;
  wire [0:0] v_9313;
  function [0:0] mux_9313(input [0:0] sel);
    case (sel) 0: mux_9313 = 1'h0; 1: mux_9313 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9314;
  wire [0:0] v_9315;
  wire [0:0] v_9316;
  wire [0:0] v_9317;
  function [0:0] mux_9317(input [0:0] sel);
    case (sel) 0: mux_9317 = 1'h0; 1: mux_9317 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9318;
  function [0:0] mux_9318(input [0:0] sel);
    case (sel) 0: mux_9318 = 1'h0; 1: mux_9318 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9319 = 1'h0;
  wire [0:0] v_9320;
  wire [0:0] v_9321;
  wire [0:0] act_9322;
  wire [0:0] v_9323;
  wire [0:0] v_9324;
  wire [0:0] v_9325;
  reg [0:0] v_9326 = 1'h0;
  wire [0:0] v_9327;
  wire [0:0] v_9328;
  wire [0:0] act_9329;
  wire [0:0] v_9330;
  wire [0:0] v_9331;
  wire [0:0] v_9332;
  reg [0:0] v_9333 = 1'h0;
  wire [0:0] v_9334;
  wire [0:0] v_9335;
  wire [0:0] act_9336;
  wire [0:0] v_9337;
  wire [0:0] v_9338;
  wire [0:0] v_9339;
  reg [0:0] v_9340 = 1'h0;
  wire [0:0] v_9341;
  wire [0:0] v_9342;
  wire [0:0] act_9343;
  wire [0:0] v_9344;
  wire [0:0] v_9345;
  wire [0:0] v_9346;
  wire [0:0] vin0_consume_en_9347;
  wire [0:0] vout_canPeek_9347;
  wire [7:0] vout_peek_9347;
  wire [0:0] v_9348;
  wire [0:0] v_9349;
  function [0:0] mux_9349(input [0:0] sel);
    case (sel) 0: mux_9349 = 1'h0; 1: mux_9349 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9350;
  wire [0:0] v_9351;
  wire [0:0] v_9352;
  wire [0:0] v_9353;
  wire [0:0] v_9354;
  function [0:0] mux_9354(input [0:0] sel);
    case (sel) 0: mux_9354 = 1'h0; 1: mux_9354 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9355;
  wire [0:0] vin0_consume_en_9356;
  wire [0:0] vout_canPeek_9356;
  wire [7:0] vout_peek_9356;
  wire [0:0] v_9357;
  wire [0:0] v_9358;
  function [0:0] mux_9358(input [0:0] sel);
    case (sel) 0: mux_9358 = 1'h0; 1: mux_9358 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9359;
  function [0:0] mux_9359(input [0:0] sel);
    case (sel) 0: mux_9359 = 1'h0; 1: mux_9359 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9360;
  wire [0:0] v_9361;
  wire [0:0] v_9362;
  wire [0:0] v_9363;
  wire [0:0] v_9364;
  wire [0:0] v_9365;
  wire [0:0] v_9366;
  function [0:0] mux_9366(input [0:0] sel);
    case (sel) 0: mux_9366 = 1'h0; 1: mux_9366 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9367;
  wire [0:0] v_9368;
  wire [0:0] v_9369;
  wire [0:0] v_9370;
  wire [0:0] v_9371;
  function [0:0] mux_9371(input [0:0] sel);
    case (sel) 0: mux_9371 = 1'h0; 1: mux_9371 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9372;
  wire [0:0] v_9373;
  wire [0:0] v_9374;
  wire [0:0] v_9375;
  function [0:0] mux_9375(input [0:0] sel);
    case (sel) 0: mux_9375 = 1'h0; 1: mux_9375 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9376;
  function [0:0] mux_9376(input [0:0] sel);
    case (sel) 0: mux_9376 = 1'h0; 1: mux_9376 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9377 = 1'h0;
  wire [0:0] v_9378;
  wire [0:0] v_9379;
  wire [0:0] act_9380;
  wire [0:0] v_9381;
  wire [0:0] v_9382;
  wire [0:0] v_9383;
  wire [0:0] vin0_consume_en_9384;
  wire [0:0] vout_canPeek_9384;
  wire [7:0] vout_peek_9384;
  wire [0:0] v_9385;
  wire [0:0] v_9386;
  function [0:0] mux_9386(input [0:0] sel);
    case (sel) 0: mux_9386 = 1'h0; 1: mux_9386 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9387;
  wire [0:0] v_9388;
  wire [0:0] v_9389;
  wire [0:0] v_9390;
  wire [0:0] v_9391;
  function [0:0] mux_9391(input [0:0] sel);
    case (sel) 0: mux_9391 = 1'h0; 1: mux_9391 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9392;
  wire [0:0] vin0_consume_en_9393;
  wire [0:0] vout_canPeek_9393;
  wire [7:0] vout_peek_9393;
  wire [0:0] v_9394;
  wire [0:0] v_9395;
  function [0:0] mux_9395(input [0:0] sel);
    case (sel) 0: mux_9395 = 1'h0; 1: mux_9395 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9396;
  function [0:0] mux_9396(input [0:0] sel);
    case (sel) 0: mux_9396 = 1'h0; 1: mux_9396 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9397;
  wire [0:0] v_9398;
  wire [0:0] v_9399;
  wire [0:0] v_9400;
  wire [0:0] v_9401;
  wire [0:0] v_9402;
  wire [0:0] v_9403;
  function [0:0] mux_9403(input [0:0] sel);
    case (sel) 0: mux_9403 = 1'h0; 1: mux_9403 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9404;
  function [0:0] mux_9404(input [0:0] sel);
    case (sel) 0: mux_9404 = 1'h0; 1: mux_9404 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9405;
  wire [0:0] v_9406;
  wire [0:0] v_9407;
  wire [0:0] v_9408;
  function [0:0] mux_9408(input [0:0] sel);
    case (sel) 0: mux_9408 = 1'h0; 1: mux_9408 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9409;
  function [0:0] mux_9409(input [0:0] sel);
    case (sel) 0: mux_9409 = 1'h0; 1: mux_9409 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9410;
  wire [0:0] v_9411;
  wire [0:0] v_9412;
  wire [0:0] v_9413;
  wire [0:0] v_9414;
  wire [0:0] v_9415;
  function [0:0] mux_9415(input [0:0] sel);
    case (sel) 0: mux_9415 = 1'h0; 1: mux_9415 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9416;
  wire [0:0] v_9417;
  wire [0:0] v_9418;
  wire [0:0] v_9419;
  wire [0:0] v_9420;
  function [0:0] mux_9420(input [0:0] sel);
    case (sel) 0: mux_9420 = 1'h0; 1: mux_9420 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9421;
  wire [0:0] v_9422;
  wire [0:0] v_9423;
  wire [0:0] v_9424;
  function [0:0] mux_9424(input [0:0] sel);
    case (sel) 0: mux_9424 = 1'h0; 1: mux_9424 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9425;
  function [0:0] mux_9425(input [0:0] sel);
    case (sel) 0: mux_9425 = 1'h0; 1: mux_9425 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9426 = 1'h0;
  wire [0:0] v_9427;
  wire [0:0] v_9428;
  wire [0:0] act_9429;
  wire [0:0] v_9430;
  wire [0:0] v_9431;
  wire [0:0] v_9432;
  reg [0:0] v_9433 = 1'h0;
  wire [0:0] v_9434;
  wire [0:0] v_9435;
  wire [0:0] act_9436;
  wire [0:0] v_9437;
  wire [0:0] v_9438;
  wire [0:0] v_9439;
  wire [0:0] vin0_consume_en_9440;
  wire [0:0] vout_canPeek_9440;
  wire [7:0] vout_peek_9440;
  wire [0:0] v_9441;
  wire [0:0] v_9442;
  function [0:0] mux_9442(input [0:0] sel);
    case (sel) 0: mux_9442 = 1'h0; 1: mux_9442 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9443;
  wire [0:0] v_9444;
  wire [0:0] v_9445;
  wire [0:0] v_9446;
  wire [0:0] v_9447;
  function [0:0] mux_9447(input [0:0] sel);
    case (sel) 0: mux_9447 = 1'h0; 1: mux_9447 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9448;
  wire [0:0] vin0_consume_en_9449;
  wire [0:0] vout_canPeek_9449;
  wire [7:0] vout_peek_9449;
  wire [0:0] v_9450;
  wire [0:0] v_9451;
  function [0:0] mux_9451(input [0:0] sel);
    case (sel) 0: mux_9451 = 1'h0; 1: mux_9451 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9452;
  function [0:0] mux_9452(input [0:0] sel);
    case (sel) 0: mux_9452 = 1'h0; 1: mux_9452 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9453;
  wire [0:0] v_9454;
  wire [0:0] v_9455;
  wire [0:0] v_9456;
  wire [0:0] v_9457;
  wire [0:0] v_9458;
  wire [0:0] v_9459;
  function [0:0] mux_9459(input [0:0] sel);
    case (sel) 0: mux_9459 = 1'h0; 1: mux_9459 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9460;
  wire [0:0] v_9461;
  wire [0:0] v_9462;
  wire [0:0] v_9463;
  wire [0:0] v_9464;
  function [0:0] mux_9464(input [0:0] sel);
    case (sel) 0: mux_9464 = 1'h0; 1: mux_9464 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9465;
  wire [0:0] v_9466;
  wire [0:0] v_9467;
  wire [0:0] v_9468;
  function [0:0] mux_9468(input [0:0] sel);
    case (sel) 0: mux_9468 = 1'h0; 1: mux_9468 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9469;
  function [0:0] mux_9469(input [0:0] sel);
    case (sel) 0: mux_9469 = 1'h0; 1: mux_9469 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9470 = 1'h0;
  wire [0:0] v_9471;
  wire [0:0] v_9472;
  wire [0:0] act_9473;
  wire [0:0] v_9474;
  wire [0:0] v_9475;
  wire [0:0] v_9476;
  wire [0:0] vin0_consume_en_9477;
  wire [0:0] vout_canPeek_9477;
  wire [7:0] vout_peek_9477;
  wire [0:0] v_9478;
  wire [0:0] v_9479;
  function [0:0] mux_9479(input [0:0] sel);
    case (sel) 0: mux_9479 = 1'h0; 1: mux_9479 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9480;
  wire [0:0] v_9481;
  wire [0:0] v_9482;
  wire [0:0] v_9483;
  wire [0:0] v_9484;
  function [0:0] mux_9484(input [0:0] sel);
    case (sel) 0: mux_9484 = 1'h0; 1: mux_9484 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9485;
  wire [0:0] vin0_consume_en_9486;
  wire [0:0] vout_canPeek_9486;
  wire [7:0] vout_peek_9486;
  wire [0:0] v_9487;
  wire [0:0] v_9488;
  function [0:0] mux_9488(input [0:0] sel);
    case (sel) 0: mux_9488 = 1'h0; 1: mux_9488 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9489;
  function [0:0] mux_9489(input [0:0] sel);
    case (sel) 0: mux_9489 = 1'h0; 1: mux_9489 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9490;
  wire [0:0] v_9491;
  wire [0:0] v_9492;
  wire [0:0] v_9493;
  wire [0:0] v_9494;
  wire [0:0] v_9495;
  wire [0:0] v_9496;
  function [0:0] mux_9496(input [0:0] sel);
    case (sel) 0: mux_9496 = 1'h0; 1: mux_9496 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9497;
  function [0:0] mux_9497(input [0:0] sel);
    case (sel) 0: mux_9497 = 1'h0; 1: mux_9497 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9498;
  wire [0:0] v_9499;
  wire [0:0] v_9500;
  wire [0:0] v_9501;
  function [0:0] mux_9501(input [0:0] sel);
    case (sel) 0: mux_9501 = 1'h0; 1: mux_9501 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9502;
  function [0:0] mux_9502(input [0:0] sel);
    case (sel) 0: mux_9502 = 1'h0; 1: mux_9502 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9503;
  wire [0:0] v_9504;
  wire [0:0] v_9505;
  wire [0:0] v_9506;
  wire [0:0] v_9507;
  wire [0:0] v_9508;
  function [0:0] mux_9508(input [0:0] sel);
    case (sel) 0: mux_9508 = 1'h0; 1: mux_9508 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9509;
  function [0:0] mux_9509(input [0:0] sel);
    case (sel) 0: mux_9509 = 1'h0; 1: mux_9509 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9510;
  wire [0:0] v_9511;
  wire [0:0] v_9512;
  wire [0:0] v_9513;
  function [0:0] mux_9513(input [0:0] sel);
    case (sel) 0: mux_9513 = 1'h0; 1: mux_9513 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9514;
  function [0:0] mux_9514(input [0:0] sel);
    case (sel) 0: mux_9514 = 1'h0; 1: mux_9514 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9515;
  wire [0:0] v_9516;
  wire [0:0] v_9517;
  wire [0:0] v_9518;
  wire [0:0] v_9519;
  wire [0:0] v_9520;
  function [0:0] mux_9520(input [0:0] sel);
    case (sel) 0: mux_9520 = 1'h0; 1: mux_9520 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9521;
  wire [0:0] v_9522;
  wire [0:0] v_9523;
  wire [0:0] v_9524;
  wire [0:0] v_9525;
  function [0:0] mux_9525(input [0:0] sel);
    case (sel) 0: mux_9525 = 1'h0; 1: mux_9525 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9526;
  wire [0:0] v_9527;
  wire [0:0] v_9528;
  wire [0:0] v_9529;
  function [0:0] mux_9529(input [0:0] sel);
    case (sel) 0: mux_9529 = 1'h0; 1: mux_9529 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9530;
  function [0:0] mux_9530(input [0:0] sel);
    case (sel) 0: mux_9530 = 1'h0; 1: mux_9530 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9531 = 1'h0;
  wire [0:0] v_9532;
  wire [0:0] v_9533;
  wire [0:0] act_9534;
  wire [0:0] v_9535;
  wire [0:0] v_9536;
  wire [0:0] v_9537;
  reg [0:0] v_9538 = 1'h0;
  wire [0:0] v_9539;
  wire [0:0] v_9540;
  wire [0:0] act_9541;
  wire [0:0] v_9542;
  wire [0:0] v_9543;
  wire [0:0] v_9544;
  reg [0:0] v_9545 = 1'h0;
  wire [0:0] v_9546;
  wire [0:0] v_9547;
  wire [0:0] act_9548;
  wire [0:0] v_9549;
  wire [0:0] v_9550;
  wire [0:0] v_9551;
  wire [0:0] vin0_consume_en_9552;
  wire [0:0] vout_canPeek_9552;
  wire [7:0] vout_peek_9552;
  wire [0:0] v_9553;
  wire [0:0] v_9554;
  function [0:0] mux_9554(input [0:0] sel);
    case (sel) 0: mux_9554 = 1'h0; 1: mux_9554 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9555;
  wire [0:0] v_9556;
  wire [0:0] v_9557;
  wire [0:0] v_9558;
  wire [0:0] v_9559;
  function [0:0] mux_9559(input [0:0] sel);
    case (sel) 0: mux_9559 = 1'h0; 1: mux_9559 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9560;
  wire [0:0] vin0_consume_en_9561;
  wire [0:0] vout_canPeek_9561;
  wire [7:0] vout_peek_9561;
  wire [0:0] v_9562;
  wire [0:0] v_9563;
  function [0:0] mux_9563(input [0:0] sel);
    case (sel) 0: mux_9563 = 1'h0; 1: mux_9563 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9564;
  function [0:0] mux_9564(input [0:0] sel);
    case (sel) 0: mux_9564 = 1'h0; 1: mux_9564 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9565;
  wire [0:0] v_9566;
  wire [0:0] v_9567;
  wire [0:0] v_9568;
  wire [0:0] v_9569;
  wire [0:0] v_9570;
  wire [0:0] v_9571;
  function [0:0] mux_9571(input [0:0] sel);
    case (sel) 0: mux_9571 = 1'h0; 1: mux_9571 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9572;
  wire [0:0] v_9573;
  wire [0:0] v_9574;
  wire [0:0] v_9575;
  wire [0:0] v_9576;
  function [0:0] mux_9576(input [0:0] sel);
    case (sel) 0: mux_9576 = 1'h0; 1: mux_9576 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9577;
  wire [0:0] v_9578;
  wire [0:0] v_9579;
  wire [0:0] v_9580;
  function [0:0] mux_9580(input [0:0] sel);
    case (sel) 0: mux_9580 = 1'h0; 1: mux_9580 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9581;
  function [0:0] mux_9581(input [0:0] sel);
    case (sel) 0: mux_9581 = 1'h0; 1: mux_9581 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9582 = 1'h0;
  wire [0:0] v_9583;
  wire [0:0] v_9584;
  wire [0:0] act_9585;
  wire [0:0] v_9586;
  wire [0:0] v_9587;
  wire [0:0] v_9588;
  wire [0:0] vin0_consume_en_9589;
  wire [0:0] vout_canPeek_9589;
  wire [7:0] vout_peek_9589;
  wire [0:0] v_9590;
  wire [0:0] v_9591;
  function [0:0] mux_9591(input [0:0] sel);
    case (sel) 0: mux_9591 = 1'h0; 1: mux_9591 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9592;
  wire [0:0] v_9593;
  wire [0:0] v_9594;
  wire [0:0] v_9595;
  wire [0:0] v_9596;
  function [0:0] mux_9596(input [0:0] sel);
    case (sel) 0: mux_9596 = 1'h0; 1: mux_9596 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9597;
  wire [0:0] vin0_consume_en_9598;
  wire [0:0] vout_canPeek_9598;
  wire [7:0] vout_peek_9598;
  wire [0:0] v_9599;
  wire [0:0] v_9600;
  function [0:0] mux_9600(input [0:0] sel);
    case (sel) 0: mux_9600 = 1'h0; 1: mux_9600 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9601;
  function [0:0] mux_9601(input [0:0] sel);
    case (sel) 0: mux_9601 = 1'h0; 1: mux_9601 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9602;
  wire [0:0] v_9603;
  wire [0:0] v_9604;
  wire [0:0] v_9605;
  wire [0:0] v_9606;
  wire [0:0] v_9607;
  wire [0:0] v_9608;
  function [0:0] mux_9608(input [0:0] sel);
    case (sel) 0: mux_9608 = 1'h0; 1: mux_9608 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9609;
  function [0:0] mux_9609(input [0:0] sel);
    case (sel) 0: mux_9609 = 1'h0; 1: mux_9609 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9610;
  wire [0:0] v_9611;
  wire [0:0] v_9612;
  wire [0:0] v_9613;
  function [0:0] mux_9613(input [0:0] sel);
    case (sel) 0: mux_9613 = 1'h0; 1: mux_9613 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9614;
  function [0:0] mux_9614(input [0:0] sel);
    case (sel) 0: mux_9614 = 1'h0; 1: mux_9614 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9615;
  wire [0:0] v_9616;
  wire [0:0] v_9617;
  wire [0:0] v_9618;
  wire [0:0] v_9619;
  wire [0:0] v_9620;
  function [0:0] mux_9620(input [0:0] sel);
    case (sel) 0: mux_9620 = 1'h0; 1: mux_9620 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9621;
  wire [0:0] v_9622;
  wire [0:0] v_9623;
  wire [0:0] v_9624;
  wire [0:0] v_9625;
  function [0:0] mux_9625(input [0:0] sel);
    case (sel) 0: mux_9625 = 1'h0; 1: mux_9625 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9626;
  wire [0:0] v_9627;
  wire [0:0] v_9628;
  wire [0:0] v_9629;
  function [0:0] mux_9629(input [0:0] sel);
    case (sel) 0: mux_9629 = 1'h0; 1: mux_9629 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9630;
  function [0:0] mux_9630(input [0:0] sel);
    case (sel) 0: mux_9630 = 1'h0; 1: mux_9630 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9631 = 1'h0;
  wire [0:0] v_9632;
  wire [0:0] v_9633;
  wire [0:0] act_9634;
  wire [0:0] v_9635;
  wire [0:0] v_9636;
  wire [0:0] v_9637;
  reg [0:0] v_9638 = 1'h0;
  wire [0:0] v_9639;
  wire [0:0] v_9640;
  wire [0:0] act_9641;
  wire [0:0] v_9642;
  wire [0:0] v_9643;
  wire [0:0] v_9644;
  wire [0:0] vin0_consume_en_9645;
  wire [0:0] vout_canPeek_9645;
  wire [7:0] vout_peek_9645;
  wire [0:0] v_9646;
  wire [0:0] v_9647;
  function [0:0] mux_9647(input [0:0] sel);
    case (sel) 0: mux_9647 = 1'h0; 1: mux_9647 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9648;
  wire [0:0] v_9649;
  wire [0:0] v_9650;
  wire [0:0] v_9651;
  wire [0:0] v_9652;
  function [0:0] mux_9652(input [0:0] sel);
    case (sel) 0: mux_9652 = 1'h0; 1: mux_9652 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9653;
  wire [0:0] vin0_consume_en_9654;
  wire [0:0] vout_canPeek_9654;
  wire [7:0] vout_peek_9654;
  wire [0:0] v_9655;
  wire [0:0] v_9656;
  function [0:0] mux_9656(input [0:0] sel);
    case (sel) 0: mux_9656 = 1'h0; 1: mux_9656 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9657;
  function [0:0] mux_9657(input [0:0] sel);
    case (sel) 0: mux_9657 = 1'h0; 1: mux_9657 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9658;
  wire [0:0] v_9659;
  wire [0:0] v_9660;
  wire [0:0] v_9661;
  wire [0:0] v_9662;
  wire [0:0] v_9663;
  wire [0:0] v_9664;
  function [0:0] mux_9664(input [0:0] sel);
    case (sel) 0: mux_9664 = 1'h0; 1: mux_9664 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9665;
  wire [0:0] v_9666;
  wire [0:0] v_9667;
  wire [0:0] v_9668;
  wire [0:0] v_9669;
  function [0:0] mux_9669(input [0:0] sel);
    case (sel) 0: mux_9669 = 1'h0; 1: mux_9669 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9670;
  wire [0:0] v_9671;
  wire [0:0] v_9672;
  wire [0:0] v_9673;
  function [0:0] mux_9673(input [0:0] sel);
    case (sel) 0: mux_9673 = 1'h0; 1: mux_9673 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9674;
  function [0:0] mux_9674(input [0:0] sel);
    case (sel) 0: mux_9674 = 1'h0; 1: mux_9674 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9675 = 1'h0;
  wire [0:0] v_9676;
  wire [0:0] v_9677;
  wire [0:0] act_9678;
  wire [0:0] v_9679;
  wire [0:0] v_9680;
  wire [0:0] v_9681;
  wire [0:0] vin0_consume_en_9682;
  wire [0:0] vout_canPeek_9682;
  wire [7:0] vout_peek_9682;
  wire [0:0] v_9683;
  wire [0:0] v_9684;
  function [0:0] mux_9684(input [0:0] sel);
    case (sel) 0: mux_9684 = 1'h0; 1: mux_9684 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9685;
  wire [0:0] v_9686;
  wire [0:0] v_9687;
  wire [0:0] v_9688;
  wire [0:0] v_9689;
  function [0:0] mux_9689(input [0:0] sel);
    case (sel) 0: mux_9689 = 1'h0; 1: mux_9689 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9690;
  wire [0:0] vin0_consume_en_9691;
  wire [0:0] vout_canPeek_9691;
  wire [7:0] vout_peek_9691;
  wire [0:0] v_9692;
  wire [0:0] v_9693;
  function [0:0] mux_9693(input [0:0] sel);
    case (sel) 0: mux_9693 = 1'h0; 1: mux_9693 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9694;
  function [0:0] mux_9694(input [0:0] sel);
    case (sel) 0: mux_9694 = 1'h0; 1: mux_9694 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9695;
  wire [0:0] v_9696;
  wire [0:0] v_9697;
  wire [0:0] v_9698;
  wire [0:0] v_9699;
  wire [0:0] v_9700;
  wire [0:0] v_9701;
  function [0:0] mux_9701(input [0:0] sel);
    case (sel) 0: mux_9701 = 1'h0; 1: mux_9701 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9702;
  function [0:0] mux_9702(input [0:0] sel);
    case (sel) 0: mux_9702 = 1'h0; 1: mux_9702 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9703;
  wire [0:0] v_9704;
  wire [0:0] v_9705;
  wire [0:0] v_9706;
  function [0:0] mux_9706(input [0:0] sel);
    case (sel) 0: mux_9706 = 1'h0; 1: mux_9706 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9707;
  function [0:0] mux_9707(input [0:0] sel);
    case (sel) 0: mux_9707 = 1'h0; 1: mux_9707 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9708;
  wire [0:0] v_9709;
  wire [0:0] v_9710;
  wire [0:0] v_9711;
  wire [0:0] v_9712;
  wire [0:0] v_9713;
  function [0:0] mux_9713(input [0:0] sel);
    case (sel) 0: mux_9713 = 1'h0; 1: mux_9713 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9714;
  function [0:0] mux_9714(input [0:0] sel);
    case (sel) 0: mux_9714 = 1'h0; 1: mux_9714 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9715;
  wire [0:0] v_9716;
  wire [0:0] v_9717;
  wire [0:0] v_9718;
  function [0:0] mux_9718(input [0:0] sel);
    case (sel) 0: mux_9718 = 1'h0; 1: mux_9718 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9719;
  function [0:0] mux_9719(input [0:0] sel);
    case (sel) 0: mux_9719 = 1'h0; 1: mux_9719 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9720;
  wire [0:0] v_9721;
  wire [0:0] v_9722;
  wire [0:0] v_9723;
  wire [0:0] v_9724;
  wire [0:0] v_9725;
  function [0:0] mux_9725(input [0:0] sel);
    case (sel) 0: mux_9725 = 1'h0; 1: mux_9725 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9726;
  function [0:0] mux_9726(input [0:0] sel);
    case (sel) 0: mux_9726 = 1'h0; 1: mux_9726 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9727;
  wire [0:0] v_9728;
  wire [0:0] v_9729;
  wire [0:0] v_9730;
  function [0:0] mux_9730(input [0:0] sel);
    case (sel) 0: mux_9730 = 1'h0; 1: mux_9730 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9731;
  function [0:0] mux_9731(input [0:0] sel);
    case (sel) 0: mux_9731 = 1'h0; 1: mux_9731 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9732;
  wire [0:0] v_9733;
  wire [0:0] v_9734;
  wire [0:0] v_9735;
  wire [0:0] v_9736;
  wire [0:0] v_9737;
  function [0:0] mux_9737(input [0:0] sel);
    case (sel) 0: mux_9737 = 1'h0; 1: mux_9737 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9738;
  function [0:0] mux_9738(input [0:0] sel);
    case (sel) 0: mux_9738 = 1'h0; 1: mux_9738 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9739;
  wire [0:0] v_9740;
  wire [0:0] v_9741;
  wire [0:0] v_9742;
  function [0:0] mux_9742(input [0:0] sel);
    case (sel) 0: mux_9742 = 1'h0; 1: mux_9742 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9743;
  function [0:0] mux_9743(input [0:0] sel);
    case (sel) 0: mux_9743 = 1'h0; 1: mux_9743 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9744;
  wire [0:0] v_9745;
  wire [0:0] v_9746;
  wire [0:0] v_9747;
  wire [0:0] v_9748;
  wire [0:0] v_9749;
  function [0:0] mux_9749(input [0:0] sel);
    case (sel) 0: mux_9749 = 1'h0; 1: mux_9749 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9750;
  function [0:0] mux_9750(input [0:0] sel);
    case (sel) 0: mux_9750 = 1'h0; 1: mux_9750 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9751;
  wire [0:0] v_9752;
  wire [0:0] v_9753;
  wire [0:0] v_9754;
  function [0:0] mux_9754(input [0:0] sel);
    case (sel) 0: mux_9754 = 1'h0; 1: mux_9754 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9755;
  function [0:0] mux_9755(input [0:0] sel);
    case (sel) 0: mux_9755 = 1'h0; 1: mux_9755 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9756;
  wire [0:0] v_9757;
  wire [0:0] v_9758;
  wire [0:0] v_9759;
  wire [0:0] v_9760;
  wire [0:0] v_9761;
  function [0:0] mux_9761(input [0:0] sel);
    case (sel) 0: mux_9761 = 1'h0; 1: mux_9761 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9762;
  wire [0:0] v_9763;
  wire [0:0] v_9764;
  wire [0:0] v_9765;
  wire [0:0] v_9766;
  function [0:0] mux_9766(input [0:0] sel);
    case (sel) 0: mux_9766 = 1'h0; 1: mux_9766 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9767;
  wire [0:0] v_9768;
  wire [0:0] v_9769;
  wire [0:0] v_9770;
  function [0:0] mux_9770(input [0:0] sel);
    case (sel) 0: mux_9770 = 1'h0; 1: mux_9770 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9771;
  function [0:0] mux_9771(input [0:0] sel);
    case (sel) 0: mux_9771 = 1'h0; 1: mux_9771 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9772 = 1'h0;
  wire [0:0] v_9773;
  wire [0:0] v_9774;
  wire [0:0] act_9775;
  wire [0:0] v_9776;
  wire [0:0] v_9777;
  wire [0:0] v_9778;
  reg [0:0] v_9779 = 1'h0;
  wire [0:0] v_9780;
  wire [0:0] v_9781;
  wire [0:0] act_9782;
  wire [0:0] v_9783;
  wire [0:0] v_9784;
  wire [0:0] v_9785;
  reg [0:0] v_9786 = 1'h0;
  wire [0:0] v_9787;
  wire [0:0] v_9788;
  wire [0:0] act_9789;
  wire [0:0] v_9790;
  wire [0:0] v_9791;
  wire [0:0] v_9792;
  reg [0:0] v_9793 = 1'h0;
  wire [0:0] v_9794;
  wire [0:0] v_9795;
  wire [0:0] act_9796;
  wire [0:0] v_9797;
  wire [0:0] v_9798;
  wire [0:0] v_9799;
  reg [0:0] v_9800 = 1'h0;
  wire [0:0] v_9801;
  wire [0:0] v_9802;
  wire [0:0] act_9803;
  wire [0:0] v_9804;
  wire [0:0] v_9805;
  wire [0:0] v_9806;
  reg [0:0] v_9807 = 1'h0;
  wire [0:0] v_9808;
  wire [0:0] v_9809;
  wire [0:0] act_9810;
  wire [0:0] v_9811;
  wire [0:0] v_9812;
  wire [0:0] v_9813;
  wire [0:0] vin0_consume_en_9814;
  wire [0:0] vout_canPeek_9814;
  wire [7:0] vout_peek_9814;
  wire [0:0] v_9815;
  wire [0:0] v_9816;
  function [0:0] mux_9816(input [0:0] sel);
    case (sel) 0: mux_9816 = 1'h0; 1: mux_9816 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9817;
  wire [0:0] v_9818;
  wire [0:0] v_9819;
  wire [0:0] v_9820;
  wire [0:0] v_9821;
  function [0:0] mux_9821(input [0:0] sel);
    case (sel) 0: mux_9821 = 1'h0; 1: mux_9821 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9822;
  wire [0:0] vin0_consume_en_9823;
  wire [0:0] vout_canPeek_9823;
  wire [7:0] vout_peek_9823;
  wire [0:0] v_9824;
  wire [0:0] v_9825;
  function [0:0] mux_9825(input [0:0] sel);
    case (sel) 0: mux_9825 = 1'h0; 1: mux_9825 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9826;
  function [0:0] mux_9826(input [0:0] sel);
    case (sel) 0: mux_9826 = 1'h0; 1: mux_9826 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9827;
  wire [0:0] v_9828;
  wire [0:0] v_9829;
  wire [0:0] v_9830;
  wire [0:0] v_9831;
  wire [0:0] v_9832;
  wire [0:0] v_9833;
  function [0:0] mux_9833(input [0:0] sel);
    case (sel) 0: mux_9833 = 1'h0; 1: mux_9833 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9834;
  wire [0:0] v_9835;
  wire [0:0] v_9836;
  wire [0:0] v_9837;
  wire [0:0] v_9838;
  function [0:0] mux_9838(input [0:0] sel);
    case (sel) 0: mux_9838 = 1'h0; 1: mux_9838 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9839;
  wire [0:0] v_9840;
  wire [0:0] v_9841;
  wire [0:0] v_9842;
  function [0:0] mux_9842(input [0:0] sel);
    case (sel) 0: mux_9842 = 1'h0; 1: mux_9842 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9843;
  function [0:0] mux_9843(input [0:0] sel);
    case (sel) 0: mux_9843 = 1'h0; 1: mux_9843 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9844 = 1'h0;
  wire [0:0] v_9845;
  wire [0:0] v_9846;
  wire [0:0] act_9847;
  wire [0:0] v_9848;
  wire [0:0] v_9849;
  wire [0:0] v_9850;
  wire [0:0] vin0_consume_en_9851;
  wire [0:0] vout_canPeek_9851;
  wire [7:0] vout_peek_9851;
  wire [0:0] v_9852;
  wire [0:0] v_9853;
  function [0:0] mux_9853(input [0:0] sel);
    case (sel) 0: mux_9853 = 1'h0; 1: mux_9853 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9854;
  wire [0:0] v_9855;
  wire [0:0] v_9856;
  wire [0:0] v_9857;
  wire [0:0] v_9858;
  function [0:0] mux_9858(input [0:0] sel);
    case (sel) 0: mux_9858 = 1'h0; 1: mux_9858 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9859;
  wire [0:0] vin0_consume_en_9860;
  wire [0:0] vout_canPeek_9860;
  wire [7:0] vout_peek_9860;
  wire [0:0] v_9861;
  wire [0:0] v_9862;
  function [0:0] mux_9862(input [0:0] sel);
    case (sel) 0: mux_9862 = 1'h0; 1: mux_9862 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9863;
  function [0:0] mux_9863(input [0:0] sel);
    case (sel) 0: mux_9863 = 1'h0; 1: mux_9863 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9864;
  wire [0:0] v_9865;
  wire [0:0] v_9866;
  wire [0:0] v_9867;
  wire [0:0] v_9868;
  wire [0:0] v_9869;
  wire [0:0] v_9870;
  function [0:0] mux_9870(input [0:0] sel);
    case (sel) 0: mux_9870 = 1'h0; 1: mux_9870 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9871;
  function [0:0] mux_9871(input [0:0] sel);
    case (sel) 0: mux_9871 = 1'h0; 1: mux_9871 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9872;
  wire [0:0] v_9873;
  wire [0:0] v_9874;
  wire [0:0] v_9875;
  function [0:0] mux_9875(input [0:0] sel);
    case (sel) 0: mux_9875 = 1'h0; 1: mux_9875 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9876;
  function [0:0] mux_9876(input [0:0] sel);
    case (sel) 0: mux_9876 = 1'h0; 1: mux_9876 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9877;
  wire [0:0] v_9878;
  wire [0:0] v_9879;
  wire [0:0] v_9880;
  wire [0:0] v_9881;
  wire [0:0] v_9882;
  function [0:0] mux_9882(input [0:0] sel);
    case (sel) 0: mux_9882 = 1'h0; 1: mux_9882 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9883;
  wire [0:0] v_9884;
  wire [0:0] v_9885;
  wire [0:0] v_9886;
  wire [0:0] v_9887;
  function [0:0] mux_9887(input [0:0] sel);
    case (sel) 0: mux_9887 = 1'h0; 1: mux_9887 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9888;
  wire [0:0] v_9889;
  wire [0:0] v_9890;
  wire [0:0] v_9891;
  function [0:0] mux_9891(input [0:0] sel);
    case (sel) 0: mux_9891 = 1'h0; 1: mux_9891 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9892;
  function [0:0] mux_9892(input [0:0] sel);
    case (sel) 0: mux_9892 = 1'h0; 1: mux_9892 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9893 = 1'h0;
  wire [0:0] v_9894;
  wire [0:0] v_9895;
  wire [0:0] act_9896;
  wire [0:0] v_9897;
  wire [0:0] v_9898;
  wire [0:0] v_9899;
  reg [0:0] v_9900 = 1'h0;
  wire [0:0] v_9901;
  wire [0:0] v_9902;
  wire [0:0] act_9903;
  wire [0:0] v_9904;
  wire [0:0] v_9905;
  wire [0:0] v_9906;
  wire [0:0] vin0_consume_en_9907;
  wire [0:0] vout_canPeek_9907;
  wire [7:0] vout_peek_9907;
  wire [0:0] v_9908;
  wire [0:0] v_9909;
  function [0:0] mux_9909(input [0:0] sel);
    case (sel) 0: mux_9909 = 1'h0; 1: mux_9909 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9910;
  wire [0:0] v_9911;
  wire [0:0] v_9912;
  wire [0:0] v_9913;
  wire [0:0] v_9914;
  function [0:0] mux_9914(input [0:0] sel);
    case (sel) 0: mux_9914 = 1'h0; 1: mux_9914 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9915;
  wire [0:0] vin0_consume_en_9916;
  wire [0:0] vout_canPeek_9916;
  wire [7:0] vout_peek_9916;
  wire [0:0] v_9917;
  wire [0:0] v_9918;
  function [0:0] mux_9918(input [0:0] sel);
    case (sel) 0: mux_9918 = 1'h0; 1: mux_9918 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9919;
  function [0:0] mux_9919(input [0:0] sel);
    case (sel) 0: mux_9919 = 1'h0; 1: mux_9919 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9920;
  wire [0:0] v_9921;
  wire [0:0] v_9922;
  wire [0:0] v_9923;
  wire [0:0] v_9924;
  wire [0:0] v_9925;
  wire [0:0] v_9926;
  function [0:0] mux_9926(input [0:0] sel);
    case (sel) 0: mux_9926 = 1'h0; 1: mux_9926 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9927;
  wire [0:0] v_9928;
  wire [0:0] v_9929;
  wire [0:0] v_9930;
  wire [0:0] v_9931;
  function [0:0] mux_9931(input [0:0] sel);
    case (sel) 0: mux_9931 = 1'h0; 1: mux_9931 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9932;
  wire [0:0] v_9933;
  wire [0:0] v_9934;
  wire [0:0] v_9935;
  function [0:0] mux_9935(input [0:0] sel);
    case (sel) 0: mux_9935 = 1'h0; 1: mux_9935 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9936;
  function [0:0] mux_9936(input [0:0] sel);
    case (sel) 0: mux_9936 = 1'h0; 1: mux_9936 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9937 = 1'h0;
  wire [0:0] v_9938;
  wire [0:0] v_9939;
  wire [0:0] act_9940;
  wire [0:0] v_9941;
  wire [0:0] v_9942;
  wire [0:0] v_9943;
  wire [0:0] vin0_consume_en_9944;
  wire [0:0] vout_canPeek_9944;
  wire [7:0] vout_peek_9944;
  wire [0:0] v_9945;
  wire [0:0] v_9946;
  function [0:0] mux_9946(input [0:0] sel);
    case (sel) 0: mux_9946 = 1'h0; 1: mux_9946 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9947;
  wire [0:0] v_9948;
  wire [0:0] v_9949;
  wire [0:0] v_9950;
  wire [0:0] v_9951;
  function [0:0] mux_9951(input [0:0] sel);
    case (sel) 0: mux_9951 = 1'h0; 1: mux_9951 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9952;
  wire [0:0] vin0_consume_en_9953;
  wire [0:0] vout_canPeek_9953;
  wire [7:0] vout_peek_9953;
  wire [0:0] v_9954;
  wire [0:0] v_9955;
  function [0:0] mux_9955(input [0:0] sel);
    case (sel) 0: mux_9955 = 1'h0; 1: mux_9955 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9956;
  function [0:0] mux_9956(input [0:0] sel);
    case (sel) 0: mux_9956 = 1'h0; 1: mux_9956 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9957;
  wire [0:0] v_9958;
  wire [0:0] v_9959;
  wire [0:0] v_9960;
  wire [0:0] v_9961;
  wire [0:0] v_9962;
  wire [0:0] v_9963;
  function [0:0] mux_9963(input [0:0] sel);
    case (sel) 0: mux_9963 = 1'h0; 1: mux_9963 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9964;
  function [0:0] mux_9964(input [0:0] sel);
    case (sel) 0: mux_9964 = 1'h0; 1: mux_9964 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9965;
  wire [0:0] v_9966;
  wire [0:0] v_9967;
  wire [0:0] v_9968;
  function [0:0] mux_9968(input [0:0] sel);
    case (sel) 0: mux_9968 = 1'h0; 1: mux_9968 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9969;
  function [0:0] mux_9969(input [0:0] sel);
    case (sel) 0: mux_9969 = 1'h0; 1: mux_9969 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9970;
  wire [0:0] v_9971;
  wire [0:0] v_9972;
  wire [0:0] v_9973;
  wire [0:0] v_9974;
  wire [0:0] v_9975;
  function [0:0] mux_9975(input [0:0] sel);
    case (sel) 0: mux_9975 = 1'h0; 1: mux_9975 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9976;
  function [0:0] mux_9976(input [0:0] sel);
    case (sel) 0: mux_9976 = 1'h0; 1: mux_9976 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9977;
  wire [0:0] v_9978;
  wire [0:0] v_9979;
  wire [0:0] v_9980;
  function [0:0] mux_9980(input [0:0] sel);
    case (sel) 0: mux_9980 = 1'h0; 1: mux_9980 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9981;
  function [0:0] mux_9981(input [0:0] sel);
    case (sel) 0: mux_9981 = 1'h0; 1: mux_9981 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9982;
  wire [0:0] v_9983;
  wire [0:0] v_9984;
  wire [0:0] v_9985;
  wire [0:0] v_9986;
  wire [0:0] v_9987;
  function [0:0] mux_9987(input [0:0] sel);
    case (sel) 0: mux_9987 = 1'h0; 1: mux_9987 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9988;
  wire [0:0] v_9989;
  wire [0:0] v_9990;
  wire [0:0] v_9991;
  wire [0:0] v_9992;
  function [0:0] mux_9992(input [0:0] sel);
    case (sel) 0: mux_9992 = 1'h0; 1: mux_9992 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9993;
  wire [0:0] v_9994;
  wire [0:0] v_9995;
  wire [0:0] v_9996;
  function [0:0] mux_9996(input [0:0] sel);
    case (sel) 0: mux_9996 = 1'h0; 1: mux_9996 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9997;
  function [0:0] mux_9997(input [0:0] sel);
    case (sel) 0: mux_9997 = 1'h0; 1: mux_9997 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9998 = 1'h0;
  wire [0:0] v_9999;
  wire [0:0] v_10000;
  wire [0:0] act_10001;
  wire [0:0] v_10002;
  wire [0:0] v_10003;
  wire [0:0] v_10004;
  reg [0:0] v_10005 = 1'h0;
  wire [0:0] v_10006;
  wire [0:0] v_10007;
  wire [0:0] act_10008;
  wire [0:0] v_10009;
  wire [0:0] v_10010;
  wire [0:0] v_10011;
  reg [0:0] v_10012 = 1'h0;
  wire [0:0] v_10013;
  wire [0:0] v_10014;
  wire [0:0] act_10015;
  wire [0:0] v_10016;
  wire [0:0] v_10017;
  wire [0:0] v_10018;
  wire [0:0] vin0_consume_en_10019;
  wire [0:0] vout_canPeek_10019;
  wire [7:0] vout_peek_10019;
  wire [0:0] v_10020;
  wire [0:0] v_10021;
  function [0:0] mux_10021(input [0:0] sel);
    case (sel) 0: mux_10021 = 1'h0; 1: mux_10021 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10022;
  wire [0:0] v_10023;
  wire [0:0] v_10024;
  wire [0:0] v_10025;
  wire [0:0] v_10026;
  function [0:0] mux_10026(input [0:0] sel);
    case (sel) 0: mux_10026 = 1'h0; 1: mux_10026 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10027;
  wire [0:0] vin0_consume_en_10028;
  wire [0:0] vout_canPeek_10028;
  wire [7:0] vout_peek_10028;
  wire [0:0] v_10029;
  wire [0:0] v_10030;
  function [0:0] mux_10030(input [0:0] sel);
    case (sel) 0: mux_10030 = 1'h0; 1: mux_10030 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10031;
  function [0:0] mux_10031(input [0:0] sel);
    case (sel) 0: mux_10031 = 1'h0; 1: mux_10031 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10032;
  wire [0:0] v_10033;
  wire [0:0] v_10034;
  wire [0:0] v_10035;
  wire [0:0] v_10036;
  wire [0:0] v_10037;
  wire [0:0] v_10038;
  function [0:0] mux_10038(input [0:0] sel);
    case (sel) 0: mux_10038 = 1'h0; 1: mux_10038 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10039;
  wire [0:0] v_10040;
  wire [0:0] v_10041;
  wire [0:0] v_10042;
  wire [0:0] v_10043;
  function [0:0] mux_10043(input [0:0] sel);
    case (sel) 0: mux_10043 = 1'h0; 1: mux_10043 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10044;
  wire [0:0] v_10045;
  wire [0:0] v_10046;
  wire [0:0] v_10047;
  function [0:0] mux_10047(input [0:0] sel);
    case (sel) 0: mux_10047 = 1'h0; 1: mux_10047 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10048;
  function [0:0] mux_10048(input [0:0] sel);
    case (sel) 0: mux_10048 = 1'h0; 1: mux_10048 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_10049 = 1'h0;
  wire [0:0] v_10050;
  wire [0:0] v_10051;
  wire [0:0] act_10052;
  wire [0:0] v_10053;
  wire [0:0] v_10054;
  wire [0:0] v_10055;
  wire [0:0] vin0_consume_en_10056;
  wire [0:0] vout_canPeek_10056;
  wire [7:0] vout_peek_10056;
  wire [0:0] v_10057;
  wire [0:0] v_10058;
  function [0:0] mux_10058(input [0:0] sel);
    case (sel) 0: mux_10058 = 1'h0; 1: mux_10058 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10059;
  wire [0:0] v_10060;
  wire [0:0] v_10061;
  wire [0:0] v_10062;
  wire [0:0] v_10063;
  function [0:0] mux_10063(input [0:0] sel);
    case (sel) 0: mux_10063 = 1'h0; 1: mux_10063 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10064;
  wire [0:0] vin0_consume_en_10065;
  wire [0:0] vout_canPeek_10065;
  wire [7:0] vout_peek_10065;
  wire [0:0] v_10066;
  wire [0:0] v_10067;
  function [0:0] mux_10067(input [0:0] sel);
    case (sel) 0: mux_10067 = 1'h0; 1: mux_10067 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10068;
  function [0:0] mux_10068(input [0:0] sel);
    case (sel) 0: mux_10068 = 1'h0; 1: mux_10068 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10069;
  wire [0:0] v_10070;
  wire [0:0] v_10071;
  wire [0:0] v_10072;
  wire [0:0] v_10073;
  wire [0:0] v_10074;
  wire [0:0] v_10075;
  function [0:0] mux_10075(input [0:0] sel);
    case (sel) 0: mux_10075 = 1'h0; 1: mux_10075 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10076;
  function [0:0] mux_10076(input [0:0] sel);
    case (sel) 0: mux_10076 = 1'h0; 1: mux_10076 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10077;
  wire [0:0] v_10078;
  wire [0:0] v_10079;
  wire [0:0] v_10080;
  function [0:0] mux_10080(input [0:0] sel);
    case (sel) 0: mux_10080 = 1'h0; 1: mux_10080 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10081;
  function [0:0] mux_10081(input [0:0] sel);
    case (sel) 0: mux_10081 = 1'h0; 1: mux_10081 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10082;
  wire [0:0] v_10083;
  wire [0:0] v_10084;
  wire [0:0] v_10085;
  wire [0:0] v_10086;
  wire [0:0] v_10087;
  function [0:0] mux_10087(input [0:0] sel);
    case (sel) 0: mux_10087 = 1'h0; 1: mux_10087 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10088;
  wire [0:0] v_10089;
  wire [0:0] v_10090;
  wire [0:0] v_10091;
  wire [0:0] v_10092;
  function [0:0] mux_10092(input [0:0] sel);
    case (sel) 0: mux_10092 = 1'h0; 1: mux_10092 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10093;
  wire [0:0] v_10094;
  wire [0:0] v_10095;
  wire [0:0] v_10096;
  function [0:0] mux_10096(input [0:0] sel);
    case (sel) 0: mux_10096 = 1'h0; 1: mux_10096 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10097;
  function [0:0] mux_10097(input [0:0] sel);
    case (sel) 0: mux_10097 = 1'h0; 1: mux_10097 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_10098 = 1'h0;
  wire [0:0] v_10099;
  wire [0:0] v_10100;
  wire [0:0] act_10101;
  wire [0:0] v_10102;
  wire [0:0] v_10103;
  wire [0:0] v_10104;
  reg [0:0] v_10105 = 1'h0;
  wire [0:0] v_10106;
  wire [0:0] v_10107;
  wire [0:0] act_10108;
  wire [0:0] v_10109;
  wire [0:0] v_10110;
  wire [0:0] v_10111;
  wire [0:0] vin0_consume_en_10112;
  wire [0:0] vout_canPeek_10112;
  wire [7:0] vout_peek_10112;
  wire [0:0] v_10113;
  wire [0:0] v_10114;
  function [0:0] mux_10114(input [0:0] sel);
    case (sel) 0: mux_10114 = 1'h0; 1: mux_10114 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10115;
  wire [0:0] v_10116;
  wire [0:0] v_10117;
  wire [0:0] v_10118;
  wire [0:0] v_10119;
  function [0:0] mux_10119(input [0:0] sel);
    case (sel) 0: mux_10119 = 1'h0; 1: mux_10119 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10120;
  wire [0:0] vin0_consume_en_10121;
  wire [0:0] vout_canPeek_10121;
  wire [7:0] vout_peek_10121;
  wire [0:0] v_10122;
  wire [0:0] v_10123;
  function [0:0] mux_10123(input [0:0] sel);
    case (sel) 0: mux_10123 = 1'h0; 1: mux_10123 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10124;
  function [0:0] mux_10124(input [0:0] sel);
    case (sel) 0: mux_10124 = 1'h0; 1: mux_10124 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10125;
  wire [0:0] v_10126;
  wire [0:0] v_10127;
  wire [0:0] v_10128;
  wire [0:0] v_10129;
  wire [0:0] v_10130;
  wire [0:0] v_10131;
  function [0:0] mux_10131(input [0:0] sel);
    case (sel) 0: mux_10131 = 1'h0; 1: mux_10131 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10132;
  wire [0:0] v_10133;
  wire [0:0] v_10134;
  wire [0:0] v_10135;
  wire [0:0] v_10136;
  function [0:0] mux_10136(input [0:0] sel);
    case (sel) 0: mux_10136 = 1'h0; 1: mux_10136 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10137;
  wire [0:0] v_10138;
  wire [0:0] v_10139;
  wire [0:0] v_10140;
  function [0:0] mux_10140(input [0:0] sel);
    case (sel) 0: mux_10140 = 1'h0; 1: mux_10140 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10141;
  function [0:0] mux_10141(input [0:0] sel);
    case (sel) 0: mux_10141 = 1'h0; 1: mux_10141 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_10142 = 1'h0;
  wire [0:0] v_10143;
  wire [0:0] v_10144;
  wire [0:0] act_10145;
  wire [0:0] v_10146;
  wire [0:0] v_10147;
  wire [0:0] v_10148;
  wire [0:0] vin0_consume_en_10149;
  wire [0:0] vout_canPeek_10149;
  wire [7:0] vout_peek_10149;
  wire [0:0] v_10150;
  wire [0:0] v_10151;
  function [0:0] mux_10151(input [0:0] sel);
    case (sel) 0: mux_10151 = 1'h0; 1: mux_10151 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10152;
  wire [0:0] v_10153;
  wire [0:0] v_10154;
  wire [0:0] v_10155;
  wire [0:0] v_10156;
  function [0:0] mux_10156(input [0:0] sel);
    case (sel) 0: mux_10156 = 1'h0; 1: mux_10156 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10157;
  wire [0:0] vin0_consume_en_10158;
  wire [0:0] vout_canPeek_10158;
  wire [7:0] vout_peek_10158;
  wire [0:0] v_10159;
  wire [0:0] v_10160;
  function [0:0] mux_10160(input [0:0] sel);
    case (sel) 0: mux_10160 = 1'h0; 1: mux_10160 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10161;
  function [0:0] mux_10161(input [0:0] sel);
    case (sel) 0: mux_10161 = 1'h0; 1: mux_10161 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10162;
  wire [0:0] v_10163;
  wire [0:0] v_10164;
  wire [0:0] v_10165;
  wire [0:0] v_10166;
  wire [0:0] v_10167;
  wire [0:0] v_10168;
  function [0:0] mux_10168(input [0:0] sel);
    case (sel) 0: mux_10168 = 1'h0; 1: mux_10168 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10169;
  function [0:0] mux_10169(input [0:0] sel);
    case (sel) 0: mux_10169 = 1'h0; 1: mux_10169 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10170;
  wire [0:0] v_10171;
  wire [0:0] v_10172;
  wire [0:0] v_10173;
  function [0:0] mux_10173(input [0:0] sel);
    case (sel) 0: mux_10173 = 1'h0; 1: mux_10173 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10174;
  function [0:0] mux_10174(input [0:0] sel);
    case (sel) 0: mux_10174 = 1'h0; 1: mux_10174 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10175;
  wire [0:0] v_10176;
  wire [0:0] v_10177;
  wire [0:0] v_10178;
  wire [0:0] v_10179;
  wire [0:0] v_10180;
  function [0:0] mux_10180(input [0:0] sel);
    case (sel) 0: mux_10180 = 1'h0; 1: mux_10180 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10181;
  function [0:0] mux_10181(input [0:0] sel);
    case (sel) 0: mux_10181 = 1'h0; 1: mux_10181 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10182;
  wire [0:0] v_10183;
  wire [0:0] v_10184;
  wire [0:0] v_10185;
  function [0:0] mux_10185(input [0:0] sel);
    case (sel) 0: mux_10185 = 1'h0; 1: mux_10185 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10186;
  function [0:0] mux_10186(input [0:0] sel);
    case (sel) 0: mux_10186 = 1'h0; 1: mux_10186 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10187;
  wire [0:0] v_10188;
  wire [0:0] v_10189;
  wire [0:0] v_10190;
  wire [0:0] v_10191;
  wire [0:0] v_10192;
  function [0:0] mux_10192(input [0:0] sel);
    case (sel) 0: mux_10192 = 1'h0; 1: mux_10192 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10193;
  function [0:0] mux_10193(input [0:0] sel);
    case (sel) 0: mux_10193 = 1'h0; 1: mux_10193 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10194;
  wire [0:0] v_10195;
  wire [0:0] v_10196;
  wire [0:0] v_10197;
  function [0:0] mux_10197(input [0:0] sel);
    case (sel) 0: mux_10197 = 1'h0; 1: mux_10197 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10198;
  function [0:0] mux_10198(input [0:0] sel);
    case (sel) 0: mux_10198 = 1'h0; 1: mux_10198 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10199;
  wire [0:0] v_10200;
  wire [0:0] v_10201;
  wire [0:0] v_10202;
  wire [0:0] v_10203;
  wire [0:0] v_10204;
  function [0:0] mux_10204(input [0:0] sel);
    case (sel) 0: mux_10204 = 1'h0; 1: mux_10204 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10205;
  wire [0:0] v_10206;
  wire [0:0] v_10207;
  wire [0:0] v_10208;
  wire [0:0] v_10209;
  function [0:0] mux_10209(input [0:0] sel);
    case (sel) 0: mux_10209 = 1'h0; 1: mux_10209 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10210;
  wire [0:0] v_10211;
  wire [0:0] v_10212;
  wire [0:0] v_10213;
  function [0:0] mux_10213(input [0:0] sel);
    case (sel) 0: mux_10213 = 1'h0; 1: mux_10213 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10214;
  function [0:0] mux_10214(input [0:0] sel);
    case (sel) 0: mux_10214 = 1'h0; 1: mux_10214 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_10215 = 1'h0;
  wire [0:0] v_10216;
  wire [0:0] v_10217;
  wire [0:0] act_10218;
  wire [0:0] v_10219;
  wire [0:0] v_10220;
  wire [0:0] v_10221;
  reg [0:0] v_10222 = 1'h0;
  wire [0:0] v_10223;
  wire [0:0] v_10224;
  wire [0:0] act_10225;
  wire [0:0] v_10226;
  wire [0:0] v_10227;
  wire [0:0] v_10228;
  reg [0:0] v_10229 = 1'h0;
  wire [0:0] v_10230;
  wire [0:0] v_10231;
  wire [0:0] act_10232;
  wire [0:0] v_10233;
  wire [0:0] v_10234;
  wire [0:0] v_10235;
  reg [0:0] v_10236 = 1'h0;
  wire [0:0] v_10237;
  wire [0:0] v_10238;
  wire [0:0] act_10239;
  wire [0:0] v_10240;
  wire [0:0] v_10241;
  wire [0:0] v_10242;
  wire [0:0] vin0_consume_en_10243;
  wire [0:0] vout_canPeek_10243;
  wire [7:0] vout_peek_10243;
  wire [0:0] v_10244;
  wire [0:0] v_10245;
  function [0:0] mux_10245(input [0:0] sel);
    case (sel) 0: mux_10245 = 1'h0; 1: mux_10245 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10246;
  wire [0:0] v_10247;
  wire [0:0] v_10248;
  wire [0:0] v_10249;
  wire [0:0] v_10250;
  function [0:0] mux_10250(input [0:0] sel);
    case (sel) 0: mux_10250 = 1'h0; 1: mux_10250 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10251;
  wire [0:0] vin0_consume_en_10252;
  wire [0:0] vout_canPeek_10252;
  wire [7:0] vout_peek_10252;
  wire [0:0] v_10253;
  wire [0:0] v_10254;
  function [0:0] mux_10254(input [0:0] sel);
    case (sel) 0: mux_10254 = 1'h0; 1: mux_10254 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10255;
  function [0:0] mux_10255(input [0:0] sel);
    case (sel) 0: mux_10255 = 1'h0; 1: mux_10255 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10256;
  wire [0:0] v_10257;
  wire [0:0] v_10258;
  wire [0:0] v_10259;
  wire [0:0] v_10260;
  wire [0:0] v_10261;
  wire [0:0] v_10262;
  function [0:0] mux_10262(input [0:0] sel);
    case (sel) 0: mux_10262 = 1'h0; 1: mux_10262 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10263;
  wire [0:0] v_10264;
  wire [0:0] v_10265;
  wire [0:0] v_10266;
  wire [0:0] v_10267;
  function [0:0] mux_10267(input [0:0] sel);
    case (sel) 0: mux_10267 = 1'h0; 1: mux_10267 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10268;
  wire [0:0] v_10269;
  wire [0:0] v_10270;
  wire [0:0] v_10271;
  function [0:0] mux_10271(input [0:0] sel);
    case (sel) 0: mux_10271 = 1'h0; 1: mux_10271 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10272;
  function [0:0] mux_10272(input [0:0] sel);
    case (sel) 0: mux_10272 = 1'h0; 1: mux_10272 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_10273 = 1'h0;
  wire [0:0] v_10274;
  wire [0:0] v_10275;
  wire [0:0] act_10276;
  wire [0:0] v_10277;
  wire [0:0] v_10278;
  wire [0:0] v_10279;
  wire [0:0] vin0_consume_en_10280;
  wire [0:0] vout_canPeek_10280;
  wire [7:0] vout_peek_10280;
  wire [0:0] v_10281;
  wire [0:0] v_10282;
  function [0:0] mux_10282(input [0:0] sel);
    case (sel) 0: mux_10282 = 1'h0; 1: mux_10282 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10283;
  wire [0:0] v_10284;
  wire [0:0] v_10285;
  wire [0:0] v_10286;
  wire [0:0] v_10287;
  function [0:0] mux_10287(input [0:0] sel);
    case (sel) 0: mux_10287 = 1'h0; 1: mux_10287 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10288;
  wire [0:0] vin0_consume_en_10289;
  wire [0:0] vout_canPeek_10289;
  wire [7:0] vout_peek_10289;
  wire [0:0] v_10290;
  wire [0:0] v_10291;
  function [0:0] mux_10291(input [0:0] sel);
    case (sel) 0: mux_10291 = 1'h0; 1: mux_10291 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10292;
  function [0:0] mux_10292(input [0:0] sel);
    case (sel) 0: mux_10292 = 1'h0; 1: mux_10292 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10293;
  wire [0:0] v_10294;
  wire [0:0] v_10295;
  wire [0:0] v_10296;
  wire [0:0] v_10297;
  wire [0:0] v_10298;
  wire [0:0] v_10299;
  function [0:0] mux_10299(input [0:0] sel);
    case (sel) 0: mux_10299 = 1'h0; 1: mux_10299 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10300;
  function [0:0] mux_10300(input [0:0] sel);
    case (sel) 0: mux_10300 = 1'h0; 1: mux_10300 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10301;
  wire [0:0] v_10302;
  wire [0:0] v_10303;
  wire [0:0] v_10304;
  function [0:0] mux_10304(input [0:0] sel);
    case (sel) 0: mux_10304 = 1'h0; 1: mux_10304 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10305;
  function [0:0] mux_10305(input [0:0] sel);
    case (sel) 0: mux_10305 = 1'h0; 1: mux_10305 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10306;
  wire [0:0] v_10307;
  wire [0:0] v_10308;
  wire [0:0] v_10309;
  wire [0:0] v_10310;
  wire [0:0] v_10311;
  function [0:0] mux_10311(input [0:0] sel);
    case (sel) 0: mux_10311 = 1'h0; 1: mux_10311 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10312;
  wire [0:0] v_10313;
  wire [0:0] v_10314;
  wire [0:0] v_10315;
  wire [0:0] v_10316;
  function [0:0] mux_10316(input [0:0] sel);
    case (sel) 0: mux_10316 = 1'h0; 1: mux_10316 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10317;
  wire [0:0] v_10318;
  wire [0:0] v_10319;
  wire [0:0] v_10320;
  function [0:0] mux_10320(input [0:0] sel);
    case (sel) 0: mux_10320 = 1'h0; 1: mux_10320 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10321;
  function [0:0] mux_10321(input [0:0] sel);
    case (sel) 0: mux_10321 = 1'h0; 1: mux_10321 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_10322 = 1'h0;
  wire [0:0] v_10323;
  wire [0:0] v_10324;
  wire [0:0] act_10325;
  wire [0:0] v_10326;
  wire [0:0] v_10327;
  wire [0:0] v_10328;
  reg [0:0] v_10329 = 1'h0;
  wire [0:0] v_10330;
  wire [0:0] v_10331;
  wire [0:0] act_10332;
  wire [0:0] v_10333;
  wire [0:0] v_10334;
  wire [0:0] v_10335;
  wire [0:0] vin0_consume_en_10336;
  wire [0:0] vout_canPeek_10336;
  wire [7:0] vout_peek_10336;
  wire [0:0] v_10337;
  wire [0:0] v_10338;
  function [0:0] mux_10338(input [0:0] sel);
    case (sel) 0: mux_10338 = 1'h0; 1: mux_10338 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10339;
  wire [0:0] v_10340;
  wire [0:0] v_10341;
  wire [0:0] v_10342;
  wire [0:0] v_10343;
  function [0:0] mux_10343(input [0:0] sel);
    case (sel) 0: mux_10343 = 1'h0; 1: mux_10343 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10344;
  wire [0:0] vin0_consume_en_10345;
  wire [0:0] vout_canPeek_10345;
  wire [7:0] vout_peek_10345;
  wire [0:0] v_10346;
  wire [0:0] v_10347;
  function [0:0] mux_10347(input [0:0] sel);
    case (sel) 0: mux_10347 = 1'h0; 1: mux_10347 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10348;
  function [0:0] mux_10348(input [0:0] sel);
    case (sel) 0: mux_10348 = 1'h0; 1: mux_10348 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10349;
  wire [0:0] v_10350;
  wire [0:0] v_10351;
  wire [0:0] v_10352;
  wire [0:0] v_10353;
  wire [0:0] v_10354;
  wire [0:0] v_10355;
  function [0:0] mux_10355(input [0:0] sel);
    case (sel) 0: mux_10355 = 1'h0; 1: mux_10355 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10356;
  wire [0:0] v_10357;
  wire [0:0] v_10358;
  wire [0:0] v_10359;
  wire [0:0] v_10360;
  function [0:0] mux_10360(input [0:0] sel);
    case (sel) 0: mux_10360 = 1'h0; 1: mux_10360 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10361;
  wire [0:0] v_10362;
  wire [0:0] v_10363;
  wire [0:0] v_10364;
  function [0:0] mux_10364(input [0:0] sel);
    case (sel) 0: mux_10364 = 1'h0; 1: mux_10364 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10365;
  function [0:0] mux_10365(input [0:0] sel);
    case (sel) 0: mux_10365 = 1'h0; 1: mux_10365 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_10366 = 1'h0;
  wire [0:0] v_10367;
  wire [0:0] v_10368;
  wire [0:0] act_10369;
  wire [0:0] v_10370;
  wire [0:0] v_10371;
  wire [0:0] v_10372;
  wire [0:0] vin0_consume_en_10373;
  wire [0:0] vout_canPeek_10373;
  wire [7:0] vout_peek_10373;
  wire [0:0] v_10374;
  wire [0:0] v_10375;
  function [0:0] mux_10375(input [0:0] sel);
    case (sel) 0: mux_10375 = 1'h0; 1: mux_10375 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10376;
  wire [0:0] v_10377;
  wire [0:0] v_10378;
  wire [0:0] v_10379;
  wire [0:0] v_10380;
  function [0:0] mux_10380(input [0:0] sel);
    case (sel) 0: mux_10380 = 1'h0; 1: mux_10380 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10381;
  wire [0:0] vin0_consume_en_10382;
  wire [0:0] vout_canPeek_10382;
  wire [7:0] vout_peek_10382;
  wire [0:0] v_10383;
  wire [0:0] v_10384;
  function [0:0] mux_10384(input [0:0] sel);
    case (sel) 0: mux_10384 = 1'h0; 1: mux_10384 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10385;
  function [0:0] mux_10385(input [0:0] sel);
    case (sel) 0: mux_10385 = 1'h0; 1: mux_10385 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10386;
  wire [0:0] v_10387;
  wire [0:0] v_10388;
  wire [0:0] v_10389;
  wire [0:0] v_10390;
  wire [0:0] v_10391;
  wire [0:0] v_10392;
  function [0:0] mux_10392(input [0:0] sel);
    case (sel) 0: mux_10392 = 1'h0; 1: mux_10392 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10393;
  function [0:0] mux_10393(input [0:0] sel);
    case (sel) 0: mux_10393 = 1'h0; 1: mux_10393 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10394;
  wire [0:0] v_10395;
  wire [0:0] v_10396;
  wire [0:0] v_10397;
  function [0:0] mux_10397(input [0:0] sel);
    case (sel) 0: mux_10397 = 1'h0; 1: mux_10397 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10398;
  function [0:0] mux_10398(input [0:0] sel);
    case (sel) 0: mux_10398 = 1'h0; 1: mux_10398 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10399;
  wire [0:0] v_10400;
  wire [0:0] v_10401;
  wire [0:0] v_10402;
  wire [0:0] v_10403;
  wire [0:0] v_10404;
  function [0:0] mux_10404(input [0:0] sel);
    case (sel) 0: mux_10404 = 1'h0; 1: mux_10404 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10405;
  function [0:0] mux_10405(input [0:0] sel);
    case (sel) 0: mux_10405 = 1'h0; 1: mux_10405 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10406;
  wire [0:0] v_10407;
  wire [0:0] v_10408;
  wire [0:0] v_10409;
  function [0:0] mux_10409(input [0:0] sel);
    case (sel) 0: mux_10409 = 1'h0; 1: mux_10409 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10410;
  function [0:0] mux_10410(input [0:0] sel);
    case (sel) 0: mux_10410 = 1'h0; 1: mux_10410 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10411;
  wire [0:0] v_10412;
  wire [0:0] v_10413;
  wire [0:0] v_10414;
  wire [0:0] v_10415;
  wire [0:0] v_10416;
  function [0:0] mux_10416(input [0:0] sel);
    case (sel) 0: mux_10416 = 1'h0; 1: mux_10416 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10417;
  wire [0:0] v_10418;
  wire [0:0] v_10419;
  wire [0:0] v_10420;
  wire [0:0] v_10421;
  function [0:0] mux_10421(input [0:0] sel);
    case (sel) 0: mux_10421 = 1'h0; 1: mux_10421 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10422;
  wire [0:0] v_10423;
  wire [0:0] v_10424;
  wire [0:0] v_10425;
  function [0:0] mux_10425(input [0:0] sel);
    case (sel) 0: mux_10425 = 1'h0; 1: mux_10425 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10426;
  function [0:0] mux_10426(input [0:0] sel);
    case (sel) 0: mux_10426 = 1'h0; 1: mux_10426 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_10427 = 1'h0;
  wire [0:0] v_10428;
  wire [0:0] v_10429;
  wire [0:0] act_10430;
  wire [0:0] v_10431;
  wire [0:0] v_10432;
  wire [0:0] v_10433;
  reg [0:0] v_10434 = 1'h0;
  wire [0:0] v_10435;
  wire [0:0] v_10436;
  wire [0:0] act_10437;
  wire [0:0] v_10438;
  wire [0:0] v_10439;
  wire [0:0] v_10440;
  reg [0:0] v_10441 = 1'h0;
  wire [0:0] v_10442;
  wire [0:0] v_10443;
  wire [0:0] act_10444;
  wire [0:0] v_10445;
  wire [0:0] v_10446;
  wire [0:0] v_10447;
  wire [0:0] vin0_consume_en_10448;
  wire [0:0] vout_canPeek_10448;
  wire [7:0] vout_peek_10448;
  wire [0:0] v_10449;
  wire [0:0] v_10450;
  function [0:0] mux_10450(input [0:0] sel);
    case (sel) 0: mux_10450 = 1'h0; 1: mux_10450 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10451;
  wire [0:0] v_10452;
  wire [0:0] v_10453;
  wire [0:0] v_10454;
  wire [0:0] v_10455;
  function [0:0] mux_10455(input [0:0] sel);
    case (sel) 0: mux_10455 = 1'h0; 1: mux_10455 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10456;
  wire [0:0] vin0_consume_en_10457;
  wire [0:0] vout_canPeek_10457;
  wire [7:0] vout_peek_10457;
  wire [0:0] v_10458;
  wire [0:0] v_10459;
  function [0:0] mux_10459(input [0:0] sel);
    case (sel) 0: mux_10459 = 1'h0; 1: mux_10459 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10460;
  function [0:0] mux_10460(input [0:0] sel);
    case (sel) 0: mux_10460 = 1'h0; 1: mux_10460 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10461;
  wire [0:0] v_10462;
  wire [0:0] v_10463;
  wire [0:0] v_10464;
  wire [0:0] v_10465;
  wire [0:0] v_10466;
  wire [0:0] v_10467;
  function [0:0] mux_10467(input [0:0] sel);
    case (sel) 0: mux_10467 = 1'h0; 1: mux_10467 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10468;
  wire [0:0] v_10469;
  wire [0:0] v_10470;
  wire [0:0] v_10471;
  wire [0:0] v_10472;
  function [0:0] mux_10472(input [0:0] sel);
    case (sel) 0: mux_10472 = 1'h0; 1: mux_10472 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10473;
  wire [0:0] v_10474;
  wire [0:0] v_10475;
  wire [0:0] v_10476;
  function [0:0] mux_10476(input [0:0] sel);
    case (sel) 0: mux_10476 = 1'h0; 1: mux_10476 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10477;
  function [0:0] mux_10477(input [0:0] sel);
    case (sel) 0: mux_10477 = 1'h0; 1: mux_10477 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_10478 = 1'h0;
  wire [0:0] v_10479;
  wire [0:0] v_10480;
  wire [0:0] act_10481;
  wire [0:0] v_10482;
  wire [0:0] v_10483;
  wire [0:0] v_10484;
  wire [0:0] vin0_consume_en_10485;
  wire [0:0] vout_canPeek_10485;
  wire [7:0] vout_peek_10485;
  wire [0:0] v_10486;
  wire [0:0] v_10487;
  function [0:0] mux_10487(input [0:0] sel);
    case (sel) 0: mux_10487 = 1'h0; 1: mux_10487 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10488;
  wire [0:0] v_10489;
  wire [0:0] v_10490;
  wire [0:0] v_10491;
  wire [0:0] v_10492;
  function [0:0] mux_10492(input [0:0] sel);
    case (sel) 0: mux_10492 = 1'h0; 1: mux_10492 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10493;
  wire [0:0] vin0_consume_en_10494;
  wire [0:0] vout_canPeek_10494;
  wire [7:0] vout_peek_10494;
  wire [0:0] v_10495;
  wire [0:0] v_10496;
  function [0:0] mux_10496(input [0:0] sel);
    case (sel) 0: mux_10496 = 1'h0; 1: mux_10496 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10497;
  function [0:0] mux_10497(input [0:0] sel);
    case (sel) 0: mux_10497 = 1'h0; 1: mux_10497 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10498;
  wire [0:0] v_10499;
  wire [0:0] v_10500;
  wire [0:0] v_10501;
  wire [0:0] v_10502;
  wire [0:0] v_10503;
  wire [0:0] v_10504;
  function [0:0] mux_10504(input [0:0] sel);
    case (sel) 0: mux_10504 = 1'h0; 1: mux_10504 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10505;
  function [0:0] mux_10505(input [0:0] sel);
    case (sel) 0: mux_10505 = 1'h0; 1: mux_10505 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10506;
  wire [0:0] v_10507;
  wire [0:0] v_10508;
  wire [0:0] v_10509;
  function [0:0] mux_10509(input [0:0] sel);
    case (sel) 0: mux_10509 = 1'h0; 1: mux_10509 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10510;
  function [0:0] mux_10510(input [0:0] sel);
    case (sel) 0: mux_10510 = 1'h0; 1: mux_10510 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10511;
  wire [0:0] v_10512;
  wire [0:0] v_10513;
  wire [0:0] v_10514;
  wire [0:0] v_10515;
  wire [0:0] v_10516;
  function [0:0] mux_10516(input [0:0] sel);
    case (sel) 0: mux_10516 = 1'h0; 1: mux_10516 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10517;
  wire [0:0] v_10518;
  wire [0:0] v_10519;
  wire [0:0] v_10520;
  wire [0:0] v_10521;
  function [0:0] mux_10521(input [0:0] sel);
    case (sel) 0: mux_10521 = 1'h0; 1: mux_10521 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10522;
  wire [0:0] v_10523;
  wire [0:0] v_10524;
  wire [0:0] v_10525;
  function [0:0] mux_10525(input [0:0] sel);
    case (sel) 0: mux_10525 = 1'h0; 1: mux_10525 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10526;
  function [0:0] mux_10526(input [0:0] sel);
    case (sel) 0: mux_10526 = 1'h0; 1: mux_10526 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_10527 = 1'h0;
  wire [0:0] v_10528;
  wire [0:0] v_10529;
  wire [0:0] act_10530;
  wire [0:0] v_10531;
  wire [0:0] v_10532;
  wire [0:0] v_10533;
  reg [0:0] v_10534 = 1'h0;
  wire [0:0] v_10535;
  wire [0:0] v_10536;
  wire [0:0] act_10537;
  wire [0:0] v_10538;
  wire [0:0] v_10539;
  wire [0:0] v_10540;
  wire [0:0] vin0_consume_en_10541;
  wire [0:0] vout_canPeek_10541;
  wire [7:0] vout_peek_10541;
  wire [0:0] v_10542;
  wire [0:0] v_10543;
  function [0:0] mux_10543(input [0:0] sel);
    case (sel) 0: mux_10543 = 1'h0; 1: mux_10543 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10544;
  wire [0:0] v_10545;
  wire [0:0] v_10546;
  wire [0:0] v_10547;
  wire [0:0] v_10548;
  function [0:0] mux_10548(input [0:0] sel);
    case (sel) 0: mux_10548 = 1'h0; 1: mux_10548 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10549;
  wire [0:0] vin0_consume_en_10550;
  wire [0:0] vout_canPeek_10550;
  wire [7:0] vout_peek_10550;
  wire [0:0] v_10551;
  wire [0:0] v_10552;
  function [0:0] mux_10552(input [0:0] sel);
    case (sel) 0: mux_10552 = 1'h0; 1: mux_10552 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10553;
  function [0:0] mux_10553(input [0:0] sel);
    case (sel) 0: mux_10553 = 1'h0; 1: mux_10553 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10554;
  wire [0:0] v_10555;
  wire [0:0] v_10556;
  wire [0:0] v_10557;
  wire [0:0] v_10558;
  wire [0:0] v_10559;
  wire [0:0] v_10560;
  function [0:0] mux_10560(input [0:0] sel);
    case (sel) 0: mux_10560 = 1'h0; 1: mux_10560 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10561;
  wire [0:0] v_10562;
  wire [0:0] v_10563;
  wire [0:0] v_10564;
  wire [0:0] v_10565;
  function [0:0] mux_10565(input [0:0] sel);
    case (sel) 0: mux_10565 = 1'h0; 1: mux_10565 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10566;
  wire [0:0] v_10567;
  wire [0:0] v_10568;
  wire [0:0] v_10569;
  function [0:0] mux_10569(input [0:0] sel);
    case (sel) 0: mux_10569 = 1'h0; 1: mux_10569 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10570;
  function [0:0] mux_10570(input [0:0] sel);
    case (sel) 0: mux_10570 = 1'h0; 1: mux_10570 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_10571 = 1'h0;
  wire [0:0] v_10572;
  wire [0:0] v_10573;
  wire [0:0] act_10574;
  wire [0:0] v_10575;
  wire [0:0] v_10576;
  wire [0:0] v_10577;
  wire [0:0] vin0_consume_en_10578;
  wire [0:0] vout_canPeek_10578;
  wire [7:0] vout_peek_10578;
  wire [0:0] v_10579;
  wire [0:0] v_10580;
  function [0:0] mux_10580(input [0:0] sel);
    case (sel) 0: mux_10580 = 1'h0; 1: mux_10580 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10581;
  wire [0:0] v_10582;
  wire [0:0] v_10583;
  wire [0:0] v_10584;
  wire [0:0] v_10585;
  function [0:0] mux_10585(input [0:0] sel);
    case (sel) 0: mux_10585 = 1'h0; 1: mux_10585 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10586;
  wire [0:0] vin0_consume_en_10587;
  wire [0:0] vout_canPeek_10587;
  wire [7:0] vout_peek_10587;
  wire [0:0] v_10588;
  wire [0:0] v_10589;
  function [0:0] mux_10589(input [0:0] sel);
    case (sel) 0: mux_10589 = 1'h0; 1: mux_10589 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10590;
  function [0:0] mux_10590(input [0:0] sel);
    case (sel) 0: mux_10590 = 1'h0; 1: mux_10590 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10591;
  wire [0:0] v_10592;
  wire [0:0] v_10593;
  wire [0:0] v_10594;
  wire [0:0] v_10595;
  wire [0:0] v_10596;
  wire [0:0] v_10597;
  function [0:0] mux_10597(input [0:0] sel);
    case (sel) 0: mux_10597 = 1'h0; 1: mux_10597 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10598;
  function [0:0] mux_10598(input [0:0] sel);
    case (sel) 0: mux_10598 = 1'h0; 1: mux_10598 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10599;
  wire [0:0] v_10600;
  wire [0:0] v_10601;
  wire [0:0] v_10602;
  function [0:0] mux_10602(input [0:0] sel);
    case (sel) 0: mux_10602 = 1'h0; 1: mux_10602 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10603;
  function [0:0] mux_10603(input [0:0] sel);
    case (sel) 0: mux_10603 = 1'h0; 1: mux_10603 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10604;
  wire [0:0] v_10605;
  wire [0:0] v_10606;
  wire [0:0] v_10607;
  wire [0:0] v_10608;
  wire [0:0] v_10609;
  function [0:0] mux_10609(input [0:0] sel);
    case (sel) 0: mux_10609 = 1'h0; 1: mux_10609 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10610;
  function [0:0] mux_10610(input [0:0] sel);
    case (sel) 0: mux_10610 = 1'h0; 1: mux_10610 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10611;
  wire [0:0] v_10612;
  wire [0:0] v_10613;
  wire [0:0] v_10614;
  function [0:0] mux_10614(input [0:0] sel);
    case (sel) 0: mux_10614 = 1'h0; 1: mux_10614 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10615;
  function [0:0] mux_10615(input [0:0] sel);
    case (sel) 0: mux_10615 = 1'h0; 1: mux_10615 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10616;
  wire [0:0] v_10617;
  wire [0:0] v_10618;
  wire [0:0] v_10619;
  wire [0:0] v_10620;
  wire [0:0] v_10621;
  function [0:0] mux_10621(input [0:0] sel);
    case (sel) 0: mux_10621 = 1'h0; 1: mux_10621 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10622;
  function [0:0] mux_10622(input [0:0] sel);
    case (sel) 0: mux_10622 = 1'h0; 1: mux_10622 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10623;
  wire [0:0] v_10624;
  wire [0:0] v_10625;
  wire [0:0] v_10626;
  function [0:0] mux_10626(input [0:0] sel);
    case (sel) 0: mux_10626 = 1'h0; 1: mux_10626 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10627;
  function [0:0] mux_10627(input [0:0] sel);
    case (sel) 0: mux_10627 = 1'h0; 1: mux_10627 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10628;
  wire [0:0] v_10629;
  wire [0:0] v_10630;
  wire [0:0] v_10631;
  wire [0:0] v_10632;
  wire [0:0] v_10633;
  function [0:0] mux_10633(input [0:0] sel);
    case (sel) 0: mux_10633 = 1'h0; 1: mux_10633 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10634;
  function [0:0] mux_10634(input [0:0] sel);
    case (sel) 0: mux_10634 = 1'h0; 1: mux_10634 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10635;
  wire [0:0] v_10636;
  wire [0:0] v_10637;
  wire [0:0] v_10638;
  function [0:0] mux_10638(input [0:0] sel);
    case (sel) 0: mux_10638 = 1'h0; 1: mux_10638 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10639;
  function [0:0] mux_10639(input [0:0] sel);
    case (sel) 0: mux_10639 = 1'h0; 1: mux_10639 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10640;
  wire [0:0] v_10641;
  wire [0:0] v_10642;
  wire [0:0] v_10643;
  wire [0:0] v_10644;
  wire [0:0] v_10645;
  function [0:0] mux_10645(input [0:0] sel);
    case (sel) 0: mux_10645 = 1'h0; 1: mux_10645 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10646;
  wire [0:0] v_10647;
  wire [0:0] v_10648;
  wire [0:0] v_10649;
  wire [0:0] v_10650;
  function [0:0] mux_10650(input [0:0] sel);
    case (sel) 0: mux_10650 = 1'h0; 1: mux_10650 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10651;
  wire [0:0] v_10652;
  wire [0:0] v_10653;
  wire [0:0] v_10654;
  function [0:0] mux_10654(input [0:0] sel);
    case (sel) 0: mux_10654 = 1'h0; 1: mux_10654 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10655;
  function [0:0] mux_10655(input [0:0] sel);
    case (sel) 0: mux_10655 = 1'h0; 1: mux_10655 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_10656 = 1'h0;
  wire [0:0] v_10657;
  wire [0:0] v_10658;
  wire [0:0] act_10659;
  wire [0:0] v_10660;
  wire [0:0] v_10661;
  wire [0:0] v_10662;
  reg [0:0] v_10663 = 1'h0;
  wire [0:0] v_10664;
  wire [0:0] v_10665;
  wire [0:0] act_10666;
  wire [0:0] v_10667;
  wire [0:0] v_10668;
  wire [0:0] v_10669;
  reg [0:0] v_10670 = 1'h0;
  wire [0:0] v_10671;
  wire [0:0] v_10672;
  wire [0:0] act_10673;
  wire [0:0] v_10674;
  wire [0:0] v_10675;
  wire [0:0] v_10676;
  reg [0:0] v_10677 = 1'h0;
  wire [0:0] v_10678;
  wire [0:0] v_10679;
  wire [0:0] act_10680;
  wire [0:0] v_10681;
  wire [0:0] v_10682;
  wire [0:0] v_10683;
  reg [0:0] v_10684 = 1'h0;
  wire [0:0] v_10685;
  wire [0:0] v_10686;
  wire [0:0] act_10687;
  wire [0:0] v_10688;
  wire [0:0] v_10689;
  wire [0:0] v_10690;
  wire [0:0] vin0_consume_en_10691;
  wire [0:0] vout_canPeek_10691;
  wire [7:0] vout_peek_10691;
  wire [0:0] v_10692;
  wire [0:0] v_10693;
  function [0:0] mux_10693(input [0:0] sel);
    case (sel) 0: mux_10693 = 1'h0; 1: mux_10693 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10694;
  wire [0:0] v_10695;
  wire [0:0] v_10696;
  wire [0:0] v_10697;
  wire [0:0] v_10698;
  function [0:0] mux_10698(input [0:0] sel);
    case (sel) 0: mux_10698 = 1'h0; 1: mux_10698 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10699;
  wire [0:0] vin0_consume_en_10700;
  wire [0:0] vout_canPeek_10700;
  wire [7:0] vout_peek_10700;
  wire [0:0] v_10701;
  wire [0:0] v_10702;
  function [0:0] mux_10702(input [0:0] sel);
    case (sel) 0: mux_10702 = 1'h0; 1: mux_10702 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10703;
  function [0:0] mux_10703(input [0:0] sel);
    case (sel) 0: mux_10703 = 1'h0; 1: mux_10703 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10704;
  wire [0:0] v_10705;
  wire [0:0] v_10706;
  wire [0:0] v_10707;
  wire [0:0] v_10708;
  wire [0:0] v_10709;
  wire [0:0] v_10710;
  function [0:0] mux_10710(input [0:0] sel);
    case (sel) 0: mux_10710 = 1'h0; 1: mux_10710 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10711;
  wire [0:0] v_10712;
  wire [0:0] v_10713;
  wire [0:0] v_10714;
  wire [0:0] v_10715;
  function [0:0] mux_10715(input [0:0] sel);
    case (sel) 0: mux_10715 = 1'h0; 1: mux_10715 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10716;
  wire [0:0] v_10717;
  wire [0:0] v_10718;
  wire [0:0] v_10719;
  function [0:0] mux_10719(input [0:0] sel);
    case (sel) 0: mux_10719 = 1'h0; 1: mux_10719 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10720;
  function [0:0] mux_10720(input [0:0] sel);
    case (sel) 0: mux_10720 = 1'h0; 1: mux_10720 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_10721 = 1'h0;
  wire [0:0] v_10722;
  wire [0:0] v_10723;
  wire [0:0] act_10724;
  wire [0:0] v_10725;
  wire [0:0] v_10726;
  wire [0:0] v_10727;
  wire [0:0] vin0_consume_en_10728;
  wire [0:0] vout_canPeek_10728;
  wire [7:0] vout_peek_10728;
  wire [0:0] v_10729;
  wire [0:0] v_10730;
  function [0:0] mux_10730(input [0:0] sel);
    case (sel) 0: mux_10730 = 1'h0; 1: mux_10730 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10731;
  wire [0:0] v_10732;
  wire [0:0] v_10733;
  wire [0:0] v_10734;
  wire [0:0] v_10735;
  function [0:0] mux_10735(input [0:0] sel);
    case (sel) 0: mux_10735 = 1'h0; 1: mux_10735 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10736;
  wire [0:0] vin0_consume_en_10737;
  wire [0:0] vout_canPeek_10737;
  wire [7:0] vout_peek_10737;
  wire [0:0] v_10738;
  wire [0:0] v_10739;
  function [0:0] mux_10739(input [0:0] sel);
    case (sel) 0: mux_10739 = 1'h0; 1: mux_10739 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10740;
  function [0:0] mux_10740(input [0:0] sel);
    case (sel) 0: mux_10740 = 1'h0; 1: mux_10740 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10741;
  wire [0:0] v_10742;
  wire [0:0] v_10743;
  wire [0:0] v_10744;
  wire [0:0] v_10745;
  wire [0:0] v_10746;
  wire [0:0] v_10747;
  function [0:0] mux_10747(input [0:0] sel);
    case (sel) 0: mux_10747 = 1'h0; 1: mux_10747 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10748;
  function [0:0] mux_10748(input [0:0] sel);
    case (sel) 0: mux_10748 = 1'h0; 1: mux_10748 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10749;
  wire [0:0] v_10750;
  wire [0:0] v_10751;
  wire [0:0] v_10752;
  function [0:0] mux_10752(input [0:0] sel);
    case (sel) 0: mux_10752 = 1'h0; 1: mux_10752 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10753;
  function [0:0] mux_10753(input [0:0] sel);
    case (sel) 0: mux_10753 = 1'h0; 1: mux_10753 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10754;
  wire [0:0] v_10755;
  wire [0:0] v_10756;
  wire [0:0] v_10757;
  wire [0:0] v_10758;
  wire [0:0] v_10759;
  function [0:0] mux_10759(input [0:0] sel);
    case (sel) 0: mux_10759 = 1'h0; 1: mux_10759 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10760;
  wire [0:0] v_10761;
  wire [0:0] v_10762;
  wire [0:0] v_10763;
  wire [0:0] v_10764;
  function [0:0] mux_10764(input [0:0] sel);
    case (sel) 0: mux_10764 = 1'h0; 1: mux_10764 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10765;
  wire [0:0] v_10766;
  wire [0:0] v_10767;
  wire [0:0] v_10768;
  function [0:0] mux_10768(input [0:0] sel);
    case (sel) 0: mux_10768 = 1'h0; 1: mux_10768 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10769;
  function [0:0] mux_10769(input [0:0] sel);
    case (sel) 0: mux_10769 = 1'h0; 1: mux_10769 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_10770 = 1'h0;
  wire [0:0] v_10771;
  wire [0:0] v_10772;
  wire [0:0] act_10773;
  wire [0:0] v_10774;
  wire [0:0] v_10775;
  wire [0:0] v_10776;
  reg [0:0] v_10777 = 1'h0;
  wire [0:0] v_10778;
  wire [0:0] v_10779;
  wire [0:0] act_10780;
  wire [0:0] v_10781;
  wire [0:0] v_10782;
  wire [0:0] v_10783;
  wire [0:0] vin0_consume_en_10784;
  wire [0:0] vout_canPeek_10784;
  wire [7:0] vout_peek_10784;
  wire [0:0] v_10785;
  wire [0:0] v_10786;
  function [0:0] mux_10786(input [0:0] sel);
    case (sel) 0: mux_10786 = 1'h0; 1: mux_10786 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10787;
  wire [0:0] v_10788;
  wire [0:0] v_10789;
  wire [0:0] v_10790;
  wire [0:0] v_10791;
  function [0:0] mux_10791(input [0:0] sel);
    case (sel) 0: mux_10791 = 1'h0; 1: mux_10791 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10792;
  wire [0:0] vin0_consume_en_10793;
  wire [0:0] vout_canPeek_10793;
  wire [7:0] vout_peek_10793;
  wire [0:0] v_10794;
  wire [0:0] v_10795;
  function [0:0] mux_10795(input [0:0] sel);
    case (sel) 0: mux_10795 = 1'h0; 1: mux_10795 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10796;
  function [0:0] mux_10796(input [0:0] sel);
    case (sel) 0: mux_10796 = 1'h0; 1: mux_10796 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10797;
  wire [0:0] v_10798;
  wire [0:0] v_10799;
  wire [0:0] v_10800;
  wire [0:0] v_10801;
  wire [0:0] v_10802;
  wire [0:0] v_10803;
  function [0:0] mux_10803(input [0:0] sel);
    case (sel) 0: mux_10803 = 1'h0; 1: mux_10803 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10804;
  wire [0:0] v_10805;
  wire [0:0] v_10806;
  wire [0:0] v_10807;
  wire [0:0] v_10808;
  function [0:0] mux_10808(input [0:0] sel);
    case (sel) 0: mux_10808 = 1'h0; 1: mux_10808 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10809;
  wire [0:0] v_10810;
  wire [0:0] v_10811;
  wire [0:0] v_10812;
  function [0:0] mux_10812(input [0:0] sel);
    case (sel) 0: mux_10812 = 1'h0; 1: mux_10812 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10813;
  function [0:0] mux_10813(input [0:0] sel);
    case (sel) 0: mux_10813 = 1'h0; 1: mux_10813 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_10814 = 1'h0;
  wire [0:0] v_10815;
  wire [0:0] v_10816;
  wire [0:0] act_10817;
  wire [0:0] v_10818;
  wire [0:0] v_10819;
  wire [0:0] v_10820;
  wire [0:0] vin0_consume_en_10821;
  wire [0:0] vout_canPeek_10821;
  wire [7:0] vout_peek_10821;
  wire [0:0] v_10822;
  wire [0:0] v_10823;
  function [0:0] mux_10823(input [0:0] sel);
    case (sel) 0: mux_10823 = 1'h0; 1: mux_10823 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10824;
  wire [0:0] v_10825;
  wire [0:0] v_10826;
  wire [0:0] v_10827;
  wire [0:0] v_10828;
  function [0:0] mux_10828(input [0:0] sel);
    case (sel) 0: mux_10828 = 1'h0; 1: mux_10828 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10829;
  wire [0:0] vin0_consume_en_10830;
  wire [0:0] vout_canPeek_10830;
  wire [7:0] vout_peek_10830;
  wire [0:0] v_10831;
  wire [0:0] v_10832;
  function [0:0] mux_10832(input [0:0] sel);
    case (sel) 0: mux_10832 = 1'h0; 1: mux_10832 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10833;
  function [0:0] mux_10833(input [0:0] sel);
    case (sel) 0: mux_10833 = 1'h0; 1: mux_10833 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10834;
  wire [0:0] v_10835;
  wire [0:0] v_10836;
  wire [0:0] v_10837;
  wire [0:0] v_10838;
  wire [0:0] v_10839;
  wire [0:0] v_10840;
  function [0:0] mux_10840(input [0:0] sel);
    case (sel) 0: mux_10840 = 1'h0; 1: mux_10840 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10841;
  function [0:0] mux_10841(input [0:0] sel);
    case (sel) 0: mux_10841 = 1'h0; 1: mux_10841 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10842;
  wire [0:0] v_10843;
  wire [0:0] v_10844;
  wire [0:0] v_10845;
  function [0:0] mux_10845(input [0:0] sel);
    case (sel) 0: mux_10845 = 1'h0; 1: mux_10845 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10846;
  function [0:0] mux_10846(input [0:0] sel);
    case (sel) 0: mux_10846 = 1'h0; 1: mux_10846 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10847;
  wire [0:0] v_10848;
  wire [0:0] v_10849;
  wire [0:0] v_10850;
  wire [0:0] v_10851;
  wire [0:0] v_10852;
  function [0:0] mux_10852(input [0:0] sel);
    case (sel) 0: mux_10852 = 1'h0; 1: mux_10852 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10853;
  function [0:0] mux_10853(input [0:0] sel);
    case (sel) 0: mux_10853 = 1'h0; 1: mux_10853 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10854;
  wire [0:0] v_10855;
  wire [0:0] v_10856;
  wire [0:0] v_10857;
  function [0:0] mux_10857(input [0:0] sel);
    case (sel) 0: mux_10857 = 1'h0; 1: mux_10857 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10858;
  function [0:0] mux_10858(input [0:0] sel);
    case (sel) 0: mux_10858 = 1'h0; 1: mux_10858 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10859;
  wire [0:0] v_10860;
  wire [0:0] v_10861;
  wire [0:0] v_10862;
  wire [0:0] v_10863;
  wire [0:0] v_10864;
  function [0:0] mux_10864(input [0:0] sel);
    case (sel) 0: mux_10864 = 1'h0; 1: mux_10864 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10865;
  wire [0:0] v_10866;
  wire [0:0] v_10867;
  wire [0:0] v_10868;
  wire [0:0] v_10869;
  function [0:0] mux_10869(input [0:0] sel);
    case (sel) 0: mux_10869 = 1'h0; 1: mux_10869 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10870;
  wire [0:0] v_10871;
  wire [0:0] v_10872;
  wire [0:0] v_10873;
  function [0:0] mux_10873(input [0:0] sel);
    case (sel) 0: mux_10873 = 1'h0; 1: mux_10873 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10874;
  function [0:0] mux_10874(input [0:0] sel);
    case (sel) 0: mux_10874 = 1'h0; 1: mux_10874 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_10875 = 1'h0;
  wire [0:0] v_10876;
  wire [0:0] v_10877;
  wire [0:0] act_10878;
  wire [0:0] v_10879;
  wire [0:0] v_10880;
  wire [0:0] v_10881;
  reg [0:0] v_10882 = 1'h0;
  wire [0:0] v_10883;
  wire [0:0] v_10884;
  wire [0:0] act_10885;
  wire [0:0] v_10886;
  wire [0:0] v_10887;
  wire [0:0] v_10888;
  reg [0:0] v_10889 = 1'h0;
  wire [0:0] v_10890;
  wire [0:0] v_10891;
  wire [0:0] act_10892;
  wire [0:0] v_10893;
  wire [0:0] v_10894;
  wire [0:0] v_10895;
  wire [0:0] vin0_consume_en_10896;
  wire [0:0] vout_canPeek_10896;
  wire [7:0] vout_peek_10896;
  wire [0:0] v_10897;
  wire [0:0] v_10898;
  function [0:0] mux_10898(input [0:0] sel);
    case (sel) 0: mux_10898 = 1'h0; 1: mux_10898 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10899;
  wire [0:0] v_10900;
  wire [0:0] v_10901;
  wire [0:0] v_10902;
  wire [0:0] v_10903;
  function [0:0] mux_10903(input [0:0] sel);
    case (sel) 0: mux_10903 = 1'h0; 1: mux_10903 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10904;
  wire [0:0] vin0_consume_en_10905;
  wire [0:0] vout_canPeek_10905;
  wire [7:0] vout_peek_10905;
  wire [0:0] v_10906;
  wire [0:0] v_10907;
  function [0:0] mux_10907(input [0:0] sel);
    case (sel) 0: mux_10907 = 1'h0; 1: mux_10907 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10908;
  function [0:0] mux_10908(input [0:0] sel);
    case (sel) 0: mux_10908 = 1'h0; 1: mux_10908 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10909;
  wire [0:0] v_10910;
  wire [0:0] v_10911;
  wire [0:0] v_10912;
  wire [0:0] v_10913;
  wire [0:0] v_10914;
  wire [0:0] v_10915;
  function [0:0] mux_10915(input [0:0] sel);
    case (sel) 0: mux_10915 = 1'h0; 1: mux_10915 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10916;
  wire [0:0] v_10917;
  wire [0:0] v_10918;
  wire [0:0] v_10919;
  wire [0:0] v_10920;
  function [0:0] mux_10920(input [0:0] sel);
    case (sel) 0: mux_10920 = 1'h0; 1: mux_10920 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10921;
  wire [0:0] v_10922;
  wire [0:0] v_10923;
  wire [0:0] v_10924;
  function [0:0] mux_10924(input [0:0] sel);
    case (sel) 0: mux_10924 = 1'h0; 1: mux_10924 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10925;
  function [0:0] mux_10925(input [0:0] sel);
    case (sel) 0: mux_10925 = 1'h0; 1: mux_10925 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_10926 = 1'h0;
  wire [0:0] v_10927;
  wire [0:0] v_10928;
  wire [0:0] act_10929;
  wire [0:0] v_10930;
  wire [0:0] v_10931;
  wire [0:0] v_10932;
  wire [0:0] vin0_consume_en_10933;
  wire [0:0] vout_canPeek_10933;
  wire [7:0] vout_peek_10933;
  wire [0:0] v_10934;
  wire [0:0] v_10935;
  function [0:0] mux_10935(input [0:0] sel);
    case (sel) 0: mux_10935 = 1'h0; 1: mux_10935 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10936;
  wire [0:0] v_10937;
  wire [0:0] v_10938;
  wire [0:0] v_10939;
  wire [0:0] v_10940;
  function [0:0] mux_10940(input [0:0] sel);
    case (sel) 0: mux_10940 = 1'h0; 1: mux_10940 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10941;
  wire [0:0] vin0_consume_en_10942;
  wire [0:0] vout_canPeek_10942;
  wire [7:0] vout_peek_10942;
  wire [0:0] v_10943;
  wire [0:0] v_10944;
  function [0:0] mux_10944(input [0:0] sel);
    case (sel) 0: mux_10944 = 1'h0; 1: mux_10944 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10945;
  function [0:0] mux_10945(input [0:0] sel);
    case (sel) 0: mux_10945 = 1'h0; 1: mux_10945 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10946;
  wire [0:0] v_10947;
  wire [0:0] v_10948;
  wire [0:0] v_10949;
  wire [0:0] v_10950;
  wire [0:0] v_10951;
  wire [0:0] v_10952;
  function [0:0] mux_10952(input [0:0] sel);
    case (sel) 0: mux_10952 = 1'h0; 1: mux_10952 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10953;
  function [0:0] mux_10953(input [0:0] sel);
    case (sel) 0: mux_10953 = 1'h0; 1: mux_10953 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10954;
  wire [0:0] v_10955;
  wire [0:0] v_10956;
  wire [0:0] v_10957;
  function [0:0] mux_10957(input [0:0] sel);
    case (sel) 0: mux_10957 = 1'h0; 1: mux_10957 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10958;
  function [0:0] mux_10958(input [0:0] sel);
    case (sel) 0: mux_10958 = 1'h0; 1: mux_10958 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10959;
  wire [0:0] v_10960;
  wire [0:0] v_10961;
  wire [0:0] v_10962;
  wire [0:0] v_10963;
  wire [0:0] v_10964;
  function [0:0] mux_10964(input [0:0] sel);
    case (sel) 0: mux_10964 = 1'h0; 1: mux_10964 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10965;
  wire [0:0] v_10966;
  wire [0:0] v_10967;
  wire [0:0] v_10968;
  wire [0:0] v_10969;
  function [0:0] mux_10969(input [0:0] sel);
    case (sel) 0: mux_10969 = 1'h0; 1: mux_10969 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10970;
  wire [0:0] v_10971;
  wire [0:0] v_10972;
  wire [0:0] v_10973;
  function [0:0] mux_10973(input [0:0] sel);
    case (sel) 0: mux_10973 = 1'h0; 1: mux_10973 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10974;
  function [0:0] mux_10974(input [0:0] sel);
    case (sel) 0: mux_10974 = 1'h0; 1: mux_10974 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_10975 = 1'h0;
  wire [0:0] v_10976;
  wire [0:0] v_10977;
  wire [0:0] act_10978;
  wire [0:0] v_10979;
  wire [0:0] v_10980;
  wire [0:0] v_10981;
  reg [0:0] v_10982 = 1'h0;
  wire [0:0] v_10983;
  wire [0:0] v_10984;
  wire [0:0] act_10985;
  wire [0:0] v_10986;
  wire [0:0] v_10987;
  wire [0:0] v_10988;
  wire [0:0] vin0_consume_en_10989;
  wire [0:0] vout_canPeek_10989;
  wire [7:0] vout_peek_10989;
  wire [0:0] v_10990;
  wire [0:0] v_10991;
  function [0:0] mux_10991(input [0:0] sel);
    case (sel) 0: mux_10991 = 1'h0; 1: mux_10991 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_10992;
  wire [0:0] v_10993;
  wire [0:0] v_10994;
  wire [0:0] v_10995;
  wire [0:0] v_10996;
  function [0:0] mux_10996(input [0:0] sel);
    case (sel) 0: mux_10996 = 1'h0; 1: mux_10996 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_10997;
  wire [0:0] vin0_consume_en_10998;
  wire [0:0] vout_canPeek_10998;
  wire [7:0] vout_peek_10998;
  wire [0:0] v_10999;
  wire [0:0] v_11000;
  function [0:0] mux_11000(input [0:0] sel);
    case (sel) 0: mux_11000 = 1'h0; 1: mux_11000 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11001;
  function [0:0] mux_11001(input [0:0] sel);
    case (sel) 0: mux_11001 = 1'h0; 1: mux_11001 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11002;
  wire [0:0] v_11003;
  wire [0:0] v_11004;
  wire [0:0] v_11005;
  wire [0:0] v_11006;
  wire [0:0] v_11007;
  wire [0:0] v_11008;
  function [0:0] mux_11008(input [0:0] sel);
    case (sel) 0: mux_11008 = 1'h0; 1: mux_11008 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11009;
  wire [0:0] v_11010;
  wire [0:0] v_11011;
  wire [0:0] v_11012;
  wire [0:0] v_11013;
  function [0:0] mux_11013(input [0:0] sel);
    case (sel) 0: mux_11013 = 1'h0; 1: mux_11013 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11014;
  wire [0:0] v_11015;
  wire [0:0] v_11016;
  wire [0:0] v_11017;
  function [0:0] mux_11017(input [0:0] sel);
    case (sel) 0: mux_11017 = 1'h0; 1: mux_11017 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11018;
  function [0:0] mux_11018(input [0:0] sel);
    case (sel) 0: mux_11018 = 1'h0; 1: mux_11018 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_11019 = 1'h0;
  wire [0:0] v_11020;
  wire [0:0] v_11021;
  wire [0:0] act_11022;
  wire [0:0] v_11023;
  wire [0:0] v_11024;
  wire [0:0] v_11025;
  wire [0:0] vin0_consume_en_11026;
  wire [0:0] vout_canPeek_11026;
  wire [7:0] vout_peek_11026;
  wire [0:0] v_11027;
  wire [0:0] v_11028;
  function [0:0] mux_11028(input [0:0] sel);
    case (sel) 0: mux_11028 = 1'h0; 1: mux_11028 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11029;
  wire [0:0] v_11030;
  wire [0:0] v_11031;
  wire [0:0] v_11032;
  wire [0:0] v_11033;
  function [0:0] mux_11033(input [0:0] sel);
    case (sel) 0: mux_11033 = 1'h0; 1: mux_11033 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11034;
  wire [0:0] vin0_consume_en_11035;
  wire [0:0] vout_canPeek_11035;
  wire [7:0] vout_peek_11035;
  wire [0:0] v_11036;
  wire [0:0] v_11037;
  function [0:0] mux_11037(input [0:0] sel);
    case (sel) 0: mux_11037 = 1'h0; 1: mux_11037 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11038;
  function [0:0] mux_11038(input [0:0] sel);
    case (sel) 0: mux_11038 = 1'h0; 1: mux_11038 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11039;
  wire [0:0] v_11040;
  wire [0:0] v_11041;
  wire [0:0] v_11042;
  wire [0:0] v_11043;
  wire [0:0] v_11044;
  wire [0:0] v_11045;
  function [0:0] mux_11045(input [0:0] sel);
    case (sel) 0: mux_11045 = 1'h0; 1: mux_11045 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11046;
  function [0:0] mux_11046(input [0:0] sel);
    case (sel) 0: mux_11046 = 1'h0; 1: mux_11046 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11047;
  wire [0:0] v_11048;
  wire [0:0] v_11049;
  wire [0:0] v_11050;
  function [0:0] mux_11050(input [0:0] sel);
    case (sel) 0: mux_11050 = 1'h0; 1: mux_11050 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11051;
  function [0:0] mux_11051(input [0:0] sel);
    case (sel) 0: mux_11051 = 1'h0; 1: mux_11051 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11052;
  wire [0:0] v_11053;
  wire [0:0] v_11054;
  wire [0:0] v_11055;
  wire [0:0] v_11056;
  wire [0:0] v_11057;
  function [0:0] mux_11057(input [0:0] sel);
    case (sel) 0: mux_11057 = 1'h0; 1: mux_11057 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11058;
  function [0:0] mux_11058(input [0:0] sel);
    case (sel) 0: mux_11058 = 1'h0; 1: mux_11058 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11059;
  wire [0:0] v_11060;
  wire [0:0] v_11061;
  wire [0:0] v_11062;
  function [0:0] mux_11062(input [0:0] sel);
    case (sel) 0: mux_11062 = 1'h0; 1: mux_11062 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11063;
  function [0:0] mux_11063(input [0:0] sel);
    case (sel) 0: mux_11063 = 1'h0; 1: mux_11063 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11064;
  wire [0:0] v_11065;
  wire [0:0] v_11066;
  wire [0:0] v_11067;
  wire [0:0] v_11068;
  wire [0:0] v_11069;
  function [0:0] mux_11069(input [0:0] sel);
    case (sel) 0: mux_11069 = 1'h0; 1: mux_11069 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11070;
  function [0:0] mux_11070(input [0:0] sel);
    case (sel) 0: mux_11070 = 1'h0; 1: mux_11070 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11071;
  wire [0:0] v_11072;
  wire [0:0] v_11073;
  wire [0:0] v_11074;
  function [0:0] mux_11074(input [0:0] sel);
    case (sel) 0: mux_11074 = 1'h0; 1: mux_11074 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11075;
  function [0:0] mux_11075(input [0:0] sel);
    case (sel) 0: mux_11075 = 1'h0; 1: mux_11075 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11076;
  wire [0:0] v_11077;
  wire [0:0] v_11078;
  wire [0:0] v_11079;
  wire [0:0] v_11080;
  wire [0:0] v_11081;
  function [0:0] mux_11081(input [0:0] sel);
    case (sel) 0: mux_11081 = 1'h0; 1: mux_11081 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11082;
  wire [0:0] v_11083;
  wire [0:0] v_11084;
  wire [0:0] v_11085;
  wire [0:0] v_11086;
  function [0:0] mux_11086(input [0:0] sel);
    case (sel) 0: mux_11086 = 1'h0; 1: mux_11086 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11087;
  wire [0:0] v_11088;
  wire [0:0] v_11089;
  wire [0:0] v_11090;
  function [0:0] mux_11090(input [0:0] sel);
    case (sel) 0: mux_11090 = 1'h0; 1: mux_11090 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11091;
  function [0:0] mux_11091(input [0:0] sel);
    case (sel) 0: mux_11091 = 1'h0; 1: mux_11091 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_11092 = 1'h0;
  wire [0:0] v_11093;
  wire [0:0] v_11094;
  wire [0:0] act_11095;
  wire [0:0] v_11096;
  wire [0:0] v_11097;
  wire [0:0] v_11098;
  reg [0:0] v_11099 = 1'h0;
  wire [0:0] v_11100;
  wire [0:0] v_11101;
  wire [0:0] act_11102;
  wire [0:0] v_11103;
  wire [0:0] v_11104;
  wire [0:0] v_11105;
  reg [0:0] v_11106 = 1'h0;
  wire [0:0] v_11107;
  wire [0:0] v_11108;
  wire [0:0] act_11109;
  wire [0:0] v_11110;
  wire [0:0] v_11111;
  wire [0:0] v_11112;
  reg [0:0] v_11113 = 1'h0;
  wire [0:0] v_11114;
  wire [0:0] v_11115;
  wire [0:0] act_11116;
  wire [0:0] v_11117;
  wire [0:0] v_11118;
  wire [0:0] v_11119;
  wire [0:0] vin0_consume_en_11120;
  wire [0:0] vout_canPeek_11120;
  wire [7:0] vout_peek_11120;
  wire [0:0] v_11121;
  wire [0:0] v_11122;
  function [0:0] mux_11122(input [0:0] sel);
    case (sel) 0: mux_11122 = 1'h0; 1: mux_11122 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11123;
  wire [0:0] v_11124;
  wire [0:0] v_11125;
  wire [0:0] v_11126;
  wire [0:0] v_11127;
  function [0:0] mux_11127(input [0:0] sel);
    case (sel) 0: mux_11127 = 1'h0; 1: mux_11127 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11128;
  wire [0:0] vin0_consume_en_11129;
  wire [0:0] vout_canPeek_11129;
  wire [7:0] vout_peek_11129;
  wire [0:0] v_11130;
  wire [0:0] v_11131;
  function [0:0] mux_11131(input [0:0] sel);
    case (sel) 0: mux_11131 = 1'h0; 1: mux_11131 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11132;
  function [0:0] mux_11132(input [0:0] sel);
    case (sel) 0: mux_11132 = 1'h0; 1: mux_11132 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11133;
  wire [0:0] v_11134;
  wire [0:0] v_11135;
  wire [0:0] v_11136;
  wire [0:0] v_11137;
  wire [0:0] v_11138;
  wire [0:0] v_11139;
  function [0:0] mux_11139(input [0:0] sel);
    case (sel) 0: mux_11139 = 1'h0; 1: mux_11139 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11140;
  wire [0:0] v_11141;
  wire [0:0] v_11142;
  wire [0:0] v_11143;
  wire [0:0] v_11144;
  function [0:0] mux_11144(input [0:0] sel);
    case (sel) 0: mux_11144 = 1'h0; 1: mux_11144 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11145;
  wire [0:0] v_11146;
  wire [0:0] v_11147;
  wire [0:0] v_11148;
  function [0:0] mux_11148(input [0:0] sel);
    case (sel) 0: mux_11148 = 1'h0; 1: mux_11148 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11149;
  function [0:0] mux_11149(input [0:0] sel);
    case (sel) 0: mux_11149 = 1'h0; 1: mux_11149 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_11150 = 1'h0;
  wire [0:0] v_11151;
  wire [0:0] v_11152;
  wire [0:0] act_11153;
  wire [0:0] v_11154;
  wire [0:0] v_11155;
  wire [0:0] v_11156;
  wire [0:0] vin0_consume_en_11157;
  wire [0:0] vout_canPeek_11157;
  wire [7:0] vout_peek_11157;
  wire [0:0] v_11158;
  wire [0:0] v_11159;
  function [0:0] mux_11159(input [0:0] sel);
    case (sel) 0: mux_11159 = 1'h0; 1: mux_11159 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11160;
  wire [0:0] v_11161;
  wire [0:0] v_11162;
  wire [0:0] v_11163;
  wire [0:0] v_11164;
  function [0:0] mux_11164(input [0:0] sel);
    case (sel) 0: mux_11164 = 1'h0; 1: mux_11164 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11165;
  wire [0:0] vin0_consume_en_11166;
  wire [0:0] vout_canPeek_11166;
  wire [7:0] vout_peek_11166;
  wire [0:0] v_11167;
  wire [0:0] v_11168;
  function [0:0] mux_11168(input [0:0] sel);
    case (sel) 0: mux_11168 = 1'h0; 1: mux_11168 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11169;
  function [0:0] mux_11169(input [0:0] sel);
    case (sel) 0: mux_11169 = 1'h0; 1: mux_11169 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11170;
  wire [0:0] v_11171;
  wire [0:0] v_11172;
  wire [0:0] v_11173;
  wire [0:0] v_11174;
  wire [0:0] v_11175;
  wire [0:0] v_11176;
  function [0:0] mux_11176(input [0:0] sel);
    case (sel) 0: mux_11176 = 1'h0; 1: mux_11176 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11177;
  function [0:0] mux_11177(input [0:0] sel);
    case (sel) 0: mux_11177 = 1'h0; 1: mux_11177 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11178;
  wire [0:0] v_11179;
  wire [0:0] v_11180;
  wire [0:0] v_11181;
  function [0:0] mux_11181(input [0:0] sel);
    case (sel) 0: mux_11181 = 1'h0; 1: mux_11181 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11182;
  function [0:0] mux_11182(input [0:0] sel);
    case (sel) 0: mux_11182 = 1'h0; 1: mux_11182 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11183;
  wire [0:0] v_11184;
  wire [0:0] v_11185;
  wire [0:0] v_11186;
  wire [0:0] v_11187;
  wire [0:0] v_11188;
  function [0:0] mux_11188(input [0:0] sel);
    case (sel) 0: mux_11188 = 1'h0; 1: mux_11188 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11189;
  wire [0:0] v_11190;
  wire [0:0] v_11191;
  wire [0:0] v_11192;
  wire [0:0] v_11193;
  function [0:0] mux_11193(input [0:0] sel);
    case (sel) 0: mux_11193 = 1'h0; 1: mux_11193 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11194;
  wire [0:0] v_11195;
  wire [0:0] v_11196;
  wire [0:0] v_11197;
  function [0:0] mux_11197(input [0:0] sel);
    case (sel) 0: mux_11197 = 1'h0; 1: mux_11197 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11198;
  function [0:0] mux_11198(input [0:0] sel);
    case (sel) 0: mux_11198 = 1'h0; 1: mux_11198 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_11199 = 1'h0;
  wire [0:0] v_11200;
  wire [0:0] v_11201;
  wire [0:0] act_11202;
  wire [0:0] v_11203;
  wire [0:0] v_11204;
  wire [0:0] v_11205;
  reg [0:0] v_11206 = 1'h0;
  wire [0:0] v_11207;
  wire [0:0] v_11208;
  wire [0:0] act_11209;
  wire [0:0] v_11210;
  wire [0:0] v_11211;
  wire [0:0] v_11212;
  wire [0:0] vin0_consume_en_11213;
  wire [0:0] vout_canPeek_11213;
  wire [7:0] vout_peek_11213;
  wire [0:0] v_11214;
  wire [0:0] v_11215;
  function [0:0] mux_11215(input [0:0] sel);
    case (sel) 0: mux_11215 = 1'h0; 1: mux_11215 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11216;
  wire [0:0] v_11217;
  wire [0:0] v_11218;
  wire [0:0] v_11219;
  wire [0:0] v_11220;
  function [0:0] mux_11220(input [0:0] sel);
    case (sel) 0: mux_11220 = 1'h0; 1: mux_11220 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11221;
  wire [0:0] vin0_consume_en_11222;
  wire [0:0] vout_canPeek_11222;
  wire [7:0] vout_peek_11222;
  wire [0:0] v_11223;
  wire [0:0] v_11224;
  function [0:0] mux_11224(input [0:0] sel);
    case (sel) 0: mux_11224 = 1'h0; 1: mux_11224 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11225;
  function [0:0] mux_11225(input [0:0] sel);
    case (sel) 0: mux_11225 = 1'h0; 1: mux_11225 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11226;
  wire [0:0] v_11227;
  wire [0:0] v_11228;
  wire [0:0] v_11229;
  wire [0:0] v_11230;
  wire [0:0] v_11231;
  wire [0:0] v_11232;
  function [0:0] mux_11232(input [0:0] sel);
    case (sel) 0: mux_11232 = 1'h0; 1: mux_11232 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11233;
  wire [0:0] v_11234;
  wire [0:0] v_11235;
  wire [0:0] v_11236;
  wire [0:0] v_11237;
  function [0:0] mux_11237(input [0:0] sel);
    case (sel) 0: mux_11237 = 1'h0; 1: mux_11237 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11238;
  wire [0:0] v_11239;
  wire [0:0] v_11240;
  wire [0:0] v_11241;
  function [0:0] mux_11241(input [0:0] sel);
    case (sel) 0: mux_11241 = 1'h0; 1: mux_11241 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11242;
  function [0:0] mux_11242(input [0:0] sel);
    case (sel) 0: mux_11242 = 1'h0; 1: mux_11242 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_11243 = 1'h0;
  wire [0:0] v_11244;
  wire [0:0] v_11245;
  wire [0:0] act_11246;
  wire [0:0] v_11247;
  wire [0:0] v_11248;
  wire [0:0] v_11249;
  wire [0:0] vin0_consume_en_11250;
  wire [0:0] vout_canPeek_11250;
  wire [7:0] vout_peek_11250;
  wire [0:0] v_11251;
  wire [0:0] v_11252;
  function [0:0] mux_11252(input [0:0] sel);
    case (sel) 0: mux_11252 = 1'h0; 1: mux_11252 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11253;
  wire [0:0] v_11254;
  wire [0:0] v_11255;
  wire [0:0] v_11256;
  wire [0:0] v_11257;
  function [0:0] mux_11257(input [0:0] sel);
    case (sel) 0: mux_11257 = 1'h0; 1: mux_11257 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11258;
  wire [0:0] vin0_consume_en_11259;
  wire [0:0] vout_canPeek_11259;
  wire [7:0] vout_peek_11259;
  wire [0:0] v_11260;
  wire [0:0] v_11261;
  function [0:0] mux_11261(input [0:0] sel);
    case (sel) 0: mux_11261 = 1'h0; 1: mux_11261 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11262;
  function [0:0] mux_11262(input [0:0] sel);
    case (sel) 0: mux_11262 = 1'h0; 1: mux_11262 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11263;
  wire [0:0] v_11264;
  wire [0:0] v_11265;
  wire [0:0] v_11266;
  wire [0:0] v_11267;
  wire [0:0] v_11268;
  wire [0:0] v_11269;
  function [0:0] mux_11269(input [0:0] sel);
    case (sel) 0: mux_11269 = 1'h0; 1: mux_11269 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11270;
  function [0:0] mux_11270(input [0:0] sel);
    case (sel) 0: mux_11270 = 1'h0; 1: mux_11270 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11271;
  wire [0:0] v_11272;
  wire [0:0] v_11273;
  wire [0:0] v_11274;
  function [0:0] mux_11274(input [0:0] sel);
    case (sel) 0: mux_11274 = 1'h0; 1: mux_11274 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11275;
  function [0:0] mux_11275(input [0:0] sel);
    case (sel) 0: mux_11275 = 1'h0; 1: mux_11275 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11276;
  wire [0:0] v_11277;
  wire [0:0] v_11278;
  wire [0:0] v_11279;
  wire [0:0] v_11280;
  wire [0:0] v_11281;
  function [0:0] mux_11281(input [0:0] sel);
    case (sel) 0: mux_11281 = 1'h0; 1: mux_11281 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11282;
  function [0:0] mux_11282(input [0:0] sel);
    case (sel) 0: mux_11282 = 1'h0; 1: mux_11282 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11283;
  wire [0:0] v_11284;
  wire [0:0] v_11285;
  wire [0:0] v_11286;
  function [0:0] mux_11286(input [0:0] sel);
    case (sel) 0: mux_11286 = 1'h0; 1: mux_11286 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11287;
  function [0:0] mux_11287(input [0:0] sel);
    case (sel) 0: mux_11287 = 1'h0; 1: mux_11287 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11288;
  wire [0:0] v_11289;
  wire [0:0] v_11290;
  wire [0:0] v_11291;
  wire [0:0] v_11292;
  wire [0:0] v_11293;
  function [0:0] mux_11293(input [0:0] sel);
    case (sel) 0: mux_11293 = 1'h0; 1: mux_11293 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11294;
  wire [0:0] v_11295;
  wire [0:0] v_11296;
  wire [0:0] v_11297;
  wire [0:0] v_11298;
  function [0:0] mux_11298(input [0:0] sel);
    case (sel) 0: mux_11298 = 1'h0; 1: mux_11298 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11299;
  wire [0:0] v_11300;
  wire [0:0] v_11301;
  wire [0:0] v_11302;
  function [0:0] mux_11302(input [0:0] sel);
    case (sel) 0: mux_11302 = 1'h0; 1: mux_11302 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11303;
  function [0:0] mux_11303(input [0:0] sel);
    case (sel) 0: mux_11303 = 1'h0; 1: mux_11303 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_11304 = 1'h0;
  wire [0:0] v_11305;
  wire [0:0] v_11306;
  wire [0:0] act_11307;
  wire [0:0] v_11308;
  wire [0:0] v_11309;
  wire [0:0] v_11310;
  reg [0:0] v_11311 = 1'h0;
  wire [0:0] v_11312;
  wire [0:0] v_11313;
  wire [0:0] act_11314;
  wire [0:0] v_11315;
  wire [0:0] v_11316;
  wire [0:0] v_11317;
  reg [0:0] v_11318 = 1'h0;
  wire [0:0] v_11319;
  wire [0:0] v_11320;
  wire [0:0] act_11321;
  wire [0:0] v_11322;
  wire [0:0] v_11323;
  wire [0:0] v_11324;
  wire [0:0] vin0_consume_en_11325;
  wire [0:0] vout_canPeek_11325;
  wire [7:0] vout_peek_11325;
  wire [0:0] v_11326;
  wire [0:0] v_11327;
  function [0:0] mux_11327(input [0:0] sel);
    case (sel) 0: mux_11327 = 1'h0; 1: mux_11327 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11328;
  wire [0:0] v_11329;
  wire [0:0] v_11330;
  wire [0:0] v_11331;
  wire [0:0] v_11332;
  function [0:0] mux_11332(input [0:0] sel);
    case (sel) 0: mux_11332 = 1'h0; 1: mux_11332 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11333;
  wire [0:0] vin0_consume_en_11334;
  wire [0:0] vout_canPeek_11334;
  wire [7:0] vout_peek_11334;
  wire [0:0] v_11335;
  wire [0:0] v_11336;
  function [0:0] mux_11336(input [0:0] sel);
    case (sel) 0: mux_11336 = 1'h0; 1: mux_11336 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11337;
  function [0:0] mux_11337(input [0:0] sel);
    case (sel) 0: mux_11337 = 1'h0; 1: mux_11337 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11338;
  wire [0:0] v_11339;
  wire [0:0] v_11340;
  wire [0:0] v_11341;
  wire [0:0] v_11342;
  wire [0:0] v_11343;
  wire [0:0] v_11344;
  function [0:0] mux_11344(input [0:0] sel);
    case (sel) 0: mux_11344 = 1'h0; 1: mux_11344 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11345;
  wire [0:0] v_11346;
  wire [0:0] v_11347;
  wire [0:0] v_11348;
  wire [0:0] v_11349;
  function [0:0] mux_11349(input [0:0] sel);
    case (sel) 0: mux_11349 = 1'h0; 1: mux_11349 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11350;
  wire [0:0] v_11351;
  wire [0:0] v_11352;
  wire [0:0] v_11353;
  function [0:0] mux_11353(input [0:0] sel);
    case (sel) 0: mux_11353 = 1'h0; 1: mux_11353 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11354;
  function [0:0] mux_11354(input [0:0] sel);
    case (sel) 0: mux_11354 = 1'h0; 1: mux_11354 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_11355 = 1'h0;
  wire [0:0] v_11356;
  wire [0:0] v_11357;
  wire [0:0] act_11358;
  wire [0:0] v_11359;
  wire [0:0] v_11360;
  wire [0:0] v_11361;
  wire [0:0] vin0_consume_en_11362;
  wire [0:0] vout_canPeek_11362;
  wire [7:0] vout_peek_11362;
  wire [0:0] v_11363;
  wire [0:0] v_11364;
  function [0:0] mux_11364(input [0:0] sel);
    case (sel) 0: mux_11364 = 1'h0; 1: mux_11364 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11365;
  wire [0:0] v_11366;
  wire [0:0] v_11367;
  wire [0:0] v_11368;
  wire [0:0] v_11369;
  function [0:0] mux_11369(input [0:0] sel);
    case (sel) 0: mux_11369 = 1'h0; 1: mux_11369 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11370;
  wire [0:0] vin0_consume_en_11371;
  wire [0:0] vout_canPeek_11371;
  wire [7:0] vout_peek_11371;
  wire [0:0] v_11372;
  wire [0:0] v_11373;
  function [0:0] mux_11373(input [0:0] sel);
    case (sel) 0: mux_11373 = 1'h0; 1: mux_11373 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11374;
  function [0:0] mux_11374(input [0:0] sel);
    case (sel) 0: mux_11374 = 1'h0; 1: mux_11374 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11375;
  wire [0:0] v_11376;
  wire [0:0] v_11377;
  wire [0:0] v_11378;
  wire [0:0] v_11379;
  wire [0:0] v_11380;
  wire [0:0] v_11381;
  function [0:0] mux_11381(input [0:0] sel);
    case (sel) 0: mux_11381 = 1'h0; 1: mux_11381 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11382;
  function [0:0] mux_11382(input [0:0] sel);
    case (sel) 0: mux_11382 = 1'h0; 1: mux_11382 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11383;
  wire [0:0] v_11384;
  wire [0:0] v_11385;
  wire [0:0] v_11386;
  function [0:0] mux_11386(input [0:0] sel);
    case (sel) 0: mux_11386 = 1'h0; 1: mux_11386 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11387;
  function [0:0] mux_11387(input [0:0] sel);
    case (sel) 0: mux_11387 = 1'h0; 1: mux_11387 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11388;
  wire [0:0] v_11389;
  wire [0:0] v_11390;
  wire [0:0] v_11391;
  wire [0:0] v_11392;
  wire [0:0] v_11393;
  function [0:0] mux_11393(input [0:0] sel);
    case (sel) 0: mux_11393 = 1'h0; 1: mux_11393 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11394;
  wire [0:0] v_11395;
  wire [0:0] v_11396;
  wire [0:0] v_11397;
  wire [0:0] v_11398;
  function [0:0] mux_11398(input [0:0] sel);
    case (sel) 0: mux_11398 = 1'h0; 1: mux_11398 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11399;
  wire [0:0] v_11400;
  wire [0:0] v_11401;
  wire [0:0] v_11402;
  function [0:0] mux_11402(input [0:0] sel);
    case (sel) 0: mux_11402 = 1'h0; 1: mux_11402 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11403;
  function [0:0] mux_11403(input [0:0] sel);
    case (sel) 0: mux_11403 = 1'h0; 1: mux_11403 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_11404 = 1'h0;
  wire [0:0] v_11405;
  wire [0:0] v_11406;
  wire [0:0] act_11407;
  wire [0:0] v_11408;
  wire [0:0] v_11409;
  wire [0:0] v_11410;
  reg [0:0] v_11411 = 1'h0;
  wire [0:0] v_11412;
  wire [0:0] v_11413;
  wire [0:0] act_11414;
  wire [0:0] v_11415;
  wire [0:0] v_11416;
  wire [0:0] v_11417;
  wire [0:0] vin0_consume_en_11418;
  wire [0:0] vout_canPeek_11418;
  wire [7:0] vout_peek_11418;
  wire [0:0] v_11419;
  wire [0:0] v_11420;
  function [0:0] mux_11420(input [0:0] sel);
    case (sel) 0: mux_11420 = 1'h0; 1: mux_11420 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11421;
  wire [0:0] v_11422;
  wire [0:0] v_11423;
  wire [0:0] v_11424;
  wire [0:0] v_11425;
  function [0:0] mux_11425(input [0:0] sel);
    case (sel) 0: mux_11425 = 1'h0; 1: mux_11425 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11426;
  wire [0:0] vin0_consume_en_11427;
  wire [0:0] vout_canPeek_11427;
  wire [7:0] vout_peek_11427;
  wire [0:0] v_11428;
  wire [0:0] v_11429;
  function [0:0] mux_11429(input [0:0] sel);
    case (sel) 0: mux_11429 = 1'h0; 1: mux_11429 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11430;
  function [0:0] mux_11430(input [0:0] sel);
    case (sel) 0: mux_11430 = 1'h0; 1: mux_11430 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11431;
  wire [0:0] v_11432;
  wire [0:0] v_11433;
  wire [0:0] v_11434;
  wire [0:0] v_11435;
  wire [0:0] v_11436;
  wire [0:0] v_11437;
  function [0:0] mux_11437(input [0:0] sel);
    case (sel) 0: mux_11437 = 1'h0; 1: mux_11437 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11438;
  wire [0:0] v_11439;
  wire [0:0] v_11440;
  wire [0:0] v_11441;
  wire [0:0] v_11442;
  function [0:0] mux_11442(input [0:0] sel);
    case (sel) 0: mux_11442 = 1'h0; 1: mux_11442 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11443;
  wire [0:0] v_11444;
  wire [0:0] v_11445;
  wire [0:0] v_11446;
  function [0:0] mux_11446(input [0:0] sel);
    case (sel) 0: mux_11446 = 1'h0; 1: mux_11446 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11447;
  function [0:0] mux_11447(input [0:0] sel);
    case (sel) 0: mux_11447 = 1'h0; 1: mux_11447 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_11448 = 1'h0;
  wire [0:0] v_11449;
  wire [0:0] v_11450;
  wire [0:0] act_11451;
  wire [0:0] v_11452;
  wire [0:0] v_11453;
  wire [0:0] v_11454;
  wire [0:0] vin0_consume_en_11455;
  wire [0:0] vout_canPeek_11455;
  wire [7:0] vout_peek_11455;
  wire [0:0] v_11456;
  wire [0:0] v_11457;
  function [0:0] mux_11457(input [0:0] sel);
    case (sel) 0: mux_11457 = 1'h0; 1: mux_11457 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11458;
  wire [0:0] v_11459;
  wire [0:0] v_11460;
  wire [0:0] v_11461;
  wire [0:0] v_11462;
  function [0:0] mux_11462(input [0:0] sel);
    case (sel) 0: mux_11462 = 1'h0; 1: mux_11462 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11463;
  wire [0:0] vin0_consume_en_11464;
  wire [0:0] vout_canPeek_11464;
  wire [7:0] vout_peek_11464;
  wire [0:0] v_11465;
  wire [0:0] v_11466;
  function [0:0] mux_11466(input [0:0] sel);
    case (sel) 0: mux_11466 = 1'h0; 1: mux_11466 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11467;
  function [0:0] mux_11467(input [0:0] sel);
    case (sel) 0: mux_11467 = 1'h0; 1: mux_11467 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11468;
  wire [0:0] v_11469;
  wire [0:0] v_11470;
  wire [0:0] v_11471;
  wire [0:0] v_11472;
  wire [0:0] v_11473;
  wire [0:0] v_11474;
  function [0:0] mux_11474(input [0:0] sel);
    case (sel) 0: mux_11474 = 1'h0; 1: mux_11474 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11475;
  function [0:0] mux_11475(input [0:0] sel);
    case (sel) 0: mux_11475 = 1'h0; 1: mux_11475 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11476;
  wire [0:0] v_11477;
  wire [0:0] v_11478;
  wire [0:0] v_11479;
  function [0:0] mux_11479(input [0:0] sel);
    case (sel) 0: mux_11479 = 1'h0; 1: mux_11479 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11480;
  function [0:0] mux_11480(input [0:0] sel);
    case (sel) 0: mux_11480 = 1'h0; 1: mux_11480 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11481;
  wire [0:0] v_11482;
  wire [0:0] v_11483;
  wire [0:0] v_11484;
  wire [0:0] v_11485;
  wire [0:0] v_11486;
  function [0:0] mux_11486(input [0:0] sel);
    case (sel) 0: mux_11486 = 1'h0; 1: mux_11486 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11487;
  function [0:0] mux_11487(input [0:0] sel);
    case (sel) 0: mux_11487 = 1'h0; 1: mux_11487 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11488;
  wire [0:0] v_11489;
  wire [0:0] v_11490;
  wire [0:0] v_11491;
  function [0:0] mux_11491(input [0:0] sel);
    case (sel) 0: mux_11491 = 1'h0; 1: mux_11491 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11492;
  function [0:0] mux_11492(input [0:0] sel);
    case (sel) 0: mux_11492 = 1'h0; 1: mux_11492 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11493;
  wire [0:0] v_11494;
  wire [0:0] v_11495;
  wire [0:0] v_11496;
  wire [0:0] v_11497;
  wire [0:0] v_11498;
  function [0:0] mux_11498(input [0:0] sel);
    case (sel) 0: mux_11498 = 1'h0; 1: mux_11498 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11499;
  function [0:0] mux_11499(input [0:0] sel);
    case (sel) 0: mux_11499 = 1'h0; 1: mux_11499 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11500;
  wire [0:0] v_11501;
  wire [0:0] v_11502;
  wire [0:0] v_11503;
  function [0:0] mux_11503(input [0:0] sel);
    case (sel) 0: mux_11503 = 1'h0; 1: mux_11503 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11504;
  function [0:0] mux_11504(input [0:0] sel);
    case (sel) 0: mux_11504 = 1'h0; 1: mux_11504 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11505;
  wire [0:0] v_11506;
  wire [0:0] v_11507;
  wire [0:0] v_11508;
  wire [0:0] v_11509;
  wire [0:0] v_11510;
  function [0:0] mux_11510(input [0:0] sel);
    case (sel) 0: mux_11510 = 1'h0; 1: mux_11510 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11511;
  function [0:0] mux_11511(input [0:0] sel);
    case (sel) 0: mux_11511 = 1'h0; 1: mux_11511 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11512;
  wire [0:0] v_11513;
  wire [0:0] v_11514;
  wire [0:0] v_11515;
  function [0:0] mux_11515(input [0:0] sel);
    case (sel) 0: mux_11515 = 1'h0; 1: mux_11515 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11516;
  function [0:0] mux_11516(input [0:0] sel);
    case (sel) 0: mux_11516 = 1'h0; 1: mux_11516 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11517;
  wire [0:0] v_11518;
  wire [0:0] v_11519;
  wire [0:0] v_11520;
  wire [0:0] v_11521;
  wire [0:0] v_11522;
  function [0:0] mux_11522(input [0:0] sel);
    case (sel) 0: mux_11522 = 1'h0; 1: mux_11522 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11523;
  function [0:0] mux_11523(input [0:0] sel);
    case (sel) 0: mux_11523 = 1'h0; 1: mux_11523 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11524;
  wire [0:0] v_11525;
  wire [0:0] v_11526;
  wire [0:0] v_11527;
  function [0:0] mux_11527(input [0:0] sel);
    case (sel) 0: mux_11527 = 1'h0; 1: mux_11527 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11528;
  function [0:0] mux_11528(input [0:0] sel);
    case (sel) 0: mux_11528 = 1'h0; 1: mux_11528 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11529;
  wire [0:0] v_11530;
  wire [0:0] v_11531;
  wire [0:0] v_11532;
  wire [0:0] v_11533;
  wire [0:0] v_11534;
  function [0:0] mux_11534(input [0:0] sel);
    case (sel) 0: mux_11534 = 1'h0; 1: mux_11534 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11535;
  function [0:0] mux_11535(input [0:0] sel);
    case (sel) 0: mux_11535 = 1'h0; 1: mux_11535 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11536;
  wire [0:0] v_11537;
  wire [0:0] v_11538;
  wire [0:0] v_11539;
  function [0:0] mux_11539(input [0:0] sel);
    case (sel) 0: mux_11539 = 1'h0; 1: mux_11539 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11540;
  function [0:0] mux_11540(input [0:0] sel);
    case (sel) 0: mux_11540 = 1'h0; 1: mux_11540 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11541;
  wire [0:0] v_11542;
  wire [0:0] v_11543;
  wire [0:0] v_11544;
  wire [0:0] v_11545;
  wire [0:0] v_11546;
  function [0:0] mux_11546(input [0:0] sel);
    case (sel) 0: mux_11546 = 1'h0; 1: mux_11546 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11547;
  wire [0:0] v_11548;
  wire [0:0] v_11549;
  wire [0:0] v_11550;
  wire [0:0] v_11551;
  function [0:0] mux_11551(input [0:0] sel);
    case (sel) 0: mux_11551 = 1'h0; 1: mux_11551 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11552;
  wire [0:0] v_11553;
  wire [0:0] v_11554;
  wire [0:0] v_11555;
  function [0:0] mux_11555(input [0:0] sel);
    case (sel) 0: mux_11555 = 1'h0; 1: mux_11555 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11556;
  function [0:0] mux_11556(input [0:0] sel);
    case (sel) 0: mux_11556 = 1'h0; 1: mux_11556 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_11557 = 1'h0;
  wire [0:0] v_11558;
  wire [0:0] v_11559;
  wire [0:0] act_11560;
  wire [0:0] v_11561;
  wire [0:0] v_11562;
  wire [0:0] v_11563;
  reg [0:0] v_11564 = 1'h0;
  wire [0:0] v_11565;
  wire [0:0] v_11566;
  wire [0:0] act_11567;
  wire [0:0] v_11568;
  wire [0:0] v_11569;
  wire [0:0] v_11570;
  reg [0:0] v_11571 = 1'h0;
  wire [0:0] v_11572;
  wire [0:0] v_11573;
  wire [0:0] act_11574;
  wire [0:0] v_11575;
  wire [0:0] v_11576;
  wire [0:0] v_11577;
  reg [0:0] v_11578 = 1'h0;
  wire [0:0] v_11579;
  wire [0:0] v_11580;
  wire [0:0] act_11581;
  wire [0:0] v_11582;
  wire [0:0] v_11583;
  wire [0:0] v_11584;
  reg [0:0] v_11585 = 1'h0;
  wire [0:0] v_11586;
  wire [0:0] v_11587;
  wire [0:0] act_11588;
  wire [0:0] v_11589;
  wire [0:0] v_11590;
  wire [0:0] v_11591;
  reg [0:0] v_11592 = 1'h0;
  wire [0:0] v_11593;
  wire [0:0] v_11594;
  wire [0:0] act_11595;
  wire [0:0] v_11596;
  wire [0:0] v_11597;
  wire [0:0] v_11598;
  reg [0:0] v_11599 = 1'h0;
  wire [0:0] v_11600;
  wire [0:0] v_11601;
  wire [0:0] act_11602;
  wire [0:0] v_11603;
  wire [0:0] v_11604;
  wire [0:0] v_11605;
  wire [0:0] vin0_consume_en_11606;
  wire [0:0] vout_canPeek_11606;
  wire [7:0] vout_peek_11606;
  wire [0:0] v_11607;
  wire [0:0] v_11608;
  function [0:0] mux_11608(input [0:0] sel);
    case (sel) 0: mux_11608 = 1'h0; 1: mux_11608 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11609;
  wire [0:0] v_11610;
  wire [0:0] v_11611;
  wire [0:0] v_11612;
  wire [0:0] v_11613;
  function [0:0] mux_11613(input [0:0] sel);
    case (sel) 0: mux_11613 = 1'h0; 1: mux_11613 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11614;
  wire [0:0] vin0_consume_en_11615;
  wire [0:0] vout_canPeek_11615;
  wire [7:0] vout_peek_11615;
  wire [0:0] v_11616;
  wire [0:0] v_11617;
  function [0:0] mux_11617(input [0:0] sel);
    case (sel) 0: mux_11617 = 1'h0; 1: mux_11617 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11618;
  function [0:0] mux_11618(input [0:0] sel);
    case (sel) 0: mux_11618 = 1'h0; 1: mux_11618 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11619;
  wire [0:0] v_11620;
  wire [0:0] v_11621;
  wire [0:0] v_11622;
  wire [0:0] v_11623;
  wire [0:0] v_11624;
  wire [0:0] v_11625;
  function [0:0] mux_11625(input [0:0] sel);
    case (sel) 0: mux_11625 = 1'h0; 1: mux_11625 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11626;
  wire [0:0] v_11627;
  wire [0:0] v_11628;
  wire [0:0] v_11629;
  wire [0:0] v_11630;
  function [0:0] mux_11630(input [0:0] sel);
    case (sel) 0: mux_11630 = 1'h0; 1: mux_11630 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11631;
  wire [0:0] v_11632;
  wire [0:0] v_11633;
  wire [0:0] v_11634;
  function [0:0] mux_11634(input [0:0] sel);
    case (sel) 0: mux_11634 = 1'h0; 1: mux_11634 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11635;
  function [0:0] mux_11635(input [0:0] sel);
    case (sel) 0: mux_11635 = 1'h0; 1: mux_11635 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_11636 = 1'h0;
  wire [0:0] v_11637;
  wire [0:0] v_11638;
  wire [0:0] act_11639;
  wire [0:0] v_11640;
  wire [0:0] v_11641;
  wire [0:0] v_11642;
  wire [0:0] vin0_consume_en_11643;
  wire [0:0] vout_canPeek_11643;
  wire [7:0] vout_peek_11643;
  wire [0:0] v_11644;
  wire [0:0] v_11645;
  function [0:0] mux_11645(input [0:0] sel);
    case (sel) 0: mux_11645 = 1'h0; 1: mux_11645 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11646;
  wire [0:0] v_11647;
  wire [0:0] v_11648;
  wire [0:0] v_11649;
  wire [0:0] v_11650;
  function [0:0] mux_11650(input [0:0] sel);
    case (sel) 0: mux_11650 = 1'h0; 1: mux_11650 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11651;
  wire [0:0] vin0_consume_en_11652;
  wire [0:0] vout_canPeek_11652;
  wire [7:0] vout_peek_11652;
  wire [0:0] v_11653;
  wire [0:0] v_11654;
  function [0:0] mux_11654(input [0:0] sel);
    case (sel) 0: mux_11654 = 1'h0; 1: mux_11654 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11655;
  function [0:0] mux_11655(input [0:0] sel);
    case (sel) 0: mux_11655 = 1'h0; 1: mux_11655 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11656;
  wire [0:0] v_11657;
  wire [0:0] v_11658;
  wire [0:0] v_11659;
  wire [0:0] v_11660;
  wire [0:0] v_11661;
  wire [0:0] v_11662;
  function [0:0] mux_11662(input [0:0] sel);
    case (sel) 0: mux_11662 = 1'h0; 1: mux_11662 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11663;
  function [0:0] mux_11663(input [0:0] sel);
    case (sel) 0: mux_11663 = 1'h0; 1: mux_11663 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11664;
  wire [0:0] v_11665;
  wire [0:0] v_11666;
  wire [0:0] v_11667;
  function [0:0] mux_11667(input [0:0] sel);
    case (sel) 0: mux_11667 = 1'h0; 1: mux_11667 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11668;
  function [0:0] mux_11668(input [0:0] sel);
    case (sel) 0: mux_11668 = 1'h0; 1: mux_11668 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11669;
  wire [0:0] v_11670;
  wire [0:0] v_11671;
  wire [0:0] v_11672;
  wire [0:0] v_11673;
  wire [0:0] v_11674;
  function [0:0] mux_11674(input [0:0] sel);
    case (sel) 0: mux_11674 = 1'h0; 1: mux_11674 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11675;
  wire [0:0] v_11676;
  wire [0:0] v_11677;
  wire [0:0] v_11678;
  wire [0:0] v_11679;
  function [0:0] mux_11679(input [0:0] sel);
    case (sel) 0: mux_11679 = 1'h0; 1: mux_11679 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11680;
  wire [0:0] v_11681;
  wire [0:0] v_11682;
  wire [0:0] v_11683;
  function [0:0] mux_11683(input [0:0] sel);
    case (sel) 0: mux_11683 = 1'h0; 1: mux_11683 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11684;
  function [0:0] mux_11684(input [0:0] sel);
    case (sel) 0: mux_11684 = 1'h0; 1: mux_11684 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_11685 = 1'h0;
  wire [0:0] v_11686;
  wire [0:0] v_11687;
  wire [0:0] act_11688;
  wire [0:0] v_11689;
  wire [0:0] v_11690;
  wire [0:0] v_11691;
  reg [0:0] v_11692 = 1'h0;
  wire [0:0] v_11693;
  wire [0:0] v_11694;
  wire [0:0] act_11695;
  wire [0:0] v_11696;
  wire [0:0] v_11697;
  wire [0:0] v_11698;
  wire [0:0] vin0_consume_en_11699;
  wire [0:0] vout_canPeek_11699;
  wire [7:0] vout_peek_11699;
  wire [0:0] v_11700;
  wire [0:0] v_11701;
  function [0:0] mux_11701(input [0:0] sel);
    case (sel) 0: mux_11701 = 1'h0; 1: mux_11701 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11702;
  wire [0:0] v_11703;
  wire [0:0] v_11704;
  wire [0:0] v_11705;
  wire [0:0] v_11706;
  function [0:0] mux_11706(input [0:0] sel);
    case (sel) 0: mux_11706 = 1'h0; 1: mux_11706 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11707;
  wire [0:0] vin0_consume_en_11708;
  wire [0:0] vout_canPeek_11708;
  wire [7:0] vout_peek_11708;
  wire [0:0] v_11709;
  wire [0:0] v_11710;
  function [0:0] mux_11710(input [0:0] sel);
    case (sel) 0: mux_11710 = 1'h0; 1: mux_11710 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11711;
  function [0:0] mux_11711(input [0:0] sel);
    case (sel) 0: mux_11711 = 1'h0; 1: mux_11711 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11712;
  wire [0:0] v_11713;
  wire [0:0] v_11714;
  wire [0:0] v_11715;
  wire [0:0] v_11716;
  wire [0:0] v_11717;
  wire [0:0] v_11718;
  function [0:0] mux_11718(input [0:0] sel);
    case (sel) 0: mux_11718 = 1'h0; 1: mux_11718 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11719;
  wire [0:0] v_11720;
  wire [0:0] v_11721;
  wire [0:0] v_11722;
  wire [0:0] v_11723;
  function [0:0] mux_11723(input [0:0] sel);
    case (sel) 0: mux_11723 = 1'h0; 1: mux_11723 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11724;
  wire [0:0] v_11725;
  wire [0:0] v_11726;
  wire [0:0] v_11727;
  function [0:0] mux_11727(input [0:0] sel);
    case (sel) 0: mux_11727 = 1'h0; 1: mux_11727 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11728;
  function [0:0] mux_11728(input [0:0] sel);
    case (sel) 0: mux_11728 = 1'h0; 1: mux_11728 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_11729 = 1'h0;
  wire [0:0] v_11730;
  wire [0:0] v_11731;
  wire [0:0] act_11732;
  wire [0:0] v_11733;
  wire [0:0] v_11734;
  wire [0:0] v_11735;
  wire [0:0] vin0_consume_en_11736;
  wire [0:0] vout_canPeek_11736;
  wire [7:0] vout_peek_11736;
  wire [0:0] v_11737;
  wire [0:0] v_11738;
  function [0:0] mux_11738(input [0:0] sel);
    case (sel) 0: mux_11738 = 1'h0; 1: mux_11738 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11739;
  wire [0:0] v_11740;
  wire [0:0] v_11741;
  wire [0:0] v_11742;
  wire [0:0] v_11743;
  function [0:0] mux_11743(input [0:0] sel);
    case (sel) 0: mux_11743 = 1'h0; 1: mux_11743 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11744;
  wire [0:0] vin0_consume_en_11745;
  wire [0:0] vout_canPeek_11745;
  wire [7:0] vout_peek_11745;
  wire [0:0] v_11746;
  wire [0:0] v_11747;
  function [0:0] mux_11747(input [0:0] sel);
    case (sel) 0: mux_11747 = 1'h0; 1: mux_11747 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11748;
  function [0:0] mux_11748(input [0:0] sel);
    case (sel) 0: mux_11748 = 1'h0; 1: mux_11748 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11749;
  wire [0:0] v_11750;
  wire [0:0] v_11751;
  wire [0:0] v_11752;
  wire [0:0] v_11753;
  wire [0:0] v_11754;
  wire [0:0] v_11755;
  function [0:0] mux_11755(input [0:0] sel);
    case (sel) 0: mux_11755 = 1'h0; 1: mux_11755 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11756;
  function [0:0] mux_11756(input [0:0] sel);
    case (sel) 0: mux_11756 = 1'h0; 1: mux_11756 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11757;
  wire [0:0] v_11758;
  wire [0:0] v_11759;
  wire [0:0] v_11760;
  function [0:0] mux_11760(input [0:0] sel);
    case (sel) 0: mux_11760 = 1'h0; 1: mux_11760 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11761;
  function [0:0] mux_11761(input [0:0] sel);
    case (sel) 0: mux_11761 = 1'h0; 1: mux_11761 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11762;
  wire [0:0] v_11763;
  wire [0:0] v_11764;
  wire [0:0] v_11765;
  wire [0:0] v_11766;
  wire [0:0] v_11767;
  function [0:0] mux_11767(input [0:0] sel);
    case (sel) 0: mux_11767 = 1'h0; 1: mux_11767 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11768;
  function [0:0] mux_11768(input [0:0] sel);
    case (sel) 0: mux_11768 = 1'h0; 1: mux_11768 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11769;
  wire [0:0] v_11770;
  wire [0:0] v_11771;
  wire [0:0] v_11772;
  function [0:0] mux_11772(input [0:0] sel);
    case (sel) 0: mux_11772 = 1'h0; 1: mux_11772 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11773;
  function [0:0] mux_11773(input [0:0] sel);
    case (sel) 0: mux_11773 = 1'h0; 1: mux_11773 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11774;
  wire [0:0] v_11775;
  wire [0:0] v_11776;
  wire [0:0] v_11777;
  wire [0:0] v_11778;
  wire [0:0] v_11779;
  function [0:0] mux_11779(input [0:0] sel);
    case (sel) 0: mux_11779 = 1'h0; 1: mux_11779 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11780;
  wire [0:0] v_11781;
  wire [0:0] v_11782;
  wire [0:0] v_11783;
  wire [0:0] v_11784;
  function [0:0] mux_11784(input [0:0] sel);
    case (sel) 0: mux_11784 = 1'h0; 1: mux_11784 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11785;
  wire [0:0] v_11786;
  wire [0:0] v_11787;
  wire [0:0] v_11788;
  function [0:0] mux_11788(input [0:0] sel);
    case (sel) 0: mux_11788 = 1'h0; 1: mux_11788 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11789;
  function [0:0] mux_11789(input [0:0] sel);
    case (sel) 0: mux_11789 = 1'h0; 1: mux_11789 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_11790 = 1'h0;
  wire [0:0] v_11791;
  wire [0:0] v_11792;
  wire [0:0] act_11793;
  wire [0:0] v_11794;
  wire [0:0] v_11795;
  wire [0:0] v_11796;
  reg [0:0] v_11797 = 1'h0;
  wire [0:0] v_11798;
  wire [0:0] v_11799;
  wire [0:0] act_11800;
  wire [0:0] v_11801;
  wire [0:0] v_11802;
  wire [0:0] v_11803;
  reg [0:0] v_11804 = 1'h0;
  wire [0:0] v_11805;
  wire [0:0] v_11806;
  wire [0:0] act_11807;
  wire [0:0] v_11808;
  wire [0:0] v_11809;
  wire [0:0] v_11810;
  wire [0:0] vin0_consume_en_11811;
  wire [0:0] vout_canPeek_11811;
  wire [7:0] vout_peek_11811;
  wire [0:0] v_11812;
  wire [0:0] v_11813;
  function [0:0] mux_11813(input [0:0] sel);
    case (sel) 0: mux_11813 = 1'h0; 1: mux_11813 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11814;
  wire [0:0] v_11815;
  wire [0:0] v_11816;
  wire [0:0] v_11817;
  wire [0:0] v_11818;
  function [0:0] mux_11818(input [0:0] sel);
    case (sel) 0: mux_11818 = 1'h0; 1: mux_11818 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11819;
  wire [0:0] vin0_consume_en_11820;
  wire [0:0] vout_canPeek_11820;
  wire [7:0] vout_peek_11820;
  wire [0:0] v_11821;
  wire [0:0] v_11822;
  function [0:0] mux_11822(input [0:0] sel);
    case (sel) 0: mux_11822 = 1'h0; 1: mux_11822 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11823;
  function [0:0] mux_11823(input [0:0] sel);
    case (sel) 0: mux_11823 = 1'h0; 1: mux_11823 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11824;
  wire [0:0] v_11825;
  wire [0:0] v_11826;
  wire [0:0] v_11827;
  wire [0:0] v_11828;
  wire [0:0] v_11829;
  wire [0:0] v_11830;
  function [0:0] mux_11830(input [0:0] sel);
    case (sel) 0: mux_11830 = 1'h0; 1: mux_11830 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11831;
  wire [0:0] v_11832;
  wire [0:0] v_11833;
  wire [0:0] v_11834;
  wire [0:0] v_11835;
  function [0:0] mux_11835(input [0:0] sel);
    case (sel) 0: mux_11835 = 1'h0; 1: mux_11835 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11836;
  wire [0:0] v_11837;
  wire [0:0] v_11838;
  wire [0:0] v_11839;
  function [0:0] mux_11839(input [0:0] sel);
    case (sel) 0: mux_11839 = 1'h0; 1: mux_11839 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11840;
  function [0:0] mux_11840(input [0:0] sel);
    case (sel) 0: mux_11840 = 1'h0; 1: mux_11840 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_11841 = 1'h0;
  wire [0:0] v_11842;
  wire [0:0] v_11843;
  wire [0:0] act_11844;
  wire [0:0] v_11845;
  wire [0:0] v_11846;
  wire [0:0] v_11847;
  wire [0:0] vin0_consume_en_11848;
  wire [0:0] vout_canPeek_11848;
  wire [7:0] vout_peek_11848;
  wire [0:0] v_11849;
  wire [0:0] v_11850;
  function [0:0] mux_11850(input [0:0] sel);
    case (sel) 0: mux_11850 = 1'h0; 1: mux_11850 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11851;
  wire [0:0] v_11852;
  wire [0:0] v_11853;
  wire [0:0] v_11854;
  wire [0:0] v_11855;
  function [0:0] mux_11855(input [0:0] sel);
    case (sel) 0: mux_11855 = 1'h0; 1: mux_11855 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11856;
  wire [0:0] vin0_consume_en_11857;
  wire [0:0] vout_canPeek_11857;
  wire [7:0] vout_peek_11857;
  wire [0:0] v_11858;
  wire [0:0] v_11859;
  function [0:0] mux_11859(input [0:0] sel);
    case (sel) 0: mux_11859 = 1'h0; 1: mux_11859 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11860;
  function [0:0] mux_11860(input [0:0] sel);
    case (sel) 0: mux_11860 = 1'h0; 1: mux_11860 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11861;
  wire [0:0] v_11862;
  wire [0:0] v_11863;
  wire [0:0] v_11864;
  wire [0:0] v_11865;
  wire [0:0] v_11866;
  wire [0:0] v_11867;
  function [0:0] mux_11867(input [0:0] sel);
    case (sel) 0: mux_11867 = 1'h0; 1: mux_11867 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11868;
  function [0:0] mux_11868(input [0:0] sel);
    case (sel) 0: mux_11868 = 1'h0; 1: mux_11868 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11869;
  wire [0:0] v_11870;
  wire [0:0] v_11871;
  wire [0:0] v_11872;
  function [0:0] mux_11872(input [0:0] sel);
    case (sel) 0: mux_11872 = 1'h0; 1: mux_11872 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11873;
  function [0:0] mux_11873(input [0:0] sel);
    case (sel) 0: mux_11873 = 1'h0; 1: mux_11873 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11874;
  wire [0:0] v_11875;
  wire [0:0] v_11876;
  wire [0:0] v_11877;
  wire [0:0] v_11878;
  wire [0:0] v_11879;
  function [0:0] mux_11879(input [0:0] sel);
    case (sel) 0: mux_11879 = 1'h0; 1: mux_11879 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11880;
  wire [0:0] v_11881;
  wire [0:0] v_11882;
  wire [0:0] v_11883;
  wire [0:0] v_11884;
  function [0:0] mux_11884(input [0:0] sel);
    case (sel) 0: mux_11884 = 1'h0; 1: mux_11884 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11885;
  wire [0:0] v_11886;
  wire [0:0] v_11887;
  wire [0:0] v_11888;
  function [0:0] mux_11888(input [0:0] sel);
    case (sel) 0: mux_11888 = 1'h0; 1: mux_11888 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11889;
  function [0:0] mux_11889(input [0:0] sel);
    case (sel) 0: mux_11889 = 1'h0; 1: mux_11889 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_11890 = 1'h0;
  wire [0:0] v_11891;
  wire [0:0] v_11892;
  wire [0:0] act_11893;
  wire [0:0] v_11894;
  wire [0:0] v_11895;
  wire [0:0] v_11896;
  reg [0:0] v_11897 = 1'h0;
  wire [0:0] v_11898;
  wire [0:0] v_11899;
  wire [0:0] act_11900;
  wire [0:0] v_11901;
  wire [0:0] v_11902;
  wire [0:0] v_11903;
  wire [0:0] vin0_consume_en_11904;
  wire [0:0] vout_canPeek_11904;
  wire [7:0] vout_peek_11904;
  wire [0:0] v_11905;
  wire [0:0] v_11906;
  function [0:0] mux_11906(input [0:0] sel);
    case (sel) 0: mux_11906 = 1'h0; 1: mux_11906 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11907;
  wire [0:0] v_11908;
  wire [0:0] v_11909;
  wire [0:0] v_11910;
  wire [0:0] v_11911;
  function [0:0] mux_11911(input [0:0] sel);
    case (sel) 0: mux_11911 = 1'h0; 1: mux_11911 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11912;
  wire [0:0] vin0_consume_en_11913;
  wire [0:0] vout_canPeek_11913;
  wire [7:0] vout_peek_11913;
  wire [0:0] v_11914;
  wire [0:0] v_11915;
  function [0:0] mux_11915(input [0:0] sel);
    case (sel) 0: mux_11915 = 1'h0; 1: mux_11915 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11916;
  function [0:0] mux_11916(input [0:0] sel);
    case (sel) 0: mux_11916 = 1'h0; 1: mux_11916 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11917;
  wire [0:0] v_11918;
  wire [0:0] v_11919;
  wire [0:0] v_11920;
  wire [0:0] v_11921;
  wire [0:0] v_11922;
  wire [0:0] v_11923;
  function [0:0] mux_11923(input [0:0] sel);
    case (sel) 0: mux_11923 = 1'h0; 1: mux_11923 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11924;
  wire [0:0] v_11925;
  wire [0:0] v_11926;
  wire [0:0] v_11927;
  wire [0:0] v_11928;
  function [0:0] mux_11928(input [0:0] sel);
    case (sel) 0: mux_11928 = 1'h0; 1: mux_11928 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11929;
  wire [0:0] v_11930;
  wire [0:0] v_11931;
  wire [0:0] v_11932;
  function [0:0] mux_11932(input [0:0] sel);
    case (sel) 0: mux_11932 = 1'h0; 1: mux_11932 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11933;
  function [0:0] mux_11933(input [0:0] sel);
    case (sel) 0: mux_11933 = 1'h0; 1: mux_11933 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_11934 = 1'h0;
  wire [0:0] v_11935;
  wire [0:0] v_11936;
  wire [0:0] act_11937;
  wire [0:0] v_11938;
  wire [0:0] v_11939;
  wire [0:0] v_11940;
  wire [0:0] vin0_consume_en_11941;
  wire [0:0] vout_canPeek_11941;
  wire [7:0] vout_peek_11941;
  wire [0:0] v_11942;
  wire [0:0] v_11943;
  function [0:0] mux_11943(input [0:0] sel);
    case (sel) 0: mux_11943 = 1'h0; 1: mux_11943 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11944;
  wire [0:0] v_11945;
  wire [0:0] v_11946;
  wire [0:0] v_11947;
  wire [0:0] v_11948;
  function [0:0] mux_11948(input [0:0] sel);
    case (sel) 0: mux_11948 = 1'h0; 1: mux_11948 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11949;
  wire [0:0] vin0_consume_en_11950;
  wire [0:0] vout_canPeek_11950;
  wire [7:0] vout_peek_11950;
  wire [0:0] v_11951;
  wire [0:0] v_11952;
  function [0:0] mux_11952(input [0:0] sel);
    case (sel) 0: mux_11952 = 1'h0; 1: mux_11952 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11953;
  function [0:0] mux_11953(input [0:0] sel);
    case (sel) 0: mux_11953 = 1'h0; 1: mux_11953 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11954;
  wire [0:0] v_11955;
  wire [0:0] v_11956;
  wire [0:0] v_11957;
  wire [0:0] v_11958;
  wire [0:0] v_11959;
  wire [0:0] v_11960;
  function [0:0] mux_11960(input [0:0] sel);
    case (sel) 0: mux_11960 = 1'h0; 1: mux_11960 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11961;
  function [0:0] mux_11961(input [0:0] sel);
    case (sel) 0: mux_11961 = 1'h0; 1: mux_11961 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11962;
  wire [0:0] v_11963;
  wire [0:0] v_11964;
  wire [0:0] v_11965;
  function [0:0] mux_11965(input [0:0] sel);
    case (sel) 0: mux_11965 = 1'h0; 1: mux_11965 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11966;
  function [0:0] mux_11966(input [0:0] sel);
    case (sel) 0: mux_11966 = 1'h0; 1: mux_11966 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11967;
  wire [0:0] v_11968;
  wire [0:0] v_11969;
  wire [0:0] v_11970;
  wire [0:0] v_11971;
  wire [0:0] v_11972;
  function [0:0] mux_11972(input [0:0] sel);
    case (sel) 0: mux_11972 = 1'h0; 1: mux_11972 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11973;
  function [0:0] mux_11973(input [0:0] sel);
    case (sel) 0: mux_11973 = 1'h0; 1: mux_11973 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11974;
  wire [0:0] v_11975;
  wire [0:0] v_11976;
  wire [0:0] v_11977;
  function [0:0] mux_11977(input [0:0] sel);
    case (sel) 0: mux_11977 = 1'h0; 1: mux_11977 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11978;
  function [0:0] mux_11978(input [0:0] sel);
    case (sel) 0: mux_11978 = 1'h0; 1: mux_11978 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11979;
  wire [0:0] v_11980;
  wire [0:0] v_11981;
  wire [0:0] v_11982;
  wire [0:0] v_11983;
  wire [0:0] v_11984;
  function [0:0] mux_11984(input [0:0] sel);
    case (sel) 0: mux_11984 = 1'h0; 1: mux_11984 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11985;
  function [0:0] mux_11985(input [0:0] sel);
    case (sel) 0: mux_11985 = 1'h0; 1: mux_11985 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11986;
  wire [0:0] v_11987;
  wire [0:0] v_11988;
  wire [0:0] v_11989;
  function [0:0] mux_11989(input [0:0] sel);
    case (sel) 0: mux_11989 = 1'h0; 1: mux_11989 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11990;
  function [0:0] mux_11990(input [0:0] sel);
    case (sel) 0: mux_11990 = 1'h0; 1: mux_11990 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_11991;
  wire [0:0] v_11992;
  wire [0:0] v_11993;
  wire [0:0] v_11994;
  wire [0:0] v_11995;
  wire [0:0] v_11996;
  function [0:0] mux_11996(input [0:0] sel);
    case (sel) 0: mux_11996 = 1'h0; 1: mux_11996 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_11997;
  wire [0:0] v_11998;
  wire [0:0] v_11999;
  wire [0:0] v_12000;
  wire [0:0] v_12001;
  function [0:0] mux_12001(input [0:0] sel);
    case (sel) 0: mux_12001 = 1'h0; 1: mux_12001 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12002;
  wire [0:0] v_12003;
  wire [0:0] v_12004;
  wire [0:0] v_12005;
  function [0:0] mux_12005(input [0:0] sel);
    case (sel) 0: mux_12005 = 1'h0; 1: mux_12005 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12006;
  function [0:0] mux_12006(input [0:0] sel);
    case (sel) 0: mux_12006 = 1'h0; 1: mux_12006 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_12007 = 1'h0;
  wire [0:0] v_12008;
  wire [0:0] v_12009;
  wire [0:0] act_12010;
  wire [0:0] v_12011;
  wire [0:0] v_12012;
  wire [0:0] v_12013;
  reg [0:0] v_12014 = 1'h0;
  wire [0:0] v_12015;
  wire [0:0] v_12016;
  wire [0:0] act_12017;
  wire [0:0] v_12018;
  wire [0:0] v_12019;
  wire [0:0] v_12020;
  reg [0:0] v_12021 = 1'h0;
  wire [0:0] v_12022;
  wire [0:0] v_12023;
  wire [0:0] act_12024;
  wire [0:0] v_12025;
  wire [0:0] v_12026;
  wire [0:0] v_12027;
  reg [0:0] v_12028 = 1'h0;
  wire [0:0] v_12029;
  wire [0:0] v_12030;
  wire [0:0] act_12031;
  wire [0:0] v_12032;
  wire [0:0] v_12033;
  wire [0:0] v_12034;
  wire [0:0] vin0_consume_en_12035;
  wire [0:0] vout_canPeek_12035;
  wire [7:0] vout_peek_12035;
  wire [0:0] v_12036;
  wire [0:0] v_12037;
  function [0:0] mux_12037(input [0:0] sel);
    case (sel) 0: mux_12037 = 1'h0; 1: mux_12037 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12038;
  wire [0:0] v_12039;
  wire [0:0] v_12040;
  wire [0:0] v_12041;
  wire [0:0] v_12042;
  function [0:0] mux_12042(input [0:0] sel);
    case (sel) 0: mux_12042 = 1'h0; 1: mux_12042 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12043;
  wire [0:0] vin0_consume_en_12044;
  wire [0:0] vout_canPeek_12044;
  wire [7:0] vout_peek_12044;
  wire [0:0] v_12045;
  wire [0:0] v_12046;
  function [0:0] mux_12046(input [0:0] sel);
    case (sel) 0: mux_12046 = 1'h0; 1: mux_12046 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12047;
  function [0:0] mux_12047(input [0:0] sel);
    case (sel) 0: mux_12047 = 1'h0; 1: mux_12047 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12048;
  wire [0:0] v_12049;
  wire [0:0] v_12050;
  wire [0:0] v_12051;
  wire [0:0] v_12052;
  wire [0:0] v_12053;
  wire [0:0] v_12054;
  function [0:0] mux_12054(input [0:0] sel);
    case (sel) 0: mux_12054 = 1'h0; 1: mux_12054 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12055;
  wire [0:0] v_12056;
  wire [0:0] v_12057;
  wire [0:0] v_12058;
  wire [0:0] v_12059;
  function [0:0] mux_12059(input [0:0] sel);
    case (sel) 0: mux_12059 = 1'h0; 1: mux_12059 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12060;
  wire [0:0] v_12061;
  wire [0:0] v_12062;
  wire [0:0] v_12063;
  function [0:0] mux_12063(input [0:0] sel);
    case (sel) 0: mux_12063 = 1'h0; 1: mux_12063 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12064;
  function [0:0] mux_12064(input [0:0] sel);
    case (sel) 0: mux_12064 = 1'h0; 1: mux_12064 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_12065 = 1'h0;
  wire [0:0] v_12066;
  wire [0:0] v_12067;
  wire [0:0] act_12068;
  wire [0:0] v_12069;
  wire [0:0] v_12070;
  wire [0:0] v_12071;
  wire [0:0] vin0_consume_en_12072;
  wire [0:0] vout_canPeek_12072;
  wire [7:0] vout_peek_12072;
  wire [0:0] v_12073;
  wire [0:0] v_12074;
  function [0:0] mux_12074(input [0:0] sel);
    case (sel) 0: mux_12074 = 1'h0; 1: mux_12074 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12075;
  wire [0:0] v_12076;
  wire [0:0] v_12077;
  wire [0:0] v_12078;
  wire [0:0] v_12079;
  function [0:0] mux_12079(input [0:0] sel);
    case (sel) 0: mux_12079 = 1'h0; 1: mux_12079 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12080;
  wire [0:0] vin0_consume_en_12081;
  wire [0:0] vout_canPeek_12081;
  wire [7:0] vout_peek_12081;
  wire [0:0] v_12082;
  wire [0:0] v_12083;
  function [0:0] mux_12083(input [0:0] sel);
    case (sel) 0: mux_12083 = 1'h0; 1: mux_12083 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12084;
  function [0:0] mux_12084(input [0:0] sel);
    case (sel) 0: mux_12084 = 1'h0; 1: mux_12084 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12085;
  wire [0:0] v_12086;
  wire [0:0] v_12087;
  wire [0:0] v_12088;
  wire [0:0] v_12089;
  wire [0:0] v_12090;
  wire [0:0] v_12091;
  function [0:0] mux_12091(input [0:0] sel);
    case (sel) 0: mux_12091 = 1'h0; 1: mux_12091 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12092;
  function [0:0] mux_12092(input [0:0] sel);
    case (sel) 0: mux_12092 = 1'h0; 1: mux_12092 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12093;
  wire [0:0] v_12094;
  wire [0:0] v_12095;
  wire [0:0] v_12096;
  function [0:0] mux_12096(input [0:0] sel);
    case (sel) 0: mux_12096 = 1'h0; 1: mux_12096 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12097;
  function [0:0] mux_12097(input [0:0] sel);
    case (sel) 0: mux_12097 = 1'h0; 1: mux_12097 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12098;
  wire [0:0] v_12099;
  wire [0:0] v_12100;
  wire [0:0] v_12101;
  wire [0:0] v_12102;
  wire [0:0] v_12103;
  function [0:0] mux_12103(input [0:0] sel);
    case (sel) 0: mux_12103 = 1'h0; 1: mux_12103 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12104;
  wire [0:0] v_12105;
  wire [0:0] v_12106;
  wire [0:0] v_12107;
  wire [0:0] v_12108;
  function [0:0] mux_12108(input [0:0] sel);
    case (sel) 0: mux_12108 = 1'h0; 1: mux_12108 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12109;
  wire [0:0] v_12110;
  wire [0:0] v_12111;
  wire [0:0] v_12112;
  function [0:0] mux_12112(input [0:0] sel);
    case (sel) 0: mux_12112 = 1'h0; 1: mux_12112 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12113;
  function [0:0] mux_12113(input [0:0] sel);
    case (sel) 0: mux_12113 = 1'h0; 1: mux_12113 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_12114 = 1'h0;
  wire [0:0] v_12115;
  wire [0:0] v_12116;
  wire [0:0] act_12117;
  wire [0:0] v_12118;
  wire [0:0] v_12119;
  wire [0:0] v_12120;
  reg [0:0] v_12121 = 1'h0;
  wire [0:0] v_12122;
  wire [0:0] v_12123;
  wire [0:0] act_12124;
  wire [0:0] v_12125;
  wire [0:0] v_12126;
  wire [0:0] v_12127;
  wire [0:0] vin0_consume_en_12128;
  wire [0:0] vout_canPeek_12128;
  wire [7:0] vout_peek_12128;
  wire [0:0] v_12129;
  wire [0:0] v_12130;
  function [0:0] mux_12130(input [0:0] sel);
    case (sel) 0: mux_12130 = 1'h0; 1: mux_12130 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12131;
  wire [0:0] v_12132;
  wire [0:0] v_12133;
  wire [0:0] v_12134;
  wire [0:0] v_12135;
  function [0:0] mux_12135(input [0:0] sel);
    case (sel) 0: mux_12135 = 1'h0; 1: mux_12135 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12136;
  wire [0:0] vin0_consume_en_12137;
  wire [0:0] vout_canPeek_12137;
  wire [7:0] vout_peek_12137;
  wire [0:0] v_12138;
  wire [0:0] v_12139;
  function [0:0] mux_12139(input [0:0] sel);
    case (sel) 0: mux_12139 = 1'h0; 1: mux_12139 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12140;
  function [0:0] mux_12140(input [0:0] sel);
    case (sel) 0: mux_12140 = 1'h0; 1: mux_12140 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12141;
  wire [0:0] v_12142;
  wire [0:0] v_12143;
  wire [0:0] v_12144;
  wire [0:0] v_12145;
  wire [0:0] v_12146;
  wire [0:0] v_12147;
  function [0:0] mux_12147(input [0:0] sel);
    case (sel) 0: mux_12147 = 1'h0; 1: mux_12147 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12148;
  wire [0:0] v_12149;
  wire [0:0] v_12150;
  wire [0:0] v_12151;
  wire [0:0] v_12152;
  function [0:0] mux_12152(input [0:0] sel);
    case (sel) 0: mux_12152 = 1'h0; 1: mux_12152 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12153;
  wire [0:0] v_12154;
  wire [0:0] v_12155;
  wire [0:0] v_12156;
  function [0:0] mux_12156(input [0:0] sel);
    case (sel) 0: mux_12156 = 1'h0; 1: mux_12156 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12157;
  function [0:0] mux_12157(input [0:0] sel);
    case (sel) 0: mux_12157 = 1'h0; 1: mux_12157 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_12158 = 1'h0;
  wire [0:0] v_12159;
  wire [0:0] v_12160;
  wire [0:0] act_12161;
  wire [0:0] v_12162;
  wire [0:0] v_12163;
  wire [0:0] v_12164;
  wire [0:0] vin0_consume_en_12165;
  wire [0:0] vout_canPeek_12165;
  wire [7:0] vout_peek_12165;
  wire [0:0] v_12166;
  wire [0:0] v_12167;
  function [0:0] mux_12167(input [0:0] sel);
    case (sel) 0: mux_12167 = 1'h0; 1: mux_12167 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12168;
  wire [0:0] v_12169;
  wire [0:0] v_12170;
  wire [0:0] v_12171;
  wire [0:0] v_12172;
  function [0:0] mux_12172(input [0:0] sel);
    case (sel) 0: mux_12172 = 1'h0; 1: mux_12172 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12173;
  wire [0:0] vin0_consume_en_12174;
  wire [0:0] vout_canPeek_12174;
  wire [7:0] vout_peek_12174;
  wire [0:0] v_12175;
  wire [0:0] v_12176;
  function [0:0] mux_12176(input [0:0] sel);
    case (sel) 0: mux_12176 = 1'h0; 1: mux_12176 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12177;
  function [0:0] mux_12177(input [0:0] sel);
    case (sel) 0: mux_12177 = 1'h0; 1: mux_12177 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12178;
  wire [0:0] v_12179;
  wire [0:0] v_12180;
  wire [0:0] v_12181;
  wire [0:0] v_12182;
  wire [0:0] v_12183;
  wire [0:0] v_12184;
  function [0:0] mux_12184(input [0:0] sel);
    case (sel) 0: mux_12184 = 1'h0; 1: mux_12184 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12185;
  function [0:0] mux_12185(input [0:0] sel);
    case (sel) 0: mux_12185 = 1'h0; 1: mux_12185 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12186;
  wire [0:0] v_12187;
  wire [0:0] v_12188;
  wire [0:0] v_12189;
  function [0:0] mux_12189(input [0:0] sel);
    case (sel) 0: mux_12189 = 1'h0; 1: mux_12189 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12190;
  function [0:0] mux_12190(input [0:0] sel);
    case (sel) 0: mux_12190 = 1'h0; 1: mux_12190 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12191;
  wire [0:0] v_12192;
  wire [0:0] v_12193;
  wire [0:0] v_12194;
  wire [0:0] v_12195;
  wire [0:0] v_12196;
  function [0:0] mux_12196(input [0:0] sel);
    case (sel) 0: mux_12196 = 1'h0; 1: mux_12196 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12197;
  function [0:0] mux_12197(input [0:0] sel);
    case (sel) 0: mux_12197 = 1'h0; 1: mux_12197 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12198;
  wire [0:0] v_12199;
  wire [0:0] v_12200;
  wire [0:0] v_12201;
  function [0:0] mux_12201(input [0:0] sel);
    case (sel) 0: mux_12201 = 1'h0; 1: mux_12201 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12202;
  function [0:0] mux_12202(input [0:0] sel);
    case (sel) 0: mux_12202 = 1'h0; 1: mux_12202 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12203;
  wire [0:0] v_12204;
  wire [0:0] v_12205;
  wire [0:0] v_12206;
  wire [0:0] v_12207;
  wire [0:0] v_12208;
  function [0:0] mux_12208(input [0:0] sel);
    case (sel) 0: mux_12208 = 1'h0; 1: mux_12208 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12209;
  wire [0:0] v_12210;
  wire [0:0] v_12211;
  wire [0:0] v_12212;
  wire [0:0] v_12213;
  function [0:0] mux_12213(input [0:0] sel);
    case (sel) 0: mux_12213 = 1'h0; 1: mux_12213 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12214;
  wire [0:0] v_12215;
  wire [0:0] v_12216;
  wire [0:0] v_12217;
  function [0:0] mux_12217(input [0:0] sel);
    case (sel) 0: mux_12217 = 1'h0; 1: mux_12217 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12218;
  function [0:0] mux_12218(input [0:0] sel);
    case (sel) 0: mux_12218 = 1'h0; 1: mux_12218 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_12219 = 1'h0;
  wire [0:0] v_12220;
  wire [0:0] v_12221;
  wire [0:0] act_12222;
  wire [0:0] v_12223;
  wire [0:0] v_12224;
  wire [0:0] v_12225;
  reg [0:0] v_12226 = 1'h0;
  wire [0:0] v_12227;
  wire [0:0] v_12228;
  wire [0:0] act_12229;
  wire [0:0] v_12230;
  wire [0:0] v_12231;
  wire [0:0] v_12232;
  reg [0:0] v_12233 = 1'h0;
  wire [0:0] v_12234;
  wire [0:0] v_12235;
  wire [0:0] act_12236;
  wire [0:0] v_12237;
  wire [0:0] v_12238;
  wire [0:0] v_12239;
  wire [0:0] vin0_consume_en_12240;
  wire [0:0] vout_canPeek_12240;
  wire [7:0] vout_peek_12240;
  wire [0:0] v_12241;
  wire [0:0] v_12242;
  function [0:0] mux_12242(input [0:0] sel);
    case (sel) 0: mux_12242 = 1'h0; 1: mux_12242 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12243;
  wire [0:0] v_12244;
  wire [0:0] v_12245;
  wire [0:0] v_12246;
  wire [0:0] v_12247;
  function [0:0] mux_12247(input [0:0] sel);
    case (sel) 0: mux_12247 = 1'h0; 1: mux_12247 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12248;
  wire [0:0] vin0_consume_en_12249;
  wire [0:0] vout_canPeek_12249;
  wire [7:0] vout_peek_12249;
  wire [0:0] v_12250;
  wire [0:0] v_12251;
  function [0:0] mux_12251(input [0:0] sel);
    case (sel) 0: mux_12251 = 1'h0; 1: mux_12251 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12252;
  function [0:0] mux_12252(input [0:0] sel);
    case (sel) 0: mux_12252 = 1'h0; 1: mux_12252 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12253;
  wire [0:0] v_12254;
  wire [0:0] v_12255;
  wire [0:0] v_12256;
  wire [0:0] v_12257;
  wire [0:0] v_12258;
  wire [0:0] v_12259;
  function [0:0] mux_12259(input [0:0] sel);
    case (sel) 0: mux_12259 = 1'h0; 1: mux_12259 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12260;
  wire [0:0] v_12261;
  wire [0:0] v_12262;
  wire [0:0] v_12263;
  wire [0:0] v_12264;
  function [0:0] mux_12264(input [0:0] sel);
    case (sel) 0: mux_12264 = 1'h0; 1: mux_12264 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12265;
  wire [0:0] v_12266;
  wire [0:0] v_12267;
  wire [0:0] v_12268;
  function [0:0] mux_12268(input [0:0] sel);
    case (sel) 0: mux_12268 = 1'h0; 1: mux_12268 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12269;
  function [0:0] mux_12269(input [0:0] sel);
    case (sel) 0: mux_12269 = 1'h0; 1: mux_12269 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_12270 = 1'h0;
  wire [0:0] v_12271;
  wire [0:0] v_12272;
  wire [0:0] act_12273;
  wire [0:0] v_12274;
  wire [0:0] v_12275;
  wire [0:0] v_12276;
  wire [0:0] vin0_consume_en_12277;
  wire [0:0] vout_canPeek_12277;
  wire [7:0] vout_peek_12277;
  wire [0:0] v_12278;
  wire [0:0] v_12279;
  function [0:0] mux_12279(input [0:0] sel);
    case (sel) 0: mux_12279 = 1'h0; 1: mux_12279 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12280;
  wire [0:0] v_12281;
  wire [0:0] v_12282;
  wire [0:0] v_12283;
  wire [0:0] v_12284;
  function [0:0] mux_12284(input [0:0] sel);
    case (sel) 0: mux_12284 = 1'h0; 1: mux_12284 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12285;
  wire [0:0] vin0_consume_en_12286;
  wire [0:0] vout_canPeek_12286;
  wire [7:0] vout_peek_12286;
  wire [0:0] v_12287;
  wire [0:0] v_12288;
  function [0:0] mux_12288(input [0:0] sel);
    case (sel) 0: mux_12288 = 1'h0; 1: mux_12288 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12289;
  function [0:0] mux_12289(input [0:0] sel);
    case (sel) 0: mux_12289 = 1'h0; 1: mux_12289 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12290;
  wire [0:0] v_12291;
  wire [0:0] v_12292;
  wire [0:0] v_12293;
  wire [0:0] v_12294;
  wire [0:0] v_12295;
  wire [0:0] v_12296;
  function [0:0] mux_12296(input [0:0] sel);
    case (sel) 0: mux_12296 = 1'h0; 1: mux_12296 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12297;
  function [0:0] mux_12297(input [0:0] sel);
    case (sel) 0: mux_12297 = 1'h0; 1: mux_12297 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12298;
  wire [0:0] v_12299;
  wire [0:0] v_12300;
  wire [0:0] v_12301;
  function [0:0] mux_12301(input [0:0] sel);
    case (sel) 0: mux_12301 = 1'h0; 1: mux_12301 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12302;
  function [0:0] mux_12302(input [0:0] sel);
    case (sel) 0: mux_12302 = 1'h0; 1: mux_12302 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12303;
  wire [0:0] v_12304;
  wire [0:0] v_12305;
  wire [0:0] v_12306;
  wire [0:0] v_12307;
  wire [0:0] v_12308;
  function [0:0] mux_12308(input [0:0] sel);
    case (sel) 0: mux_12308 = 1'h0; 1: mux_12308 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12309;
  wire [0:0] v_12310;
  wire [0:0] v_12311;
  wire [0:0] v_12312;
  wire [0:0] v_12313;
  function [0:0] mux_12313(input [0:0] sel);
    case (sel) 0: mux_12313 = 1'h0; 1: mux_12313 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12314;
  wire [0:0] v_12315;
  wire [0:0] v_12316;
  wire [0:0] v_12317;
  function [0:0] mux_12317(input [0:0] sel);
    case (sel) 0: mux_12317 = 1'h0; 1: mux_12317 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12318;
  function [0:0] mux_12318(input [0:0] sel);
    case (sel) 0: mux_12318 = 1'h0; 1: mux_12318 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_12319 = 1'h0;
  wire [0:0] v_12320;
  wire [0:0] v_12321;
  wire [0:0] act_12322;
  wire [0:0] v_12323;
  wire [0:0] v_12324;
  wire [0:0] v_12325;
  reg [0:0] v_12326 = 1'h0;
  wire [0:0] v_12327;
  wire [0:0] v_12328;
  wire [0:0] act_12329;
  wire [0:0] v_12330;
  wire [0:0] v_12331;
  wire [0:0] v_12332;
  wire [0:0] vin0_consume_en_12333;
  wire [0:0] vout_canPeek_12333;
  wire [7:0] vout_peek_12333;
  wire [0:0] v_12334;
  wire [0:0] v_12335;
  function [0:0] mux_12335(input [0:0] sel);
    case (sel) 0: mux_12335 = 1'h0; 1: mux_12335 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12336;
  wire [0:0] v_12337;
  wire [0:0] v_12338;
  wire [0:0] v_12339;
  wire [0:0] v_12340;
  function [0:0] mux_12340(input [0:0] sel);
    case (sel) 0: mux_12340 = 1'h0; 1: mux_12340 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12341;
  wire [0:0] vin0_consume_en_12342;
  wire [0:0] vout_canPeek_12342;
  wire [7:0] vout_peek_12342;
  wire [0:0] v_12343;
  wire [0:0] v_12344;
  function [0:0] mux_12344(input [0:0] sel);
    case (sel) 0: mux_12344 = 1'h0; 1: mux_12344 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12345;
  function [0:0] mux_12345(input [0:0] sel);
    case (sel) 0: mux_12345 = 1'h0; 1: mux_12345 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12346;
  wire [0:0] v_12347;
  wire [0:0] v_12348;
  wire [0:0] v_12349;
  wire [0:0] v_12350;
  wire [0:0] v_12351;
  wire [0:0] v_12352;
  function [0:0] mux_12352(input [0:0] sel);
    case (sel) 0: mux_12352 = 1'h0; 1: mux_12352 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12353;
  wire [0:0] v_12354;
  wire [0:0] v_12355;
  wire [0:0] v_12356;
  wire [0:0] v_12357;
  function [0:0] mux_12357(input [0:0] sel);
    case (sel) 0: mux_12357 = 1'h0; 1: mux_12357 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12358;
  wire [0:0] v_12359;
  wire [0:0] v_12360;
  wire [0:0] v_12361;
  function [0:0] mux_12361(input [0:0] sel);
    case (sel) 0: mux_12361 = 1'h0; 1: mux_12361 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12362;
  function [0:0] mux_12362(input [0:0] sel);
    case (sel) 0: mux_12362 = 1'h0; 1: mux_12362 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_12363 = 1'h0;
  wire [0:0] v_12364;
  wire [0:0] v_12365;
  wire [0:0] act_12366;
  wire [0:0] v_12367;
  wire [0:0] v_12368;
  wire [0:0] v_12369;
  wire [0:0] vin0_consume_en_12370;
  wire [0:0] vout_canPeek_12370;
  wire [7:0] vout_peek_12370;
  wire [0:0] v_12371;
  wire [0:0] v_12372;
  function [0:0] mux_12372(input [0:0] sel);
    case (sel) 0: mux_12372 = 1'h0; 1: mux_12372 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12373;
  wire [0:0] v_12374;
  wire [0:0] v_12375;
  wire [0:0] v_12376;
  wire [0:0] v_12377;
  function [0:0] mux_12377(input [0:0] sel);
    case (sel) 0: mux_12377 = 1'h0; 1: mux_12377 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12378;
  wire [0:0] vin0_consume_en_12379;
  wire [0:0] vout_canPeek_12379;
  wire [7:0] vout_peek_12379;
  wire [0:0] v_12380;
  wire [0:0] v_12381;
  function [0:0] mux_12381(input [0:0] sel);
    case (sel) 0: mux_12381 = 1'h0; 1: mux_12381 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12382;
  function [0:0] mux_12382(input [0:0] sel);
    case (sel) 0: mux_12382 = 1'h0; 1: mux_12382 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12383;
  wire [0:0] v_12384;
  wire [0:0] v_12385;
  wire [0:0] v_12386;
  wire [0:0] v_12387;
  wire [0:0] v_12388;
  wire [0:0] v_12389;
  function [0:0] mux_12389(input [0:0] sel);
    case (sel) 0: mux_12389 = 1'h0; 1: mux_12389 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12390;
  function [0:0] mux_12390(input [0:0] sel);
    case (sel) 0: mux_12390 = 1'h0; 1: mux_12390 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12391;
  wire [0:0] v_12392;
  wire [0:0] v_12393;
  wire [0:0] v_12394;
  function [0:0] mux_12394(input [0:0] sel);
    case (sel) 0: mux_12394 = 1'h0; 1: mux_12394 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12395;
  function [0:0] mux_12395(input [0:0] sel);
    case (sel) 0: mux_12395 = 1'h0; 1: mux_12395 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12396;
  wire [0:0] v_12397;
  wire [0:0] v_12398;
  wire [0:0] v_12399;
  wire [0:0] v_12400;
  wire [0:0] v_12401;
  function [0:0] mux_12401(input [0:0] sel);
    case (sel) 0: mux_12401 = 1'h0; 1: mux_12401 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12402;
  function [0:0] mux_12402(input [0:0] sel);
    case (sel) 0: mux_12402 = 1'h0; 1: mux_12402 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12403;
  wire [0:0] v_12404;
  wire [0:0] v_12405;
  wire [0:0] v_12406;
  function [0:0] mux_12406(input [0:0] sel);
    case (sel) 0: mux_12406 = 1'h0; 1: mux_12406 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12407;
  function [0:0] mux_12407(input [0:0] sel);
    case (sel) 0: mux_12407 = 1'h0; 1: mux_12407 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12408;
  wire [0:0] v_12409;
  wire [0:0] v_12410;
  wire [0:0] v_12411;
  wire [0:0] v_12412;
  wire [0:0] v_12413;
  function [0:0] mux_12413(input [0:0] sel);
    case (sel) 0: mux_12413 = 1'h0; 1: mux_12413 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12414;
  function [0:0] mux_12414(input [0:0] sel);
    case (sel) 0: mux_12414 = 1'h0; 1: mux_12414 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12415;
  wire [0:0] v_12416;
  wire [0:0] v_12417;
  wire [0:0] v_12418;
  function [0:0] mux_12418(input [0:0] sel);
    case (sel) 0: mux_12418 = 1'h0; 1: mux_12418 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12419;
  function [0:0] mux_12419(input [0:0] sel);
    case (sel) 0: mux_12419 = 1'h0; 1: mux_12419 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12420;
  wire [0:0] v_12421;
  wire [0:0] v_12422;
  wire [0:0] v_12423;
  wire [0:0] v_12424;
  wire [0:0] v_12425;
  function [0:0] mux_12425(input [0:0] sel);
    case (sel) 0: mux_12425 = 1'h0; 1: mux_12425 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12426;
  function [0:0] mux_12426(input [0:0] sel);
    case (sel) 0: mux_12426 = 1'h0; 1: mux_12426 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12427;
  wire [0:0] v_12428;
  wire [0:0] v_12429;
  wire [0:0] v_12430;
  function [0:0] mux_12430(input [0:0] sel);
    case (sel) 0: mux_12430 = 1'h0; 1: mux_12430 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12431;
  function [0:0] mux_12431(input [0:0] sel);
    case (sel) 0: mux_12431 = 1'h0; 1: mux_12431 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12432;
  wire [0:0] v_12433;
  wire [0:0] v_12434;
  wire [0:0] v_12435;
  wire [0:0] v_12436;
  wire [0:0] v_12437;
  function [0:0] mux_12437(input [0:0] sel);
    case (sel) 0: mux_12437 = 1'h0; 1: mux_12437 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12438;
  wire [0:0] v_12439;
  wire [0:0] v_12440;
  wire [0:0] v_12441;
  wire [0:0] v_12442;
  function [0:0] mux_12442(input [0:0] sel);
    case (sel) 0: mux_12442 = 1'h0; 1: mux_12442 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12443;
  wire [0:0] v_12444;
  wire [0:0] v_12445;
  wire [0:0] v_12446;
  function [0:0] mux_12446(input [0:0] sel);
    case (sel) 0: mux_12446 = 1'h0; 1: mux_12446 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12447;
  function [0:0] mux_12447(input [0:0] sel);
    case (sel) 0: mux_12447 = 1'h0; 1: mux_12447 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_12448 = 1'h0;
  wire [0:0] v_12449;
  wire [0:0] v_12450;
  wire [0:0] act_12451;
  wire [0:0] v_12452;
  wire [0:0] v_12453;
  wire [0:0] v_12454;
  reg [0:0] v_12455 = 1'h0;
  wire [0:0] v_12456;
  wire [0:0] v_12457;
  wire [0:0] act_12458;
  wire [0:0] v_12459;
  wire [0:0] v_12460;
  wire [0:0] v_12461;
  reg [0:0] v_12462 = 1'h0;
  wire [0:0] v_12463;
  wire [0:0] v_12464;
  wire [0:0] act_12465;
  wire [0:0] v_12466;
  wire [0:0] v_12467;
  wire [0:0] v_12468;
  reg [0:0] v_12469 = 1'h0;
  wire [0:0] v_12470;
  wire [0:0] v_12471;
  wire [0:0] act_12472;
  wire [0:0] v_12473;
  wire [0:0] v_12474;
  wire [0:0] v_12475;
  reg [0:0] v_12476 = 1'h0;
  wire [0:0] v_12477;
  wire [0:0] v_12478;
  wire [0:0] act_12479;
  wire [0:0] v_12480;
  wire [0:0] v_12481;
  wire [0:0] v_12482;
  wire [0:0] vin0_consume_en_12483;
  wire [0:0] vout_canPeek_12483;
  wire [7:0] vout_peek_12483;
  wire [0:0] v_12484;
  wire [0:0] v_12485;
  function [0:0] mux_12485(input [0:0] sel);
    case (sel) 0: mux_12485 = 1'h0; 1: mux_12485 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12486;
  wire [0:0] v_12487;
  wire [0:0] v_12488;
  wire [0:0] v_12489;
  wire [0:0] v_12490;
  function [0:0] mux_12490(input [0:0] sel);
    case (sel) 0: mux_12490 = 1'h0; 1: mux_12490 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12491;
  wire [0:0] vin0_consume_en_12492;
  wire [0:0] vout_canPeek_12492;
  wire [7:0] vout_peek_12492;
  wire [0:0] v_12493;
  wire [0:0] v_12494;
  function [0:0] mux_12494(input [0:0] sel);
    case (sel) 0: mux_12494 = 1'h0; 1: mux_12494 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12495;
  function [0:0] mux_12495(input [0:0] sel);
    case (sel) 0: mux_12495 = 1'h0; 1: mux_12495 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12496;
  wire [0:0] v_12497;
  wire [0:0] v_12498;
  wire [0:0] v_12499;
  wire [0:0] v_12500;
  wire [0:0] v_12501;
  wire [0:0] v_12502;
  function [0:0] mux_12502(input [0:0] sel);
    case (sel) 0: mux_12502 = 1'h0; 1: mux_12502 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12503;
  wire [0:0] v_12504;
  wire [0:0] v_12505;
  wire [0:0] v_12506;
  wire [0:0] v_12507;
  function [0:0] mux_12507(input [0:0] sel);
    case (sel) 0: mux_12507 = 1'h0; 1: mux_12507 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12508;
  wire [0:0] v_12509;
  wire [0:0] v_12510;
  wire [0:0] v_12511;
  function [0:0] mux_12511(input [0:0] sel);
    case (sel) 0: mux_12511 = 1'h0; 1: mux_12511 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12512;
  function [0:0] mux_12512(input [0:0] sel);
    case (sel) 0: mux_12512 = 1'h0; 1: mux_12512 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_12513 = 1'h0;
  wire [0:0] v_12514;
  wire [0:0] v_12515;
  wire [0:0] act_12516;
  wire [0:0] v_12517;
  wire [0:0] v_12518;
  wire [0:0] v_12519;
  wire [0:0] vin0_consume_en_12520;
  wire [0:0] vout_canPeek_12520;
  wire [7:0] vout_peek_12520;
  wire [0:0] v_12521;
  wire [0:0] v_12522;
  function [0:0] mux_12522(input [0:0] sel);
    case (sel) 0: mux_12522 = 1'h0; 1: mux_12522 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12523;
  wire [0:0] v_12524;
  wire [0:0] v_12525;
  wire [0:0] v_12526;
  wire [0:0] v_12527;
  function [0:0] mux_12527(input [0:0] sel);
    case (sel) 0: mux_12527 = 1'h0; 1: mux_12527 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12528;
  wire [0:0] vin0_consume_en_12529;
  wire [0:0] vout_canPeek_12529;
  wire [7:0] vout_peek_12529;
  wire [0:0] v_12530;
  wire [0:0] v_12531;
  function [0:0] mux_12531(input [0:0] sel);
    case (sel) 0: mux_12531 = 1'h0; 1: mux_12531 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12532;
  function [0:0] mux_12532(input [0:0] sel);
    case (sel) 0: mux_12532 = 1'h0; 1: mux_12532 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12533;
  wire [0:0] v_12534;
  wire [0:0] v_12535;
  wire [0:0] v_12536;
  wire [0:0] v_12537;
  wire [0:0] v_12538;
  wire [0:0] v_12539;
  function [0:0] mux_12539(input [0:0] sel);
    case (sel) 0: mux_12539 = 1'h0; 1: mux_12539 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12540;
  function [0:0] mux_12540(input [0:0] sel);
    case (sel) 0: mux_12540 = 1'h0; 1: mux_12540 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12541;
  wire [0:0] v_12542;
  wire [0:0] v_12543;
  wire [0:0] v_12544;
  function [0:0] mux_12544(input [0:0] sel);
    case (sel) 0: mux_12544 = 1'h0; 1: mux_12544 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12545;
  function [0:0] mux_12545(input [0:0] sel);
    case (sel) 0: mux_12545 = 1'h0; 1: mux_12545 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12546;
  wire [0:0] v_12547;
  wire [0:0] v_12548;
  wire [0:0] v_12549;
  wire [0:0] v_12550;
  wire [0:0] v_12551;
  function [0:0] mux_12551(input [0:0] sel);
    case (sel) 0: mux_12551 = 1'h0; 1: mux_12551 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12552;
  wire [0:0] v_12553;
  wire [0:0] v_12554;
  wire [0:0] v_12555;
  wire [0:0] v_12556;
  function [0:0] mux_12556(input [0:0] sel);
    case (sel) 0: mux_12556 = 1'h0; 1: mux_12556 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12557;
  wire [0:0] v_12558;
  wire [0:0] v_12559;
  wire [0:0] v_12560;
  function [0:0] mux_12560(input [0:0] sel);
    case (sel) 0: mux_12560 = 1'h0; 1: mux_12560 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12561;
  function [0:0] mux_12561(input [0:0] sel);
    case (sel) 0: mux_12561 = 1'h0; 1: mux_12561 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_12562 = 1'h0;
  wire [0:0] v_12563;
  wire [0:0] v_12564;
  wire [0:0] act_12565;
  wire [0:0] v_12566;
  wire [0:0] v_12567;
  wire [0:0] v_12568;
  reg [0:0] v_12569 = 1'h0;
  wire [0:0] v_12570;
  wire [0:0] v_12571;
  wire [0:0] act_12572;
  wire [0:0] v_12573;
  wire [0:0] v_12574;
  wire [0:0] v_12575;
  wire [0:0] vin0_consume_en_12576;
  wire [0:0] vout_canPeek_12576;
  wire [7:0] vout_peek_12576;
  wire [0:0] v_12577;
  wire [0:0] v_12578;
  function [0:0] mux_12578(input [0:0] sel);
    case (sel) 0: mux_12578 = 1'h0; 1: mux_12578 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12579;
  wire [0:0] v_12580;
  wire [0:0] v_12581;
  wire [0:0] v_12582;
  wire [0:0] v_12583;
  function [0:0] mux_12583(input [0:0] sel);
    case (sel) 0: mux_12583 = 1'h0; 1: mux_12583 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12584;
  wire [0:0] vin0_consume_en_12585;
  wire [0:0] vout_canPeek_12585;
  wire [7:0] vout_peek_12585;
  wire [0:0] v_12586;
  wire [0:0] v_12587;
  function [0:0] mux_12587(input [0:0] sel);
    case (sel) 0: mux_12587 = 1'h0; 1: mux_12587 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12588;
  function [0:0] mux_12588(input [0:0] sel);
    case (sel) 0: mux_12588 = 1'h0; 1: mux_12588 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12589;
  wire [0:0] v_12590;
  wire [0:0] v_12591;
  wire [0:0] v_12592;
  wire [0:0] v_12593;
  wire [0:0] v_12594;
  wire [0:0] v_12595;
  function [0:0] mux_12595(input [0:0] sel);
    case (sel) 0: mux_12595 = 1'h0; 1: mux_12595 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12596;
  wire [0:0] v_12597;
  wire [0:0] v_12598;
  wire [0:0] v_12599;
  wire [0:0] v_12600;
  function [0:0] mux_12600(input [0:0] sel);
    case (sel) 0: mux_12600 = 1'h0; 1: mux_12600 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12601;
  wire [0:0] v_12602;
  wire [0:0] v_12603;
  wire [0:0] v_12604;
  function [0:0] mux_12604(input [0:0] sel);
    case (sel) 0: mux_12604 = 1'h0; 1: mux_12604 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12605;
  function [0:0] mux_12605(input [0:0] sel);
    case (sel) 0: mux_12605 = 1'h0; 1: mux_12605 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_12606 = 1'h0;
  wire [0:0] v_12607;
  wire [0:0] v_12608;
  wire [0:0] act_12609;
  wire [0:0] v_12610;
  wire [0:0] v_12611;
  wire [0:0] v_12612;
  wire [0:0] vin0_consume_en_12613;
  wire [0:0] vout_canPeek_12613;
  wire [7:0] vout_peek_12613;
  wire [0:0] v_12614;
  wire [0:0] v_12615;
  function [0:0] mux_12615(input [0:0] sel);
    case (sel) 0: mux_12615 = 1'h0; 1: mux_12615 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12616;
  wire [0:0] v_12617;
  wire [0:0] v_12618;
  wire [0:0] v_12619;
  wire [0:0] v_12620;
  function [0:0] mux_12620(input [0:0] sel);
    case (sel) 0: mux_12620 = 1'h0; 1: mux_12620 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12621;
  wire [0:0] vin0_consume_en_12622;
  wire [0:0] vout_canPeek_12622;
  wire [7:0] vout_peek_12622;
  wire [0:0] v_12623;
  wire [0:0] v_12624;
  function [0:0] mux_12624(input [0:0] sel);
    case (sel) 0: mux_12624 = 1'h0; 1: mux_12624 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12625;
  function [0:0] mux_12625(input [0:0] sel);
    case (sel) 0: mux_12625 = 1'h0; 1: mux_12625 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12626;
  wire [0:0] v_12627;
  wire [0:0] v_12628;
  wire [0:0] v_12629;
  wire [0:0] v_12630;
  wire [0:0] v_12631;
  wire [0:0] v_12632;
  function [0:0] mux_12632(input [0:0] sel);
    case (sel) 0: mux_12632 = 1'h0; 1: mux_12632 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12633;
  function [0:0] mux_12633(input [0:0] sel);
    case (sel) 0: mux_12633 = 1'h0; 1: mux_12633 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12634;
  wire [0:0] v_12635;
  wire [0:0] v_12636;
  wire [0:0] v_12637;
  function [0:0] mux_12637(input [0:0] sel);
    case (sel) 0: mux_12637 = 1'h0; 1: mux_12637 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12638;
  function [0:0] mux_12638(input [0:0] sel);
    case (sel) 0: mux_12638 = 1'h0; 1: mux_12638 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12639;
  wire [0:0] v_12640;
  wire [0:0] v_12641;
  wire [0:0] v_12642;
  wire [0:0] v_12643;
  wire [0:0] v_12644;
  function [0:0] mux_12644(input [0:0] sel);
    case (sel) 0: mux_12644 = 1'h0; 1: mux_12644 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12645;
  function [0:0] mux_12645(input [0:0] sel);
    case (sel) 0: mux_12645 = 1'h0; 1: mux_12645 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12646;
  wire [0:0] v_12647;
  wire [0:0] v_12648;
  wire [0:0] v_12649;
  function [0:0] mux_12649(input [0:0] sel);
    case (sel) 0: mux_12649 = 1'h0; 1: mux_12649 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12650;
  function [0:0] mux_12650(input [0:0] sel);
    case (sel) 0: mux_12650 = 1'h0; 1: mux_12650 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12651;
  wire [0:0] v_12652;
  wire [0:0] v_12653;
  wire [0:0] v_12654;
  wire [0:0] v_12655;
  wire [0:0] v_12656;
  function [0:0] mux_12656(input [0:0] sel);
    case (sel) 0: mux_12656 = 1'h0; 1: mux_12656 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12657;
  wire [0:0] v_12658;
  wire [0:0] v_12659;
  wire [0:0] v_12660;
  wire [0:0] v_12661;
  function [0:0] mux_12661(input [0:0] sel);
    case (sel) 0: mux_12661 = 1'h0; 1: mux_12661 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12662;
  wire [0:0] v_12663;
  wire [0:0] v_12664;
  wire [0:0] v_12665;
  function [0:0] mux_12665(input [0:0] sel);
    case (sel) 0: mux_12665 = 1'h0; 1: mux_12665 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12666;
  function [0:0] mux_12666(input [0:0] sel);
    case (sel) 0: mux_12666 = 1'h0; 1: mux_12666 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_12667 = 1'h0;
  wire [0:0] v_12668;
  wire [0:0] v_12669;
  wire [0:0] act_12670;
  wire [0:0] v_12671;
  wire [0:0] v_12672;
  wire [0:0] v_12673;
  reg [0:0] v_12674 = 1'h0;
  wire [0:0] v_12675;
  wire [0:0] v_12676;
  wire [0:0] act_12677;
  wire [0:0] v_12678;
  wire [0:0] v_12679;
  wire [0:0] v_12680;
  reg [0:0] v_12681 = 1'h0;
  wire [0:0] v_12682;
  wire [0:0] v_12683;
  wire [0:0] act_12684;
  wire [0:0] v_12685;
  wire [0:0] v_12686;
  wire [0:0] v_12687;
  wire [0:0] vin0_consume_en_12688;
  wire [0:0] vout_canPeek_12688;
  wire [7:0] vout_peek_12688;
  wire [0:0] v_12689;
  wire [0:0] v_12690;
  function [0:0] mux_12690(input [0:0] sel);
    case (sel) 0: mux_12690 = 1'h0; 1: mux_12690 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12691;
  wire [0:0] v_12692;
  wire [0:0] v_12693;
  wire [0:0] v_12694;
  wire [0:0] v_12695;
  function [0:0] mux_12695(input [0:0] sel);
    case (sel) 0: mux_12695 = 1'h0; 1: mux_12695 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12696;
  wire [0:0] vin0_consume_en_12697;
  wire [0:0] vout_canPeek_12697;
  wire [7:0] vout_peek_12697;
  wire [0:0] v_12698;
  wire [0:0] v_12699;
  function [0:0] mux_12699(input [0:0] sel);
    case (sel) 0: mux_12699 = 1'h0; 1: mux_12699 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12700;
  function [0:0] mux_12700(input [0:0] sel);
    case (sel) 0: mux_12700 = 1'h0; 1: mux_12700 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12701;
  wire [0:0] v_12702;
  wire [0:0] v_12703;
  wire [0:0] v_12704;
  wire [0:0] v_12705;
  wire [0:0] v_12706;
  wire [0:0] v_12707;
  function [0:0] mux_12707(input [0:0] sel);
    case (sel) 0: mux_12707 = 1'h0; 1: mux_12707 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12708;
  wire [0:0] v_12709;
  wire [0:0] v_12710;
  wire [0:0] v_12711;
  wire [0:0] v_12712;
  function [0:0] mux_12712(input [0:0] sel);
    case (sel) 0: mux_12712 = 1'h0; 1: mux_12712 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12713;
  wire [0:0] v_12714;
  wire [0:0] v_12715;
  wire [0:0] v_12716;
  function [0:0] mux_12716(input [0:0] sel);
    case (sel) 0: mux_12716 = 1'h0; 1: mux_12716 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12717;
  function [0:0] mux_12717(input [0:0] sel);
    case (sel) 0: mux_12717 = 1'h0; 1: mux_12717 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_12718 = 1'h0;
  wire [0:0] v_12719;
  wire [0:0] v_12720;
  wire [0:0] act_12721;
  wire [0:0] v_12722;
  wire [0:0] v_12723;
  wire [0:0] v_12724;
  wire [0:0] vin0_consume_en_12725;
  wire [0:0] vout_canPeek_12725;
  wire [7:0] vout_peek_12725;
  wire [0:0] v_12726;
  wire [0:0] v_12727;
  function [0:0] mux_12727(input [0:0] sel);
    case (sel) 0: mux_12727 = 1'h0; 1: mux_12727 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12728;
  wire [0:0] v_12729;
  wire [0:0] v_12730;
  wire [0:0] v_12731;
  wire [0:0] v_12732;
  function [0:0] mux_12732(input [0:0] sel);
    case (sel) 0: mux_12732 = 1'h0; 1: mux_12732 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12733;
  wire [0:0] vin0_consume_en_12734;
  wire [0:0] vout_canPeek_12734;
  wire [7:0] vout_peek_12734;
  wire [0:0] v_12735;
  wire [0:0] v_12736;
  function [0:0] mux_12736(input [0:0] sel);
    case (sel) 0: mux_12736 = 1'h0; 1: mux_12736 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12737;
  function [0:0] mux_12737(input [0:0] sel);
    case (sel) 0: mux_12737 = 1'h0; 1: mux_12737 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12738;
  wire [0:0] v_12739;
  wire [0:0] v_12740;
  wire [0:0] v_12741;
  wire [0:0] v_12742;
  wire [0:0] v_12743;
  wire [0:0] v_12744;
  function [0:0] mux_12744(input [0:0] sel);
    case (sel) 0: mux_12744 = 1'h0; 1: mux_12744 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12745;
  function [0:0] mux_12745(input [0:0] sel);
    case (sel) 0: mux_12745 = 1'h0; 1: mux_12745 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12746;
  wire [0:0] v_12747;
  wire [0:0] v_12748;
  wire [0:0] v_12749;
  function [0:0] mux_12749(input [0:0] sel);
    case (sel) 0: mux_12749 = 1'h0; 1: mux_12749 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12750;
  function [0:0] mux_12750(input [0:0] sel);
    case (sel) 0: mux_12750 = 1'h0; 1: mux_12750 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12751;
  wire [0:0] v_12752;
  wire [0:0] v_12753;
  wire [0:0] v_12754;
  wire [0:0] v_12755;
  wire [0:0] v_12756;
  function [0:0] mux_12756(input [0:0] sel);
    case (sel) 0: mux_12756 = 1'h0; 1: mux_12756 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12757;
  wire [0:0] v_12758;
  wire [0:0] v_12759;
  wire [0:0] v_12760;
  wire [0:0] v_12761;
  function [0:0] mux_12761(input [0:0] sel);
    case (sel) 0: mux_12761 = 1'h0; 1: mux_12761 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12762;
  wire [0:0] v_12763;
  wire [0:0] v_12764;
  wire [0:0] v_12765;
  function [0:0] mux_12765(input [0:0] sel);
    case (sel) 0: mux_12765 = 1'h0; 1: mux_12765 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12766;
  function [0:0] mux_12766(input [0:0] sel);
    case (sel) 0: mux_12766 = 1'h0; 1: mux_12766 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_12767 = 1'h0;
  wire [0:0] v_12768;
  wire [0:0] v_12769;
  wire [0:0] act_12770;
  wire [0:0] v_12771;
  wire [0:0] v_12772;
  wire [0:0] v_12773;
  reg [0:0] v_12774 = 1'h0;
  wire [0:0] v_12775;
  wire [0:0] v_12776;
  wire [0:0] act_12777;
  wire [0:0] v_12778;
  wire [0:0] v_12779;
  wire [0:0] v_12780;
  wire [0:0] vin0_consume_en_12781;
  wire [0:0] vout_canPeek_12781;
  wire [7:0] vout_peek_12781;
  wire [0:0] v_12782;
  wire [0:0] v_12783;
  function [0:0] mux_12783(input [0:0] sel);
    case (sel) 0: mux_12783 = 1'h0; 1: mux_12783 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12784;
  wire [0:0] v_12785;
  wire [0:0] v_12786;
  wire [0:0] v_12787;
  wire [0:0] v_12788;
  function [0:0] mux_12788(input [0:0] sel);
    case (sel) 0: mux_12788 = 1'h0; 1: mux_12788 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12789;
  wire [0:0] vin0_consume_en_12790;
  wire [0:0] vout_canPeek_12790;
  wire [7:0] vout_peek_12790;
  wire [0:0] v_12791;
  wire [0:0] v_12792;
  function [0:0] mux_12792(input [0:0] sel);
    case (sel) 0: mux_12792 = 1'h0; 1: mux_12792 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12793;
  function [0:0] mux_12793(input [0:0] sel);
    case (sel) 0: mux_12793 = 1'h0; 1: mux_12793 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12794;
  wire [0:0] v_12795;
  wire [0:0] v_12796;
  wire [0:0] v_12797;
  wire [0:0] v_12798;
  wire [0:0] v_12799;
  wire [0:0] v_12800;
  function [0:0] mux_12800(input [0:0] sel);
    case (sel) 0: mux_12800 = 1'h0; 1: mux_12800 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12801;
  wire [0:0] v_12802;
  wire [0:0] v_12803;
  wire [0:0] v_12804;
  wire [0:0] v_12805;
  function [0:0] mux_12805(input [0:0] sel);
    case (sel) 0: mux_12805 = 1'h0; 1: mux_12805 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12806;
  wire [0:0] v_12807;
  wire [0:0] v_12808;
  wire [0:0] v_12809;
  function [0:0] mux_12809(input [0:0] sel);
    case (sel) 0: mux_12809 = 1'h0; 1: mux_12809 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12810;
  function [0:0] mux_12810(input [0:0] sel);
    case (sel) 0: mux_12810 = 1'h0; 1: mux_12810 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_12811 = 1'h0;
  wire [0:0] v_12812;
  wire [0:0] v_12813;
  wire [0:0] act_12814;
  wire [0:0] v_12815;
  wire [0:0] v_12816;
  wire [0:0] v_12817;
  wire [0:0] vin0_consume_en_12818;
  wire [0:0] vout_canPeek_12818;
  wire [7:0] vout_peek_12818;
  wire [0:0] v_12819;
  wire [0:0] v_12820;
  function [0:0] mux_12820(input [0:0] sel);
    case (sel) 0: mux_12820 = 1'h0; 1: mux_12820 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12821;
  wire [0:0] v_12822;
  wire [0:0] v_12823;
  wire [0:0] v_12824;
  wire [0:0] v_12825;
  function [0:0] mux_12825(input [0:0] sel);
    case (sel) 0: mux_12825 = 1'h0; 1: mux_12825 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12826;
  wire [0:0] vin0_consume_en_12827;
  wire [0:0] vout_canPeek_12827;
  wire [7:0] vout_peek_12827;
  wire [0:0] v_12828;
  wire [0:0] v_12829;
  function [0:0] mux_12829(input [0:0] sel);
    case (sel) 0: mux_12829 = 1'h0; 1: mux_12829 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12830;
  function [0:0] mux_12830(input [0:0] sel);
    case (sel) 0: mux_12830 = 1'h0; 1: mux_12830 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12831;
  wire [0:0] v_12832;
  wire [0:0] v_12833;
  wire [0:0] v_12834;
  wire [0:0] v_12835;
  wire [0:0] v_12836;
  wire [0:0] v_12837;
  function [0:0] mux_12837(input [0:0] sel);
    case (sel) 0: mux_12837 = 1'h0; 1: mux_12837 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12838;
  function [0:0] mux_12838(input [0:0] sel);
    case (sel) 0: mux_12838 = 1'h0; 1: mux_12838 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12839;
  wire [0:0] v_12840;
  wire [0:0] v_12841;
  wire [0:0] v_12842;
  function [0:0] mux_12842(input [0:0] sel);
    case (sel) 0: mux_12842 = 1'h0; 1: mux_12842 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12843;
  function [0:0] mux_12843(input [0:0] sel);
    case (sel) 0: mux_12843 = 1'h0; 1: mux_12843 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12844;
  wire [0:0] v_12845;
  wire [0:0] v_12846;
  wire [0:0] v_12847;
  wire [0:0] v_12848;
  wire [0:0] v_12849;
  function [0:0] mux_12849(input [0:0] sel);
    case (sel) 0: mux_12849 = 1'h0; 1: mux_12849 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12850;
  function [0:0] mux_12850(input [0:0] sel);
    case (sel) 0: mux_12850 = 1'h0; 1: mux_12850 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12851;
  wire [0:0] v_12852;
  wire [0:0] v_12853;
  wire [0:0] v_12854;
  function [0:0] mux_12854(input [0:0] sel);
    case (sel) 0: mux_12854 = 1'h0; 1: mux_12854 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12855;
  function [0:0] mux_12855(input [0:0] sel);
    case (sel) 0: mux_12855 = 1'h0; 1: mux_12855 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12856;
  wire [0:0] v_12857;
  wire [0:0] v_12858;
  wire [0:0] v_12859;
  wire [0:0] v_12860;
  wire [0:0] v_12861;
  function [0:0] mux_12861(input [0:0] sel);
    case (sel) 0: mux_12861 = 1'h0; 1: mux_12861 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12862;
  function [0:0] mux_12862(input [0:0] sel);
    case (sel) 0: mux_12862 = 1'h0; 1: mux_12862 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12863;
  wire [0:0] v_12864;
  wire [0:0] v_12865;
  wire [0:0] v_12866;
  function [0:0] mux_12866(input [0:0] sel);
    case (sel) 0: mux_12866 = 1'h0; 1: mux_12866 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12867;
  function [0:0] mux_12867(input [0:0] sel);
    case (sel) 0: mux_12867 = 1'h0; 1: mux_12867 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12868;
  wire [0:0] v_12869;
  wire [0:0] v_12870;
  wire [0:0] v_12871;
  wire [0:0] v_12872;
  wire [0:0] v_12873;
  function [0:0] mux_12873(input [0:0] sel);
    case (sel) 0: mux_12873 = 1'h0; 1: mux_12873 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12874;
  wire [0:0] v_12875;
  wire [0:0] v_12876;
  wire [0:0] v_12877;
  wire [0:0] v_12878;
  function [0:0] mux_12878(input [0:0] sel);
    case (sel) 0: mux_12878 = 1'h0; 1: mux_12878 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12879;
  wire [0:0] v_12880;
  wire [0:0] v_12881;
  wire [0:0] v_12882;
  function [0:0] mux_12882(input [0:0] sel);
    case (sel) 0: mux_12882 = 1'h0; 1: mux_12882 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12883;
  function [0:0] mux_12883(input [0:0] sel);
    case (sel) 0: mux_12883 = 1'h0; 1: mux_12883 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_12884 = 1'h0;
  wire [0:0] v_12885;
  wire [0:0] v_12886;
  wire [0:0] act_12887;
  wire [0:0] v_12888;
  wire [0:0] v_12889;
  wire [0:0] v_12890;
  reg [0:0] v_12891 = 1'h0;
  wire [0:0] v_12892;
  wire [0:0] v_12893;
  wire [0:0] act_12894;
  wire [0:0] v_12895;
  wire [0:0] v_12896;
  wire [0:0] v_12897;
  reg [0:0] v_12898 = 1'h0;
  wire [0:0] v_12899;
  wire [0:0] v_12900;
  wire [0:0] act_12901;
  wire [0:0] v_12902;
  wire [0:0] v_12903;
  wire [0:0] v_12904;
  reg [0:0] v_12905 = 1'h0;
  wire [0:0] v_12906;
  wire [0:0] v_12907;
  wire [0:0] act_12908;
  wire [0:0] v_12909;
  wire [0:0] v_12910;
  wire [0:0] v_12911;
  wire [0:0] vin0_consume_en_12912;
  wire [0:0] vout_canPeek_12912;
  wire [7:0] vout_peek_12912;
  wire [0:0] v_12913;
  wire [0:0] v_12914;
  function [0:0] mux_12914(input [0:0] sel);
    case (sel) 0: mux_12914 = 1'h0; 1: mux_12914 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12915;
  wire [0:0] v_12916;
  wire [0:0] v_12917;
  wire [0:0] v_12918;
  wire [0:0] v_12919;
  function [0:0] mux_12919(input [0:0] sel);
    case (sel) 0: mux_12919 = 1'h0; 1: mux_12919 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12920;
  wire [0:0] vin0_consume_en_12921;
  wire [0:0] vout_canPeek_12921;
  wire [7:0] vout_peek_12921;
  wire [0:0] v_12922;
  wire [0:0] v_12923;
  function [0:0] mux_12923(input [0:0] sel);
    case (sel) 0: mux_12923 = 1'h0; 1: mux_12923 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12924;
  function [0:0] mux_12924(input [0:0] sel);
    case (sel) 0: mux_12924 = 1'h0; 1: mux_12924 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12925;
  wire [0:0] v_12926;
  wire [0:0] v_12927;
  wire [0:0] v_12928;
  wire [0:0] v_12929;
  wire [0:0] v_12930;
  wire [0:0] v_12931;
  function [0:0] mux_12931(input [0:0] sel);
    case (sel) 0: mux_12931 = 1'h0; 1: mux_12931 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12932;
  wire [0:0] v_12933;
  wire [0:0] v_12934;
  wire [0:0] v_12935;
  wire [0:0] v_12936;
  function [0:0] mux_12936(input [0:0] sel);
    case (sel) 0: mux_12936 = 1'h0; 1: mux_12936 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12937;
  wire [0:0] v_12938;
  wire [0:0] v_12939;
  wire [0:0] v_12940;
  function [0:0] mux_12940(input [0:0] sel);
    case (sel) 0: mux_12940 = 1'h0; 1: mux_12940 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12941;
  function [0:0] mux_12941(input [0:0] sel);
    case (sel) 0: mux_12941 = 1'h0; 1: mux_12941 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_12942 = 1'h0;
  wire [0:0] v_12943;
  wire [0:0] v_12944;
  wire [0:0] act_12945;
  wire [0:0] v_12946;
  wire [0:0] v_12947;
  wire [0:0] v_12948;
  wire [0:0] vin0_consume_en_12949;
  wire [0:0] vout_canPeek_12949;
  wire [7:0] vout_peek_12949;
  wire [0:0] v_12950;
  wire [0:0] v_12951;
  function [0:0] mux_12951(input [0:0] sel);
    case (sel) 0: mux_12951 = 1'h0; 1: mux_12951 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12952;
  wire [0:0] v_12953;
  wire [0:0] v_12954;
  wire [0:0] v_12955;
  wire [0:0] v_12956;
  function [0:0] mux_12956(input [0:0] sel);
    case (sel) 0: mux_12956 = 1'h0; 1: mux_12956 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12957;
  wire [0:0] vin0_consume_en_12958;
  wire [0:0] vout_canPeek_12958;
  wire [7:0] vout_peek_12958;
  wire [0:0] v_12959;
  wire [0:0] v_12960;
  function [0:0] mux_12960(input [0:0] sel);
    case (sel) 0: mux_12960 = 1'h0; 1: mux_12960 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12961;
  function [0:0] mux_12961(input [0:0] sel);
    case (sel) 0: mux_12961 = 1'h0; 1: mux_12961 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12962;
  wire [0:0] v_12963;
  wire [0:0] v_12964;
  wire [0:0] v_12965;
  wire [0:0] v_12966;
  wire [0:0] v_12967;
  wire [0:0] v_12968;
  function [0:0] mux_12968(input [0:0] sel);
    case (sel) 0: mux_12968 = 1'h0; 1: mux_12968 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12969;
  function [0:0] mux_12969(input [0:0] sel);
    case (sel) 0: mux_12969 = 1'h0; 1: mux_12969 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12970;
  wire [0:0] v_12971;
  wire [0:0] v_12972;
  wire [0:0] v_12973;
  function [0:0] mux_12973(input [0:0] sel);
    case (sel) 0: mux_12973 = 1'h0; 1: mux_12973 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12974;
  function [0:0] mux_12974(input [0:0] sel);
    case (sel) 0: mux_12974 = 1'h0; 1: mux_12974 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12975;
  wire [0:0] v_12976;
  wire [0:0] v_12977;
  wire [0:0] v_12978;
  wire [0:0] v_12979;
  wire [0:0] v_12980;
  function [0:0] mux_12980(input [0:0] sel);
    case (sel) 0: mux_12980 = 1'h0; 1: mux_12980 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12981;
  wire [0:0] v_12982;
  wire [0:0] v_12983;
  wire [0:0] v_12984;
  wire [0:0] v_12985;
  function [0:0] mux_12985(input [0:0] sel);
    case (sel) 0: mux_12985 = 1'h0; 1: mux_12985 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_12986;
  wire [0:0] v_12987;
  wire [0:0] v_12988;
  wire [0:0] v_12989;
  function [0:0] mux_12989(input [0:0] sel);
    case (sel) 0: mux_12989 = 1'h0; 1: mux_12989 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_12990;
  function [0:0] mux_12990(input [0:0] sel);
    case (sel) 0: mux_12990 = 1'h0; 1: mux_12990 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_12991 = 1'h0;
  wire [0:0] v_12992;
  wire [0:0] v_12993;
  wire [0:0] act_12994;
  wire [0:0] v_12995;
  wire [0:0] v_12996;
  wire [0:0] v_12997;
  reg [0:0] v_12998 = 1'h0;
  wire [0:0] v_12999;
  wire [0:0] v_13000;
  wire [0:0] act_13001;
  wire [0:0] v_13002;
  wire [0:0] v_13003;
  wire [0:0] v_13004;
  wire [0:0] vin0_consume_en_13005;
  wire [0:0] vout_canPeek_13005;
  wire [7:0] vout_peek_13005;
  wire [0:0] v_13006;
  wire [0:0] v_13007;
  function [0:0] mux_13007(input [0:0] sel);
    case (sel) 0: mux_13007 = 1'h0; 1: mux_13007 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13008;
  wire [0:0] v_13009;
  wire [0:0] v_13010;
  wire [0:0] v_13011;
  wire [0:0] v_13012;
  function [0:0] mux_13012(input [0:0] sel);
    case (sel) 0: mux_13012 = 1'h0; 1: mux_13012 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13013;
  wire [0:0] vin0_consume_en_13014;
  wire [0:0] vout_canPeek_13014;
  wire [7:0] vout_peek_13014;
  wire [0:0] v_13015;
  wire [0:0] v_13016;
  function [0:0] mux_13016(input [0:0] sel);
    case (sel) 0: mux_13016 = 1'h0; 1: mux_13016 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13017;
  function [0:0] mux_13017(input [0:0] sel);
    case (sel) 0: mux_13017 = 1'h0; 1: mux_13017 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13018;
  wire [0:0] v_13019;
  wire [0:0] v_13020;
  wire [0:0] v_13021;
  wire [0:0] v_13022;
  wire [0:0] v_13023;
  wire [0:0] v_13024;
  function [0:0] mux_13024(input [0:0] sel);
    case (sel) 0: mux_13024 = 1'h0; 1: mux_13024 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13025;
  wire [0:0] v_13026;
  wire [0:0] v_13027;
  wire [0:0] v_13028;
  wire [0:0] v_13029;
  function [0:0] mux_13029(input [0:0] sel);
    case (sel) 0: mux_13029 = 1'h0; 1: mux_13029 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13030;
  wire [0:0] v_13031;
  wire [0:0] v_13032;
  wire [0:0] v_13033;
  function [0:0] mux_13033(input [0:0] sel);
    case (sel) 0: mux_13033 = 1'h0; 1: mux_13033 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13034;
  function [0:0] mux_13034(input [0:0] sel);
    case (sel) 0: mux_13034 = 1'h0; 1: mux_13034 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_13035 = 1'h0;
  wire [0:0] v_13036;
  wire [0:0] v_13037;
  wire [0:0] act_13038;
  wire [0:0] v_13039;
  wire [0:0] v_13040;
  wire [0:0] v_13041;
  wire [0:0] vin0_consume_en_13042;
  wire [0:0] vout_canPeek_13042;
  wire [7:0] vout_peek_13042;
  wire [0:0] v_13043;
  wire [0:0] v_13044;
  function [0:0] mux_13044(input [0:0] sel);
    case (sel) 0: mux_13044 = 1'h0; 1: mux_13044 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13045;
  wire [0:0] v_13046;
  wire [0:0] v_13047;
  wire [0:0] v_13048;
  wire [0:0] v_13049;
  function [0:0] mux_13049(input [0:0] sel);
    case (sel) 0: mux_13049 = 1'h0; 1: mux_13049 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13050;
  wire [0:0] vin0_consume_en_13051;
  wire [0:0] vout_canPeek_13051;
  wire [7:0] vout_peek_13051;
  wire [0:0] v_13052;
  wire [0:0] v_13053;
  function [0:0] mux_13053(input [0:0] sel);
    case (sel) 0: mux_13053 = 1'h0; 1: mux_13053 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13054;
  function [0:0] mux_13054(input [0:0] sel);
    case (sel) 0: mux_13054 = 1'h0; 1: mux_13054 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13055;
  wire [0:0] v_13056;
  wire [0:0] v_13057;
  wire [0:0] v_13058;
  wire [0:0] v_13059;
  wire [0:0] v_13060;
  wire [0:0] v_13061;
  function [0:0] mux_13061(input [0:0] sel);
    case (sel) 0: mux_13061 = 1'h0; 1: mux_13061 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13062;
  function [0:0] mux_13062(input [0:0] sel);
    case (sel) 0: mux_13062 = 1'h0; 1: mux_13062 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13063;
  wire [0:0] v_13064;
  wire [0:0] v_13065;
  wire [0:0] v_13066;
  function [0:0] mux_13066(input [0:0] sel);
    case (sel) 0: mux_13066 = 1'h0; 1: mux_13066 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13067;
  function [0:0] mux_13067(input [0:0] sel);
    case (sel) 0: mux_13067 = 1'h0; 1: mux_13067 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13068;
  wire [0:0] v_13069;
  wire [0:0] v_13070;
  wire [0:0] v_13071;
  wire [0:0] v_13072;
  wire [0:0] v_13073;
  function [0:0] mux_13073(input [0:0] sel);
    case (sel) 0: mux_13073 = 1'h0; 1: mux_13073 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13074;
  function [0:0] mux_13074(input [0:0] sel);
    case (sel) 0: mux_13074 = 1'h0; 1: mux_13074 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13075;
  wire [0:0] v_13076;
  wire [0:0] v_13077;
  wire [0:0] v_13078;
  function [0:0] mux_13078(input [0:0] sel);
    case (sel) 0: mux_13078 = 1'h0; 1: mux_13078 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13079;
  function [0:0] mux_13079(input [0:0] sel);
    case (sel) 0: mux_13079 = 1'h0; 1: mux_13079 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13080;
  wire [0:0] v_13081;
  wire [0:0] v_13082;
  wire [0:0] v_13083;
  wire [0:0] v_13084;
  wire [0:0] v_13085;
  function [0:0] mux_13085(input [0:0] sel);
    case (sel) 0: mux_13085 = 1'h0; 1: mux_13085 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13086;
  wire [0:0] v_13087;
  wire [0:0] v_13088;
  wire [0:0] v_13089;
  wire [0:0] v_13090;
  function [0:0] mux_13090(input [0:0] sel);
    case (sel) 0: mux_13090 = 1'h0; 1: mux_13090 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13091;
  wire [0:0] v_13092;
  wire [0:0] v_13093;
  wire [0:0] v_13094;
  function [0:0] mux_13094(input [0:0] sel);
    case (sel) 0: mux_13094 = 1'h0; 1: mux_13094 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13095;
  function [0:0] mux_13095(input [0:0] sel);
    case (sel) 0: mux_13095 = 1'h0; 1: mux_13095 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_13096 = 1'h0;
  wire [0:0] v_13097;
  wire [0:0] v_13098;
  wire [0:0] act_13099;
  wire [0:0] v_13100;
  wire [0:0] v_13101;
  wire [0:0] v_13102;
  reg [0:0] v_13103 = 1'h0;
  wire [0:0] v_13104;
  wire [0:0] v_13105;
  wire [0:0] act_13106;
  wire [0:0] v_13107;
  wire [0:0] v_13108;
  wire [0:0] v_13109;
  reg [0:0] v_13110 = 1'h0;
  wire [0:0] v_13111;
  wire [0:0] v_13112;
  wire [0:0] act_13113;
  wire [0:0] v_13114;
  wire [0:0] v_13115;
  wire [0:0] v_13116;
  wire [0:0] vin0_consume_en_13117;
  wire [0:0] vout_canPeek_13117;
  wire [7:0] vout_peek_13117;
  wire [0:0] v_13118;
  wire [0:0] v_13119;
  function [0:0] mux_13119(input [0:0] sel);
    case (sel) 0: mux_13119 = 1'h0; 1: mux_13119 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13120;
  wire [0:0] v_13121;
  wire [0:0] v_13122;
  wire [0:0] v_13123;
  wire [0:0] v_13124;
  function [0:0] mux_13124(input [0:0] sel);
    case (sel) 0: mux_13124 = 1'h0; 1: mux_13124 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13125;
  wire [0:0] vin0_consume_en_13126;
  wire [0:0] vout_canPeek_13126;
  wire [7:0] vout_peek_13126;
  wire [0:0] v_13127;
  wire [0:0] v_13128;
  function [0:0] mux_13128(input [0:0] sel);
    case (sel) 0: mux_13128 = 1'h0; 1: mux_13128 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13129;
  function [0:0] mux_13129(input [0:0] sel);
    case (sel) 0: mux_13129 = 1'h0; 1: mux_13129 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13130;
  wire [0:0] v_13131;
  wire [0:0] v_13132;
  wire [0:0] v_13133;
  wire [0:0] v_13134;
  wire [0:0] v_13135;
  wire [0:0] v_13136;
  function [0:0] mux_13136(input [0:0] sel);
    case (sel) 0: mux_13136 = 1'h0; 1: mux_13136 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13137;
  wire [0:0] v_13138;
  wire [0:0] v_13139;
  wire [0:0] v_13140;
  wire [0:0] v_13141;
  function [0:0] mux_13141(input [0:0] sel);
    case (sel) 0: mux_13141 = 1'h0; 1: mux_13141 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13142;
  wire [0:0] v_13143;
  wire [0:0] v_13144;
  wire [0:0] v_13145;
  function [0:0] mux_13145(input [0:0] sel);
    case (sel) 0: mux_13145 = 1'h0; 1: mux_13145 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13146;
  function [0:0] mux_13146(input [0:0] sel);
    case (sel) 0: mux_13146 = 1'h0; 1: mux_13146 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_13147 = 1'h0;
  wire [0:0] v_13148;
  wire [0:0] v_13149;
  wire [0:0] act_13150;
  wire [0:0] v_13151;
  wire [0:0] v_13152;
  wire [0:0] v_13153;
  wire [0:0] vin0_consume_en_13154;
  wire [0:0] vout_canPeek_13154;
  wire [7:0] vout_peek_13154;
  wire [0:0] v_13155;
  wire [0:0] v_13156;
  function [0:0] mux_13156(input [0:0] sel);
    case (sel) 0: mux_13156 = 1'h0; 1: mux_13156 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13157;
  wire [0:0] v_13158;
  wire [0:0] v_13159;
  wire [0:0] v_13160;
  wire [0:0] v_13161;
  function [0:0] mux_13161(input [0:0] sel);
    case (sel) 0: mux_13161 = 1'h0; 1: mux_13161 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13162;
  wire [0:0] vin0_consume_en_13163;
  wire [0:0] vout_canPeek_13163;
  wire [7:0] vout_peek_13163;
  wire [0:0] v_13164;
  wire [0:0] v_13165;
  function [0:0] mux_13165(input [0:0] sel);
    case (sel) 0: mux_13165 = 1'h0; 1: mux_13165 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13166;
  function [0:0] mux_13166(input [0:0] sel);
    case (sel) 0: mux_13166 = 1'h0; 1: mux_13166 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13167;
  wire [0:0] v_13168;
  wire [0:0] v_13169;
  wire [0:0] v_13170;
  wire [0:0] v_13171;
  wire [0:0] v_13172;
  wire [0:0] v_13173;
  function [0:0] mux_13173(input [0:0] sel);
    case (sel) 0: mux_13173 = 1'h0; 1: mux_13173 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13174;
  function [0:0] mux_13174(input [0:0] sel);
    case (sel) 0: mux_13174 = 1'h0; 1: mux_13174 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13175;
  wire [0:0] v_13176;
  wire [0:0] v_13177;
  wire [0:0] v_13178;
  function [0:0] mux_13178(input [0:0] sel);
    case (sel) 0: mux_13178 = 1'h0; 1: mux_13178 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13179;
  function [0:0] mux_13179(input [0:0] sel);
    case (sel) 0: mux_13179 = 1'h0; 1: mux_13179 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13180;
  wire [0:0] v_13181;
  wire [0:0] v_13182;
  wire [0:0] v_13183;
  wire [0:0] v_13184;
  wire [0:0] v_13185;
  function [0:0] mux_13185(input [0:0] sel);
    case (sel) 0: mux_13185 = 1'h0; 1: mux_13185 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13186;
  wire [0:0] v_13187;
  wire [0:0] v_13188;
  wire [0:0] v_13189;
  wire [0:0] v_13190;
  function [0:0] mux_13190(input [0:0] sel);
    case (sel) 0: mux_13190 = 1'h0; 1: mux_13190 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13191;
  wire [0:0] v_13192;
  wire [0:0] v_13193;
  wire [0:0] v_13194;
  function [0:0] mux_13194(input [0:0] sel);
    case (sel) 0: mux_13194 = 1'h0; 1: mux_13194 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13195;
  function [0:0] mux_13195(input [0:0] sel);
    case (sel) 0: mux_13195 = 1'h0; 1: mux_13195 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_13196 = 1'h0;
  wire [0:0] v_13197;
  wire [0:0] v_13198;
  wire [0:0] act_13199;
  wire [0:0] v_13200;
  wire [0:0] v_13201;
  wire [0:0] v_13202;
  reg [0:0] v_13203 = 1'h0;
  wire [0:0] v_13204;
  wire [0:0] v_13205;
  wire [0:0] act_13206;
  wire [0:0] v_13207;
  wire [0:0] v_13208;
  wire [0:0] v_13209;
  wire [0:0] vin0_consume_en_13210;
  wire [0:0] vout_canPeek_13210;
  wire [7:0] vout_peek_13210;
  wire [0:0] v_13211;
  wire [0:0] v_13212;
  function [0:0] mux_13212(input [0:0] sel);
    case (sel) 0: mux_13212 = 1'h0; 1: mux_13212 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13213;
  wire [0:0] v_13214;
  wire [0:0] v_13215;
  wire [0:0] v_13216;
  wire [0:0] v_13217;
  function [0:0] mux_13217(input [0:0] sel);
    case (sel) 0: mux_13217 = 1'h0; 1: mux_13217 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13218;
  wire [0:0] vin0_consume_en_13219;
  wire [0:0] vout_canPeek_13219;
  wire [7:0] vout_peek_13219;
  wire [0:0] v_13220;
  wire [0:0] v_13221;
  function [0:0] mux_13221(input [0:0] sel);
    case (sel) 0: mux_13221 = 1'h0; 1: mux_13221 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13222;
  function [0:0] mux_13222(input [0:0] sel);
    case (sel) 0: mux_13222 = 1'h0; 1: mux_13222 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13223;
  wire [0:0] v_13224;
  wire [0:0] v_13225;
  wire [0:0] v_13226;
  wire [0:0] v_13227;
  wire [0:0] v_13228;
  wire [0:0] v_13229;
  function [0:0] mux_13229(input [0:0] sel);
    case (sel) 0: mux_13229 = 1'h0; 1: mux_13229 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13230;
  wire [0:0] v_13231;
  wire [0:0] v_13232;
  wire [0:0] v_13233;
  wire [0:0] v_13234;
  function [0:0] mux_13234(input [0:0] sel);
    case (sel) 0: mux_13234 = 1'h0; 1: mux_13234 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13235;
  wire [0:0] v_13236;
  wire [0:0] v_13237;
  wire [0:0] v_13238;
  function [0:0] mux_13238(input [0:0] sel);
    case (sel) 0: mux_13238 = 1'h0; 1: mux_13238 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13239;
  function [0:0] mux_13239(input [0:0] sel);
    case (sel) 0: mux_13239 = 1'h0; 1: mux_13239 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_13240 = 1'h0;
  wire [0:0] v_13241;
  wire [0:0] v_13242;
  wire [0:0] act_13243;
  wire [0:0] v_13244;
  wire [0:0] v_13245;
  wire [0:0] v_13246;
  wire [0:0] vin0_consume_en_13247;
  wire [0:0] vout_canPeek_13247;
  wire [7:0] vout_peek_13247;
  wire [0:0] v_13248;
  wire [0:0] v_13249;
  function [0:0] mux_13249(input [0:0] sel);
    case (sel) 0: mux_13249 = 1'h0; 1: mux_13249 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13250;
  wire [0:0] v_13251;
  wire [0:0] v_13252;
  wire [0:0] v_13253;
  wire [0:0] v_13254;
  function [0:0] mux_13254(input [0:0] sel);
    case (sel) 0: mux_13254 = 1'h0; 1: mux_13254 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13255;
  wire [0:0] vin0_consume_en_13256;
  wire [0:0] vout_canPeek_13256;
  wire [7:0] vout_peek_13256;
  wire [0:0] v_13257;
  wire [0:0] v_13258;
  function [0:0] mux_13258(input [0:0] sel);
    case (sel) 0: mux_13258 = 1'h0; 1: mux_13258 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13259;
  function [0:0] mux_13259(input [0:0] sel);
    case (sel) 0: mux_13259 = 1'h0; 1: mux_13259 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13260;
  wire [0:0] v_13261;
  wire [0:0] v_13262;
  wire [0:0] v_13263;
  wire [0:0] v_13264;
  wire [0:0] v_13265;
  wire [0:0] v_13266;
  function [0:0] mux_13266(input [0:0] sel);
    case (sel) 0: mux_13266 = 1'h0; 1: mux_13266 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13267;
  function [0:0] mux_13267(input [0:0] sel);
    case (sel) 0: mux_13267 = 1'h0; 1: mux_13267 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13268;
  wire [0:0] v_13269;
  wire [0:0] v_13270;
  wire [0:0] v_13271;
  function [0:0] mux_13271(input [0:0] sel);
    case (sel) 0: mux_13271 = 1'h0; 1: mux_13271 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13272;
  function [0:0] mux_13272(input [0:0] sel);
    case (sel) 0: mux_13272 = 1'h0; 1: mux_13272 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13273;
  wire [0:0] v_13274;
  wire [0:0] v_13275;
  wire [0:0] v_13276;
  wire [0:0] v_13277;
  wire [0:0] v_13278;
  function [0:0] mux_13278(input [0:0] sel);
    case (sel) 0: mux_13278 = 1'h0; 1: mux_13278 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13279;
  function [0:0] mux_13279(input [0:0] sel);
    case (sel) 0: mux_13279 = 1'h0; 1: mux_13279 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13280;
  wire [0:0] v_13281;
  wire [0:0] v_13282;
  wire [0:0] v_13283;
  function [0:0] mux_13283(input [0:0] sel);
    case (sel) 0: mux_13283 = 1'h0; 1: mux_13283 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13284;
  function [0:0] mux_13284(input [0:0] sel);
    case (sel) 0: mux_13284 = 1'h0; 1: mux_13284 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13285;
  wire [0:0] v_13286;
  wire [0:0] v_13287;
  wire [0:0] v_13288;
  wire [0:0] v_13289;
  wire [0:0] v_13290;
  function [0:0] mux_13290(input [0:0] sel);
    case (sel) 0: mux_13290 = 1'h0; 1: mux_13290 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13291;
  function [0:0] mux_13291(input [0:0] sel);
    case (sel) 0: mux_13291 = 1'h0; 1: mux_13291 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13292;
  wire [0:0] v_13293;
  wire [0:0] v_13294;
  wire [0:0] v_13295;
  function [0:0] mux_13295(input [0:0] sel);
    case (sel) 0: mux_13295 = 1'h0; 1: mux_13295 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13296;
  function [0:0] mux_13296(input [0:0] sel);
    case (sel) 0: mux_13296 = 1'h0; 1: mux_13296 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13297;
  wire [0:0] v_13298;
  wire [0:0] v_13299;
  wire [0:0] v_13300;
  wire [0:0] v_13301;
  wire [0:0] v_13302;
  function [0:0] mux_13302(input [0:0] sel);
    case (sel) 0: mux_13302 = 1'h0; 1: mux_13302 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13303;
  function [0:0] mux_13303(input [0:0] sel);
    case (sel) 0: mux_13303 = 1'h0; 1: mux_13303 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13304;
  wire [0:0] v_13305;
  wire [0:0] v_13306;
  wire [0:0] v_13307;
  function [0:0] mux_13307(input [0:0] sel);
    case (sel) 0: mux_13307 = 1'h0; 1: mux_13307 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13308;
  function [0:0] mux_13308(input [0:0] sel);
    case (sel) 0: mux_13308 = 1'h0; 1: mux_13308 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13309;
  wire [0:0] v_13310;
  wire [0:0] v_13311;
  wire [0:0] v_13312;
  wire [0:0] v_13313;
  wire [0:0] v_13314;
  function [0:0] mux_13314(input [0:0] sel);
    case (sel) 0: mux_13314 = 1'h0; 1: mux_13314 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13315;
  function [0:0] mux_13315(input [0:0] sel);
    case (sel) 0: mux_13315 = 1'h0; 1: mux_13315 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13316;
  wire [0:0] v_13317;
  wire [0:0] v_13318;
  wire [0:0] v_13319;
  function [0:0] mux_13319(input [0:0] sel);
    case (sel) 0: mux_13319 = 1'h0; 1: mux_13319 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13320;
  function [0:0] mux_13320(input [0:0] sel);
    case (sel) 0: mux_13320 = 1'h0; 1: mux_13320 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13321;
  wire [0:0] v_13322;
  wire [0:0] v_13323;
  wire [0:0] v_13324;
  wire [0:0] v_13325;
  wire [0:0] v_13326;
  function [0:0] mux_13326(input [0:0] sel);
    case (sel) 0: mux_13326 = 1'h0; 1: mux_13326 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13327;
  wire [0:0] v_13328;
  wire [0:0] v_13329;
  wire [0:0] v_13330;
  wire [0:0] v_13331;
  function [0:0] mux_13331(input [0:0] sel);
    case (sel) 0: mux_13331 = 1'h0; 1: mux_13331 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13332;
  wire [0:0] v_13333;
  wire [0:0] v_13334;
  wire [0:0] v_13335;
  function [0:0] mux_13335(input [0:0] sel);
    case (sel) 0: mux_13335 = 1'h0; 1: mux_13335 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13336;
  function [0:0] mux_13336(input [0:0] sel);
    case (sel) 0: mux_13336 = 1'h0; 1: mux_13336 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_13337 = 1'h0;
  wire [0:0] v_13338;
  wire [0:0] v_13339;
  wire [0:0] act_13340;
  wire [0:0] v_13341;
  wire [0:0] v_13342;
  wire [0:0] v_13343;
  reg [0:0] v_13344 = 1'h0;
  wire [0:0] v_13345;
  wire [0:0] v_13346;
  wire [0:0] act_13347;
  wire [0:0] v_13348;
  wire [0:0] v_13349;
  wire [0:0] v_13350;
  reg [0:0] v_13351 = 1'h0;
  wire [0:0] v_13352;
  wire [0:0] v_13353;
  wire [0:0] act_13354;
  wire [0:0] v_13355;
  wire [0:0] v_13356;
  wire [0:0] v_13357;
  reg [0:0] v_13358 = 1'h0;
  wire [0:0] v_13359;
  wire [0:0] v_13360;
  wire [0:0] act_13361;
  wire [0:0] v_13362;
  wire [0:0] v_13363;
  wire [0:0] v_13364;
  reg [0:0] v_13365 = 1'h0;
  wire [0:0] v_13366;
  wire [0:0] v_13367;
  wire [0:0] act_13368;
  wire [0:0] v_13369;
  wire [0:0] v_13370;
  wire [0:0] v_13371;
  reg [0:0] v_13372 = 1'h0;
  wire [0:0] v_13373;
  wire [0:0] v_13374;
  wire [0:0] act_13375;
  wire [0:0] v_13376;
  wire [0:0] v_13377;
  wire [0:0] v_13378;
  wire [0:0] vin0_consume_en_13379;
  wire [0:0] vout_canPeek_13379;
  wire [7:0] vout_peek_13379;
  wire [0:0] v_13380;
  wire [0:0] v_13381;
  function [0:0] mux_13381(input [0:0] sel);
    case (sel) 0: mux_13381 = 1'h0; 1: mux_13381 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13382;
  wire [0:0] v_13383;
  wire [0:0] v_13384;
  wire [0:0] v_13385;
  wire [0:0] v_13386;
  function [0:0] mux_13386(input [0:0] sel);
    case (sel) 0: mux_13386 = 1'h0; 1: mux_13386 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13387;
  wire [0:0] vin0_consume_en_13388;
  wire [0:0] vout_canPeek_13388;
  wire [7:0] vout_peek_13388;
  wire [0:0] v_13389;
  wire [0:0] v_13390;
  function [0:0] mux_13390(input [0:0] sel);
    case (sel) 0: mux_13390 = 1'h0; 1: mux_13390 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13391;
  function [0:0] mux_13391(input [0:0] sel);
    case (sel) 0: mux_13391 = 1'h0; 1: mux_13391 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13392;
  wire [0:0] v_13393;
  wire [0:0] v_13394;
  wire [0:0] v_13395;
  wire [0:0] v_13396;
  wire [0:0] v_13397;
  wire [0:0] v_13398;
  function [0:0] mux_13398(input [0:0] sel);
    case (sel) 0: mux_13398 = 1'h0; 1: mux_13398 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13399;
  wire [0:0] v_13400;
  wire [0:0] v_13401;
  wire [0:0] v_13402;
  wire [0:0] v_13403;
  function [0:0] mux_13403(input [0:0] sel);
    case (sel) 0: mux_13403 = 1'h0; 1: mux_13403 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13404;
  wire [0:0] v_13405;
  wire [0:0] v_13406;
  wire [0:0] v_13407;
  function [0:0] mux_13407(input [0:0] sel);
    case (sel) 0: mux_13407 = 1'h0; 1: mux_13407 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13408;
  function [0:0] mux_13408(input [0:0] sel);
    case (sel) 0: mux_13408 = 1'h0; 1: mux_13408 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_13409 = 1'h0;
  wire [0:0] v_13410;
  wire [0:0] v_13411;
  wire [0:0] act_13412;
  wire [0:0] v_13413;
  wire [0:0] v_13414;
  wire [0:0] v_13415;
  wire [0:0] vin0_consume_en_13416;
  wire [0:0] vout_canPeek_13416;
  wire [7:0] vout_peek_13416;
  wire [0:0] v_13417;
  wire [0:0] v_13418;
  function [0:0] mux_13418(input [0:0] sel);
    case (sel) 0: mux_13418 = 1'h0; 1: mux_13418 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13419;
  wire [0:0] v_13420;
  wire [0:0] v_13421;
  wire [0:0] v_13422;
  wire [0:0] v_13423;
  function [0:0] mux_13423(input [0:0] sel);
    case (sel) 0: mux_13423 = 1'h0; 1: mux_13423 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13424;
  wire [0:0] vin0_consume_en_13425;
  wire [0:0] vout_canPeek_13425;
  wire [7:0] vout_peek_13425;
  wire [0:0] v_13426;
  wire [0:0] v_13427;
  function [0:0] mux_13427(input [0:0] sel);
    case (sel) 0: mux_13427 = 1'h0; 1: mux_13427 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13428;
  function [0:0] mux_13428(input [0:0] sel);
    case (sel) 0: mux_13428 = 1'h0; 1: mux_13428 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13429;
  wire [0:0] v_13430;
  wire [0:0] v_13431;
  wire [0:0] v_13432;
  wire [0:0] v_13433;
  wire [0:0] v_13434;
  wire [0:0] v_13435;
  function [0:0] mux_13435(input [0:0] sel);
    case (sel) 0: mux_13435 = 1'h0; 1: mux_13435 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13436;
  function [0:0] mux_13436(input [0:0] sel);
    case (sel) 0: mux_13436 = 1'h0; 1: mux_13436 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13437;
  wire [0:0] v_13438;
  wire [0:0] v_13439;
  wire [0:0] v_13440;
  function [0:0] mux_13440(input [0:0] sel);
    case (sel) 0: mux_13440 = 1'h0; 1: mux_13440 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13441;
  function [0:0] mux_13441(input [0:0] sel);
    case (sel) 0: mux_13441 = 1'h0; 1: mux_13441 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13442;
  wire [0:0] v_13443;
  wire [0:0] v_13444;
  wire [0:0] v_13445;
  wire [0:0] v_13446;
  wire [0:0] v_13447;
  function [0:0] mux_13447(input [0:0] sel);
    case (sel) 0: mux_13447 = 1'h0; 1: mux_13447 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13448;
  wire [0:0] v_13449;
  wire [0:0] v_13450;
  wire [0:0] v_13451;
  wire [0:0] v_13452;
  function [0:0] mux_13452(input [0:0] sel);
    case (sel) 0: mux_13452 = 1'h0; 1: mux_13452 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13453;
  wire [0:0] v_13454;
  wire [0:0] v_13455;
  wire [0:0] v_13456;
  function [0:0] mux_13456(input [0:0] sel);
    case (sel) 0: mux_13456 = 1'h0; 1: mux_13456 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13457;
  function [0:0] mux_13457(input [0:0] sel);
    case (sel) 0: mux_13457 = 1'h0; 1: mux_13457 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_13458 = 1'h0;
  wire [0:0] v_13459;
  wire [0:0] v_13460;
  wire [0:0] act_13461;
  wire [0:0] v_13462;
  wire [0:0] v_13463;
  wire [0:0] v_13464;
  reg [0:0] v_13465 = 1'h0;
  wire [0:0] v_13466;
  wire [0:0] v_13467;
  wire [0:0] act_13468;
  wire [0:0] v_13469;
  wire [0:0] v_13470;
  wire [0:0] v_13471;
  wire [0:0] vin0_consume_en_13472;
  wire [0:0] vout_canPeek_13472;
  wire [7:0] vout_peek_13472;
  wire [0:0] v_13473;
  wire [0:0] v_13474;
  function [0:0] mux_13474(input [0:0] sel);
    case (sel) 0: mux_13474 = 1'h0; 1: mux_13474 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13475;
  wire [0:0] v_13476;
  wire [0:0] v_13477;
  wire [0:0] v_13478;
  wire [0:0] v_13479;
  function [0:0] mux_13479(input [0:0] sel);
    case (sel) 0: mux_13479 = 1'h0; 1: mux_13479 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13480;
  wire [0:0] vin0_consume_en_13481;
  wire [0:0] vout_canPeek_13481;
  wire [7:0] vout_peek_13481;
  wire [0:0] v_13482;
  wire [0:0] v_13483;
  function [0:0] mux_13483(input [0:0] sel);
    case (sel) 0: mux_13483 = 1'h0; 1: mux_13483 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13484;
  function [0:0] mux_13484(input [0:0] sel);
    case (sel) 0: mux_13484 = 1'h0; 1: mux_13484 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13485;
  wire [0:0] v_13486;
  wire [0:0] v_13487;
  wire [0:0] v_13488;
  wire [0:0] v_13489;
  wire [0:0] v_13490;
  wire [0:0] v_13491;
  function [0:0] mux_13491(input [0:0] sel);
    case (sel) 0: mux_13491 = 1'h0; 1: mux_13491 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13492;
  wire [0:0] v_13493;
  wire [0:0] v_13494;
  wire [0:0] v_13495;
  wire [0:0] v_13496;
  function [0:0] mux_13496(input [0:0] sel);
    case (sel) 0: mux_13496 = 1'h0; 1: mux_13496 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13497;
  wire [0:0] v_13498;
  wire [0:0] v_13499;
  wire [0:0] v_13500;
  function [0:0] mux_13500(input [0:0] sel);
    case (sel) 0: mux_13500 = 1'h0; 1: mux_13500 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13501;
  function [0:0] mux_13501(input [0:0] sel);
    case (sel) 0: mux_13501 = 1'h0; 1: mux_13501 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_13502 = 1'h0;
  wire [0:0] v_13503;
  wire [0:0] v_13504;
  wire [0:0] act_13505;
  wire [0:0] v_13506;
  wire [0:0] v_13507;
  wire [0:0] v_13508;
  wire [0:0] vin0_consume_en_13509;
  wire [0:0] vout_canPeek_13509;
  wire [7:0] vout_peek_13509;
  wire [0:0] v_13510;
  wire [0:0] v_13511;
  function [0:0] mux_13511(input [0:0] sel);
    case (sel) 0: mux_13511 = 1'h0; 1: mux_13511 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13512;
  wire [0:0] v_13513;
  wire [0:0] v_13514;
  wire [0:0] v_13515;
  wire [0:0] v_13516;
  function [0:0] mux_13516(input [0:0] sel);
    case (sel) 0: mux_13516 = 1'h0; 1: mux_13516 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13517;
  wire [0:0] vin0_consume_en_13518;
  wire [0:0] vout_canPeek_13518;
  wire [7:0] vout_peek_13518;
  wire [0:0] v_13519;
  wire [0:0] v_13520;
  function [0:0] mux_13520(input [0:0] sel);
    case (sel) 0: mux_13520 = 1'h0; 1: mux_13520 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13521;
  function [0:0] mux_13521(input [0:0] sel);
    case (sel) 0: mux_13521 = 1'h0; 1: mux_13521 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13522;
  wire [0:0] v_13523;
  wire [0:0] v_13524;
  wire [0:0] v_13525;
  wire [0:0] v_13526;
  wire [0:0] v_13527;
  wire [0:0] v_13528;
  function [0:0] mux_13528(input [0:0] sel);
    case (sel) 0: mux_13528 = 1'h0; 1: mux_13528 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13529;
  function [0:0] mux_13529(input [0:0] sel);
    case (sel) 0: mux_13529 = 1'h0; 1: mux_13529 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13530;
  wire [0:0] v_13531;
  wire [0:0] v_13532;
  wire [0:0] v_13533;
  function [0:0] mux_13533(input [0:0] sel);
    case (sel) 0: mux_13533 = 1'h0; 1: mux_13533 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13534;
  function [0:0] mux_13534(input [0:0] sel);
    case (sel) 0: mux_13534 = 1'h0; 1: mux_13534 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13535;
  wire [0:0] v_13536;
  wire [0:0] v_13537;
  wire [0:0] v_13538;
  wire [0:0] v_13539;
  wire [0:0] v_13540;
  function [0:0] mux_13540(input [0:0] sel);
    case (sel) 0: mux_13540 = 1'h0; 1: mux_13540 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13541;
  function [0:0] mux_13541(input [0:0] sel);
    case (sel) 0: mux_13541 = 1'h0; 1: mux_13541 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13542;
  wire [0:0] v_13543;
  wire [0:0] v_13544;
  wire [0:0] v_13545;
  function [0:0] mux_13545(input [0:0] sel);
    case (sel) 0: mux_13545 = 1'h0; 1: mux_13545 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13546;
  function [0:0] mux_13546(input [0:0] sel);
    case (sel) 0: mux_13546 = 1'h0; 1: mux_13546 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13547;
  wire [0:0] v_13548;
  wire [0:0] v_13549;
  wire [0:0] v_13550;
  wire [0:0] v_13551;
  wire [0:0] v_13552;
  function [0:0] mux_13552(input [0:0] sel);
    case (sel) 0: mux_13552 = 1'h0; 1: mux_13552 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13553;
  wire [0:0] v_13554;
  wire [0:0] v_13555;
  wire [0:0] v_13556;
  wire [0:0] v_13557;
  function [0:0] mux_13557(input [0:0] sel);
    case (sel) 0: mux_13557 = 1'h0; 1: mux_13557 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13558;
  wire [0:0] v_13559;
  wire [0:0] v_13560;
  wire [0:0] v_13561;
  function [0:0] mux_13561(input [0:0] sel);
    case (sel) 0: mux_13561 = 1'h0; 1: mux_13561 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13562;
  function [0:0] mux_13562(input [0:0] sel);
    case (sel) 0: mux_13562 = 1'h0; 1: mux_13562 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_13563 = 1'h0;
  wire [0:0] v_13564;
  wire [0:0] v_13565;
  wire [0:0] act_13566;
  wire [0:0] v_13567;
  wire [0:0] v_13568;
  wire [0:0] v_13569;
  reg [0:0] v_13570 = 1'h0;
  wire [0:0] v_13571;
  wire [0:0] v_13572;
  wire [0:0] act_13573;
  wire [0:0] v_13574;
  wire [0:0] v_13575;
  wire [0:0] v_13576;
  reg [0:0] v_13577 = 1'h0;
  wire [0:0] v_13578;
  wire [0:0] v_13579;
  wire [0:0] act_13580;
  wire [0:0] v_13581;
  wire [0:0] v_13582;
  wire [0:0] v_13583;
  wire [0:0] vin0_consume_en_13584;
  wire [0:0] vout_canPeek_13584;
  wire [7:0] vout_peek_13584;
  wire [0:0] v_13585;
  wire [0:0] v_13586;
  function [0:0] mux_13586(input [0:0] sel);
    case (sel) 0: mux_13586 = 1'h0; 1: mux_13586 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13587;
  wire [0:0] v_13588;
  wire [0:0] v_13589;
  wire [0:0] v_13590;
  wire [0:0] v_13591;
  function [0:0] mux_13591(input [0:0] sel);
    case (sel) 0: mux_13591 = 1'h0; 1: mux_13591 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13592;
  wire [0:0] vin0_consume_en_13593;
  wire [0:0] vout_canPeek_13593;
  wire [7:0] vout_peek_13593;
  wire [0:0] v_13594;
  wire [0:0] v_13595;
  function [0:0] mux_13595(input [0:0] sel);
    case (sel) 0: mux_13595 = 1'h0; 1: mux_13595 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13596;
  function [0:0] mux_13596(input [0:0] sel);
    case (sel) 0: mux_13596 = 1'h0; 1: mux_13596 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13597;
  wire [0:0] v_13598;
  wire [0:0] v_13599;
  wire [0:0] v_13600;
  wire [0:0] v_13601;
  wire [0:0] v_13602;
  wire [0:0] v_13603;
  function [0:0] mux_13603(input [0:0] sel);
    case (sel) 0: mux_13603 = 1'h0; 1: mux_13603 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13604;
  wire [0:0] v_13605;
  wire [0:0] v_13606;
  wire [0:0] v_13607;
  wire [0:0] v_13608;
  function [0:0] mux_13608(input [0:0] sel);
    case (sel) 0: mux_13608 = 1'h0; 1: mux_13608 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13609;
  wire [0:0] v_13610;
  wire [0:0] v_13611;
  wire [0:0] v_13612;
  function [0:0] mux_13612(input [0:0] sel);
    case (sel) 0: mux_13612 = 1'h0; 1: mux_13612 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13613;
  function [0:0] mux_13613(input [0:0] sel);
    case (sel) 0: mux_13613 = 1'h0; 1: mux_13613 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_13614 = 1'h0;
  wire [0:0] v_13615;
  wire [0:0] v_13616;
  wire [0:0] act_13617;
  wire [0:0] v_13618;
  wire [0:0] v_13619;
  wire [0:0] v_13620;
  wire [0:0] vin0_consume_en_13621;
  wire [0:0] vout_canPeek_13621;
  wire [7:0] vout_peek_13621;
  wire [0:0] v_13622;
  wire [0:0] v_13623;
  function [0:0] mux_13623(input [0:0] sel);
    case (sel) 0: mux_13623 = 1'h0; 1: mux_13623 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13624;
  wire [0:0] v_13625;
  wire [0:0] v_13626;
  wire [0:0] v_13627;
  wire [0:0] v_13628;
  function [0:0] mux_13628(input [0:0] sel);
    case (sel) 0: mux_13628 = 1'h0; 1: mux_13628 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13629;
  wire [0:0] vin0_consume_en_13630;
  wire [0:0] vout_canPeek_13630;
  wire [7:0] vout_peek_13630;
  wire [0:0] v_13631;
  wire [0:0] v_13632;
  function [0:0] mux_13632(input [0:0] sel);
    case (sel) 0: mux_13632 = 1'h0; 1: mux_13632 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13633;
  function [0:0] mux_13633(input [0:0] sel);
    case (sel) 0: mux_13633 = 1'h0; 1: mux_13633 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13634;
  wire [0:0] v_13635;
  wire [0:0] v_13636;
  wire [0:0] v_13637;
  wire [0:0] v_13638;
  wire [0:0] v_13639;
  wire [0:0] v_13640;
  function [0:0] mux_13640(input [0:0] sel);
    case (sel) 0: mux_13640 = 1'h0; 1: mux_13640 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13641;
  function [0:0] mux_13641(input [0:0] sel);
    case (sel) 0: mux_13641 = 1'h0; 1: mux_13641 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13642;
  wire [0:0] v_13643;
  wire [0:0] v_13644;
  wire [0:0] v_13645;
  function [0:0] mux_13645(input [0:0] sel);
    case (sel) 0: mux_13645 = 1'h0; 1: mux_13645 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13646;
  function [0:0] mux_13646(input [0:0] sel);
    case (sel) 0: mux_13646 = 1'h0; 1: mux_13646 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13647;
  wire [0:0] v_13648;
  wire [0:0] v_13649;
  wire [0:0] v_13650;
  wire [0:0] v_13651;
  wire [0:0] v_13652;
  function [0:0] mux_13652(input [0:0] sel);
    case (sel) 0: mux_13652 = 1'h0; 1: mux_13652 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13653;
  wire [0:0] v_13654;
  wire [0:0] v_13655;
  wire [0:0] v_13656;
  wire [0:0] v_13657;
  function [0:0] mux_13657(input [0:0] sel);
    case (sel) 0: mux_13657 = 1'h0; 1: mux_13657 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13658;
  wire [0:0] v_13659;
  wire [0:0] v_13660;
  wire [0:0] v_13661;
  function [0:0] mux_13661(input [0:0] sel);
    case (sel) 0: mux_13661 = 1'h0; 1: mux_13661 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13662;
  function [0:0] mux_13662(input [0:0] sel);
    case (sel) 0: mux_13662 = 1'h0; 1: mux_13662 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_13663 = 1'h0;
  wire [0:0] v_13664;
  wire [0:0] v_13665;
  wire [0:0] act_13666;
  wire [0:0] v_13667;
  wire [0:0] v_13668;
  wire [0:0] v_13669;
  reg [0:0] v_13670 = 1'h0;
  wire [0:0] v_13671;
  wire [0:0] v_13672;
  wire [0:0] act_13673;
  wire [0:0] v_13674;
  wire [0:0] v_13675;
  wire [0:0] v_13676;
  wire [0:0] vin0_consume_en_13677;
  wire [0:0] vout_canPeek_13677;
  wire [7:0] vout_peek_13677;
  wire [0:0] v_13678;
  wire [0:0] v_13679;
  function [0:0] mux_13679(input [0:0] sel);
    case (sel) 0: mux_13679 = 1'h0; 1: mux_13679 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13680;
  wire [0:0] v_13681;
  wire [0:0] v_13682;
  wire [0:0] v_13683;
  wire [0:0] v_13684;
  function [0:0] mux_13684(input [0:0] sel);
    case (sel) 0: mux_13684 = 1'h0; 1: mux_13684 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13685;
  wire [0:0] vin0_consume_en_13686;
  wire [0:0] vout_canPeek_13686;
  wire [7:0] vout_peek_13686;
  wire [0:0] v_13687;
  wire [0:0] v_13688;
  function [0:0] mux_13688(input [0:0] sel);
    case (sel) 0: mux_13688 = 1'h0; 1: mux_13688 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13689;
  function [0:0] mux_13689(input [0:0] sel);
    case (sel) 0: mux_13689 = 1'h0; 1: mux_13689 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13690;
  wire [0:0] v_13691;
  wire [0:0] v_13692;
  wire [0:0] v_13693;
  wire [0:0] v_13694;
  wire [0:0] v_13695;
  wire [0:0] v_13696;
  function [0:0] mux_13696(input [0:0] sel);
    case (sel) 0: mux_13696 = 1'h0; 1: mux_13696 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13697;
  wire [0:0] v_13698;
  wire [0:0] v_13699;
  wire [0:0] v_13700;
  wire [0:0] v_13701;
  function [0:0] mux_13701(input [0:0] sel);
    case (sel) 0: mux_13701 = 1'h0; 1: mux_13701 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13702;
  wire [0:0] v_13703;
  wire [0:0] v_13704;
  wire [0:0] v_13705;
  function [0:0] mux_13705(input [0:0] sel);
    case (sel) 0: mux_13705 = 1'h0; 1: mux_13705 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13706;
  function [0:0] mux_13706(input [0:0] sel);
    case (sel) 0: mux_13706 = 1'h0; 1: mux_13706 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_13707 = 1'h0;
  wire [0:0] v_13708;
  wire [0:0] v_13709;
  wire [0:0] act_13710;
  wire [0:0] v_13711;
  wire [0:0] v_13712;
  wire [0:0] v_13713;
  wire [0:0] vin0_consume_en_13714;
  wire [0:0] vout_canPeek_13714;
  wire [7:0] vout_peek_13714;
  wire [0:0] v_13715;
  wire [0:0] v_13716;
  function [0:0] mux_13716(input [0:0] sel);
    case (sel) 0: mux_13716 = 1'h0; 1: mux_13716 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13717;
  wire [0:0] v_13718;
  wire [0:0] v_13719;
  wire [0:0] v_13720;
  wire [0:0] v_13721;
  function [0:0] mux_13721(input [0:0] sel);
    case (sel) 0: mux_13721 = 1'h0; 1: mux_13721 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13722;
  wire [0:0] vin0_consume_en_13723;
  wire [0:0] vout_canPeek_13723;
  wire [7:0] vout_peek_13723;
  wire [0:0] v_13724;
  wire [0:0] v_13725;
  function [0:0] mux_13725(input [0:0] sel);
    case (sel) 0: mux_13725 = 1'h0; 1: mux_13725 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13726;
  function [0:0] mux_13726(input [0:0] sel);
    case (sel) 0: mux_13726 = 1'h0; 1: mux_13726 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13727;
  wire [0:0] v_13728;
  wire [0:0] v_13729;
  wire [0:0] v_13730;
  wire [0:0] v_13731;
  wire [0:0] v_13732;
  wire [0:0] v_13733;
  function [0:0] mux_13733(input [0:0] sel);
    case (sel) 0: mux_13733 = 1'h0; 1: mux_13733 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13734;
  function [0:0] mux_13734(input [0:0] sel);
    case (sel) 0: mux_13734 = 1'h0; 1: mux_13734 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13735;
  wire [0:0] v_13736;
  wire [0:0] v_13737;
  wire [0:0] v_13738;
  function [0:0] mux_13738(input [0:0] sel);
    case (sel) 0: mux_13738 = 1'h0; 1: mux_13738 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13739;
  function [0:0] mux_13739(input [0:0] sel);
    case (sel) 0: mux_13739 = 1'h0; 1: mux_13739 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13740;
  wire [0:0] v_13741;
  wire [0:0] v_13742;
  wire [0:0] v_13743;
  wire [0:0] v_13744;
  wire [0:0] v_13745;
  function [0:0] mux_13745(input [0:0] sel);
    case (sel) 0: mux_13745 = 1'h0; 1: mux_13745 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13746;
  function [0:0] mux_13746(input [0:0] sel);
    case (sel) 0: mux_13746 = 1'h0; 1: mux_13746 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13747;
  wire [0:0] v_13748;
  wire [0:0] v_13749;
  wire [0:0] v_13750;
  function [0:0] mux_13750(input [0:0] sel);
    case (sel) 0: mux_13750 = 1'h0; 1: mux_13750 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13751;
  function [0:0] mux_13751(input [0:0] sel);
    case (sel) 0: mux_13751 = 1'h0; 1: mux_13751 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13752;
  wire [0:0] v_13753;
  wire [0:0] v_13754;
  wire [0:0] v_13755;
  wire [0:0] v_13756;
  wire [0:0] v_13757;
  function [0:0] mux_13757(input [0:0] sel);
    case (sel) 0: mux_13757 = 1'h0; 1: mux_13757 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13758;
  function [0:0] mux_13758(input [0:0] sel);
    case (sel) 0: mux_13758 = 1'h0; 1: mux_13758 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13759;
  wire [0:0] v_13760;
  wire [0:0] v_13761;
  wire [0:0] v_13762;
  function [0:0] mux_13762(input [0:0] sel);
    case (sel) 0: mux_13762 = 1'h0; 1: mux_13762 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13763;
  function [0:0] mux_13763(input [0:0] sel);
    case (sel) 0: mux_13763 = 1'h0; 1: mux_13763 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13764;
  wire [0:0] v_13765;
  wire [0:0] v_13766;
  wire [0:0] v_13767;
  wire [0:0] v_13768;
  wire [0:0] v_13769;
  function [0:0] mux_13769(input [0:0] sel);
    case (sel) 0: mux_13769 = 1'h0; 1: mux_13769 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13770;
  wire [0:0] v_13771;
  wire [0:0] v_13772;
  wire [0:0] v_13773;
  wire [0:0] v_13774;
  function [0:0] mux_13774(input [0:0] sel);
    case (sel) 0: mux_13774 = 1'h0; 1: mux_13774 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13775;
  wire [0:0] v_13776;
  wire [0:0] v_13777;
  wire [0:0] v_13778;
  function [0:0] mux_13778(input [0:0] sel);
    case (sel) 0: mux_13778 = 1'h0; 1: mux_13778 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13779;
  function [0:0] mux_13779(input [0:0] sel);
    case (sel) 0: mux_13779 = 1'h0; 1: mux_13779 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_13780 = 1'h0;
  wire [0:0] v_13781;
  wire [0:0] v_13782;
  wire [0:0] act_13783;
  wire [0:0] v_13784;
  wire [0:0] v_13785;
  wire [0:0] v_13786;
  reg [0:0] v_13787 = 1'h0;
  wire [0:0] v_13788;
  wire [0:0] v_13789;
  wire [0:0] act_13790;
  wire [0:0] v_13791;
  wire [0:0] v_13792;
  wire [0:0] v_13793;
  reg [0:0] v_13794 = 1'h0;
  wire [0:0] v_13795;
  wire [0:0] v_13796;
  wire [0:0] act_13797;
  wire [0:0] v_13798;
  wire [0:0] v_13799;
  wire [0:0] v_13800;
  reg [0:0] v_13801 = 1'h0;
  wire [0:0] v_13802;
  wire [0:0] v_13803;
  wire [0:0] act_13804;
  wire [0:0] v_13805;
  wire [0:0] v_13806;
  wire [0:0] v_13807;
  wire [0:0] vin0_consume_en_13808;
  wire [0:0] vout_canPeek_13808;
  wire [7:0] vout_peek_13808;
  wire [0:0] v_13809;
  wire [0:0] v_13810;
  function [0:0] mux_13810(input [0:0] sel);
    case (sel) 0: mux_13810 = 1'h0; 1: mux_13810 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13811;
  wire [0:0] v_13812;
  wire [0:0] v_13813;
  wire [0:0] v_13814;
  wire [0:0] v_13815;
  function [0:0] mux_13815(input [0:0] sel);
    case (sel) 0: mux_13815 = 1'h0; 1: mux_13815 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13816;
  wire [0:0] vin0_consume_en_13817;
  wire [0:0] vout_canPeek_13817;
  wire [7:0] vout_peek_13817;
  wire [0:0] v_13818;
  wire [0:0] v_13819;
  function [0:0] mux_13819(input [0:0] sel);
    case (sel) 0: mux_13819 = 1'h0; 1: mux_13819 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13820;
  function [0:0] mux_13820(input [0:0] sel);
    case (sel) 0: mux_13820 = 1'h0; 1: mux_13820 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13821;
  wire [0:0] v_13822;
  wire [0:0] v_13823;
  wire [0:0] v_13824;
  wire [0:0] v_13825;
  wire [0:0] v_13826;
  wire [0:0] v_13827;
  function [0:0] mux_13827(input [0:0] sel);
    case (sel) 0: mux_13827 = 1'h0; 1: mux_13827 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13828;
  wire [0:0] v_13829;
  wire [0:0] v_13830;
  wire [0:0] v_13831;
  wire [0:0] v_13832;
  function [0:0] mux_13832(input [0:0] sel);
    case (sel) 0: mux_13832 = 1'h0; 1: mux_13832 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13833;
  wire [0:0] v_13834;
  wire [0:0] v_13835;
  wire [0:0] v_13836;
  function [0:0] mux_13836(input [0:0] sel);
    case (sel) 0: mux_13836 = 1'h0; 1: mux_13836 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13837;
  function [0:0] mux_13837(input [0:0] sel);
    case (sel) 0: mux_13837 = 1'h0; 1: mux_13837 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_13838 = 1'h0;
  wire [0:0] v_13839;
  wire [0:0] v_13840;
  wire [0:0] act_13841;
  wire [0:0] v_13842;
  wire [0:0] v_13843;
  wire [0:0] v_13844;
  wire [0:0] vin0_consume_en_13845;
  wire [0:0] vout_canPeek_13845;
  wire [7:0] vout_peek_13845;
  wire [0:0] v_13846;
  wire [0:0] v_13847;
  function [0:0] mux_13847(input [0:0] sel);
    case (sel) 0: mux_13847 = 1'h0; 1: mux_13847 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13848;
  wire [0:0] v_13849;
  wire [0:0] v_13850;
  wire [0:0] v_13851;
  wire [0:0] v_13852;
  function [0:0] mux_13852(input [0:0] sel);
    case (sel) 0: mux_13852 = 1'h0; 1: mux_13852 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13853;
  wire [0:0] vin0_consume_en_13854;
  wire [0:0] vout_canPeek_13854;
  wire [7:0] vout_peek_13854;
  wire [0:0] v_13855;
  wire [0:0] v_13856;
  function [0:0] mux_13856(input [0:0] sel);
    case (sel) 0: mux_13856 = 1'h0; 1: mux_13856 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13857;
  function [0:0] mux_13857(input [0:0] sel);
    case (sel) 0: mux_13857 = 1'h0; 1: mux_13857 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13858;
  wire [0:0] v_13859;
  wire [0:0] v_13860;
  wire [0:0] v_13861;
  wire [0:0] v_13862;
  wire [0:0] v_13863;
  wire [0:0] v_13864;
  function [0:0] mux_13864(input [0:0] sel);
    case (sel) 0: mux_13864 = 1'h0; 1: mux_13864 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13865;
  function [0:0] mux_13865(input [0:0] sel);
    case (sel) 0: mux_13865 = 1'h0; 1: mux_13865 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13866;
  wire [0:0] v_13867;
  wire [0:0] v_13868;
  wire [0:0] v_13869;
  function [0:0] mux_13869(input [0:0] sel);
    case (sel) 0: mux_13869 = 1'h0; 1: mux_13869 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13870;
  function [0:0] mux_13870(input [0:0] sel);
    case (sel) 0: mux_13870 = 1'h0; 1: mux_13870 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13871;
  wire [0:0] v_13872;
  wire [0:0] v_13873;
  wire [0:0] v_13874;
  wire [0:0] v_13875;
  wire [0:0] v_13876;
  function [0:0] mux_13876(input [0:0] sel);
    case (sel) 0: mux_13876 = 1'h0; 1: mux_13876 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13877;
  wire [0:0] v_13878;
  wire [0:0] v_13879;
  wire [0:0] v_13880;
  wire [0:0] v_13881;
  function [0:0] mux_13881(input [0:0] sel);
    case (sel) 0: mux_13881 = 1'h0; 1: mux_13881 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13882;
  wire [0:0] v_13883;
  wire [0:0] v_13884;
  wire [0:0] v_13885;
  function [0:0] mux_13885(input [0:0] sel);
    case (sel) 0: mux_13885 = 1'h0; 1: mux_13885 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13886;
  function [0:0] mux_13886(input [0:0] sel);
    case (sel) 0: mux_13886 = 1'h0; 1: mux_13886 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_13887 = 1'h0;
  wire [0:0] v_13888;
  wire [0:0] v_13889;
  wire [0:0] act_13890;
  wire [0:0] v_13891;
  wire [0:0] v_13892;
  wire [0:0] v_13893;
  reg [0:0] v_13894 = 1'h0;
  wire [0:0] v_13895;
  wire [0:0] v_13896;
  wire [0:0] act_13897;
  wire [0:0] v_13898;
  wire [0:0] v_13899;
  wire [0:0] v_13900;
  wire [0:0] vin0_consume_en_13901;
  wire [0:0] vout_canPeek_13901;
  wire [7:0] vout_peek_13901;
  wire [0:0] v_13902;
  wire [0:0] v_13903;
  function [0:0] mux_13903(input [0:0] sel);
    case (sel) 0: mux_13903 = 1'h0; 1: mux_13903 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13904;
  wire [0:0] v_13905;
  wire [0:0] v_13906;
  wire [0:0] v_13907;
  wire [0:0] v_13908;
  function [0:0] mux_13908(input [0:0] sel);
    case (sel) 0: mux_13908 = 1'h0; 1: mux_13908 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13909;
  wire [0:0] vin0_consume_en_13910;
  wire [0:0] vout_canPeek_13910;
  wire [7:0] vout_peek_13910;
  wire [0:0] v_13911;
  wire [0:0] v_13912;
  function [0:0] mux_13912(input [0:0] sel);
    case (sel) 0: mux_13912 = 1'h0; 1: mux_13912 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13913;
  function [0:0] mux_13913(input [0:0] sel);
    case (sel) 0: mux_13913 = 1'h0; 1: mux_13913 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13914;
  wire [0:0] v_13915;
  wire [0:0] v_13916;
  wire [0:0] v_13917;
  wire [0:0] v_13918;
  wire [0:0] v_13919;
  wire [0:0] v_13920;
  function [0:0] mux_13920(input [0:0] sel);
    case (sel) 0: mux_13920 = 1'h0; 1: mux_13920 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13921;
  wire [0:0] v_13922;
  wire [0:0] v_13923;
  wire [0:0] v_13924;
  wire [0:0] v_13925;
  function [0:0] mux_13925(input [0:0] sel);
    case (sel) 0: mux_13925 = 1'h0; 1: mux_13925 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13926;
  wire [0:0] v_13927;
  wire [0:0] v_13928;
  wire [0:0] v_13929;
  function [0:0] mux_13929(input [0:0] sel);
    case (sel) 0: mux_13929 = 1'h0; 1: mux_13929 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13930;
  function [0:0] mux_13930(input [0:0] sel);
    case (sel) 0: mux_13930 = 1'h0; 1: mux_13930 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_13931 = 1'h0;
  wire [0:0] v_13932;
  wire [0:0] v_13933;
  wire [0:0] act_13934;
  wire [0:0] v_13935;
  wire [0:0] v_13936;
  wire [0:0] v_13937;
  wire [0:0] vin0_consume_en_13938;
  wire [0:0] vout_canPeek_13938;
  wire [7:0] vout_peek_13938;
  wire [0:0] v_13939;
  wire [0:0] v_13940;
  function [0:0] mux_13940(input [0:0] sel);
    case (sel) 0: mux_13940 = 1'h0; 1: mux_13940 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13941;
  wire [0:0] v_13942;
  wire [0:0] v_13943;
  wire [0:0] v_13944;
  wire [0:0] v_13945;
  function [0:0] mux_13945(input [0:0] sel);
    case (sel) 0: mux_13945 = 1'h0; 1: mux_13945 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13946;
  wire [0:0] vin0_consume_en_13947;
  wire [0:0] vout_canPeek_13947;
  wire [7:0] vout_peek_13947;
  wire [0:0] v_13948;
  wire [0:0] v_13949;
  function [0:0] mux_13949(input [0:0] sel);
    case (sel) 0: mux_13949 = 1'h0; 1: mux_13949 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13950;
  function [0:0] mux_13950(input [0:0] sel);
    case (sel) 0: mux_13950 = 1'h0; 1: mux_13950 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13951;
  wire [0:0] v_13952;
  wire [0:0] v_13953;
  wire [0:0] v_13954;
  wire [0:0] v_13955;
  wire [0:0] v_13956;
  wire [0:0] v_13957;
  function [0:0] mux_13957(input [0:0] sel);
    case (sel) 0: mux_13957 = 1'h0; 1: mux_13957 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13958;
  function [0:0] mux_13958(input [0:0] sel);
    case (sel) 0: mux_13958 = 1'h0; 1: mux_13958 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13959;
  wire [0:0] v_13960;
  wire [0:0] v_13961;
  wire [0:0] v_13962;
  function [0:0] mux_13962(input [0:0] sel);
    case (sel) 0: mux_13962 = 1'h0; 1: mux_13962 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13963;
  function [0:0] mux_13963(input [0:0] sel);
    case (sel) 0: mux_13963 = 1'h0; 1: mux_13963 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13964;
  wire [0:0] v_13965;
  wire [0:0] v_13966;
  wire [0:0] v_13967;
  wire [0:0] v_13968;
  wire [0:0] v_13969;
  function [0:0] mux_13969(input [0:0] sel);
    case (sel) 0: mux_13969 = 1'h0; 1: mux_13969 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13970;
  function [0:0] mux_13970(input [0:0] sel);
    case (sel) 0: mux_13970 = 1'h0; 1: mux_13970 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13971;
  wire [0:0] v_13972;
  wire [0:0] v_13973;
  wire [0:0] v_13974;
  function [0:0] mux_13974(input [0:0] sel);
    case (sel) 0: mux_13974 = 1'h0; 1: mux_13974 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13975;
  function [0:0] mux_13975(input [0:0] sel);
    case (sel) 0: mux_13975 = 1'h0; 1: mux_13975 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13976;
  wire [0:0] v_13977;
  wire [0:0] v_13978;
  wire [0:0] v_13979;
  wire [0:0] v_13980;
  wire [0:0] v_13981;
  function [0:0] mux_13981(input [0:0] sel);
    case (sel) 0: mux_13981 = 1'h0; 1: mux_13981 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13982;
  wire [0:0] v_13983;
  wire [0:0] v_13984;
  wire [0:0] v_13985;
  wire [0:0] v_13986;
  function [0:0] mux_13986(input [0:0] sel);
    case (sel) 0: mux_13986 = 1'h0; 1: mux_13986 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13987;
  wire [0:0] v_13988;
  wire [0:0] v_13989;
  wire [0:0] v_13990;
  function [0:0] mux_13990(input [0:0] sel);
    case (sel) 0: mux_13990 = 1'h0; 1: mux_13990 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_13991;
  function [0:0] mux_13991(input [0:0] sel);
    case (sel) 0: mux_13991 = 1'h0; 1: mux_13991 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_13992 = 1'h0;
  wire [0:0] v_13993;
  wire [0:0] v_13994;
  wire [0:0] act_13995;
  wire [0:0] v_13996;
  wire [0:0] v_13997;
  wire [0:0] v_13998;
  reg [0:0] v_13999 = 1'h0;
  wire [0:0] v_14000;
  wire [0:0] v_14001;
  wire [0:0] act_14002;
  wire [0:0] v_14003;
  wire [0:0] v_14004;
  wire [0:0] v_14005;
  reg [0:0] v_14006 = 1'h0;
  wire [0:0] v_14007;
  wire [0:0] v_14008;
  wire [0:0] act_14009;
  wire [0:0] v_14010;
  wire [0:0] v_14011;
  wire [0:0] v_14012;
  wire [0:0] vin0_consume_en_14013;
  wire [0:0] vout_canPeek_14013;
  wire [7:0] vout_peek_14013;
  wire [0:0] v_14014;
  wire [0:0] v_14015;
  function [0:0] mux_14015(input [0:0] sel);
    case (sel) 0: mux_14015 = 1'h0; 1: mux_14015 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14016;
  wire [0:0] v_14017;
  wire [0:0] v_14018;
  wire [0:0] v_14019;
  wire [0:0] v_14020;
  function [0:0] mux_14020(input [0:0] sel);
    case (sel) 0: mux_14020 = 1'h0; 1: mux_14020 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14021;
  wire [0:0] vin0_consume_en_14022;
  wire [0:0] vout_canPeek_14022;
  wire [7:0] vout_peek_14022;
  wire [0:0] v_14023;
  wire [0:0] v_14024;
  function [0:0] mux_14024(input [0:0] sel);
    case (sel) 0: mux_14024 = 1'h0; 1: mux_14024 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14025;
  function [0:0] mux_14025(input [0:0] sel);
    case (sel) 0: mux_14025 = 1'h0; 1: mux_14025 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14026;
  wire [0:0] v_14027;
  wire [0:0] v_14028;
  wire [0:0] v_14029;
  wire [0:0] v_14030;
  wire [0:0] v_14031;
  wire [0:0] v_14032;
  function [0:0] mux_14032(input [0:0] sel);
    case (sel) 0: mux_14032 = 1'h0; 1: mux_14032 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14033;
  wire [0:0] v_14034;
  wire [0:0] v_14035;
  wire [0:0] v_14036;
  wire [0:0] v_14037;
  function [0:0] mux_14037(input [0:0] sel);
    case (sel) 0: mux_14037 = 1'h0; 1: mux_14037 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14038;
  wire [0:0] v_14039;
  wire [0:0] v_14040;
  wire [0:0] v_14041;
  function [0:0] mux_14041(input [0:0] sel);
    case (sel) 0: mux_14041 = 1'h0; 1: mux_14041 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14042;
  function [0:0] mux_14042(input [0:0] sel);
    case (sel) 0: mux_14042 = 1'h0; 1: mux_14042 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_14043 = 1'h0;
  wire [0:0] v_14044;
  wire [0:0] v_14045;
  wire [0:0] act_14046;
  wire [0:0] v_14047;
  wire [0:0] v_14048;
  wire [0:0] v_14049;
  wire [0:0] vin0_consume_en_14050;
  wire [0:0] vout_canPeek_14050;
  wire [7:0] vout_peek_14050;
  wire [0:0] v_14051;
  wire [0:0] v_14052;
  function [0:0] mux_14052(input [0:0] sel);
    case (sel) 0: mux_14052 = 1'h0; 1: mux_14052 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14053;
  wire [0:0] v_14054;
  wire [0:0] v_14055;
  wire [0:0] v_14056;
  wire [0:0] v_14057;
  function [0:0] mux_14057(input [0:0] sel);
    case (sel) 0: mux_14057 = 1'h0; 1: mux_14057 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14058;
  wire [0:0] vin0_consume_en_14059;
  wire [0:0] vout_canPeek_14059;
  wire [7:0] vout_peek_14059;
  wire [0:0] v_14060;
  wire [0:0] v_14061;
  function [0:0] mux_14061(input [0:0] sel);
    case (sel) 0: mux_14061 = 1'h0; 1: mux_14061 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14062;
  function [0:0] mux_14062(input [0:0] sel);
    case (sel) 0: mux_14062 = 1'h0; 1: mux_14062 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14063;
  wire [0:0] v_14064;
  wire [0:0] v_14065;
  wire [0:0] v_14066;
  wire [0:0] v_14067;
  wire [0:0] v_14068;
  wire [0:0] v_14069;
  function [0:0] mux_14069(input [0:0] sel);
    case (sel) 0: mux_14069 = 1'h0; 1: mux_14069 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14070;
  function [0:0] mux_14070(input [0:0] sel);
    case (sel) 0: mux_14070 = 1'h0; 1: mux_14070 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14071;
  wire [0:0] v_14072;
  wire [0:0] v_14073;
  wire [0:0] v_14074;
  function [0:0] mux_14074(input [0:0] sel);
    case (sel) 0: mux_14074 = 1'h0; 1: mux_14074 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14075;
  function [0:0] mux_14075(input [0:0] sel);
    case (sel) 0: mux_14075 = 1'h0; 1: mux_14075 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14076;
  wire [0:0] v_14077;
  wire [0:0] v_14078;
  wire [0:0] v_14079;
  wire [0:0] v_14080;
  wire [0:0] v_14081;
  function [0:0] mux_14081(input [0:0] sel);
    case (sel) 0: mux_14081 = 1'h0; 1: mux_14081 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14082;
  wire [0:0] v_14083;
  wire [0:0] v_14084;
  wire [0:0] v_14085;
  wire [0:0] v_14086;
  function [0:0] mux_14086(input [0:0] sel);
    case (sel) 0: mux_14086 = 1'h0; 1: mux_14086 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14087;
  wire [0:0] v_14088;
  wire [0:0] v_14089;
  wire [0:0] v_14090;
  function [0:0] mux_14090(input [0:0] sel);
    case (sel) 0: mux_14090 = 1'h0; 1: mux_14090 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14091;
  function [0:0] mux_14091(input [0:0] sel);
    case (sel) 0: mux_14091 = 1'h0; 1: mux_14091 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_14092 = 1'h0;
  wire [0:0] v_14093;
  wire [0:0] v_14094;
  wire [0:0] act_14095;
  wire [0:0] v_14096;
  wire [0:0] v_14097;
  wire [0:0] v_14098;
  reg [0:0] v_14099 = 1'h0;
  wire [0:0] v_14100;
  wire [0:0] v_14101;
  wire [0:0] act_14102;
  wire [0:0] v_14103;
  wire [0:0] v_14104;
  wire [0:0] v_14105;
  wire [0:0] vin0_consume_en_14106;
  wire [0:0] vout_canPeek_14106;
  wire [7:0] vout_peek_14106;
  wire [0:0] v_14107;
  wire [0:0] v_14108;
  function [0:0] mux_14108(input [0:0] sel);
    case (sel) 0: mux_14108 = 1'h0; 1: mux_14108 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14109;
  wire [0:0] v_14110;
  wire [0:0] v_14111;
  wire [0:0] v_14112;
  wire [0:0] v_14113;
  function [0:0] mux_14113(input [0:0] sel);
    case (sel) 0: mux_14113 = 1'h0; 1: mux_14113 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14114;
  wire [0:0] vin0_consume_en_14115;
  wire [0:0] vout_canPeek_14115;
  wire [7:0] vout_peek_14115;
  wire [0:0] v_14116;
  wire [0:0] v_14117;
  function [0:0] mux_14117(input [0:0] sel);
    case (sel) 0: mux_14117 = 1'h0; 1: mux_14117 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14118;
  function [0:0] mux_14118(input [0:0] sel);
    case (sel) 0: mux_14118 = 1'h0; 1: mux_14118 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14119;
  wire [0:0] v_14120;
  wire [0:0] v_14121;
  wire [0:0] v_14122;
  wire [0:0] v_14123;
  wire [0:0] v_14124;
  wire [0:0] v_14125;
  function [0:0] mux_14125(input [0:0] sel);
    case (sel) 0: mux_14125 = 1'h0; 1: mux_14125 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14126;
  wire [0:0] v_14127;
  wire [0:0] v_14128;
  wire [0:0] v_14129;
  wire [0:0] v_14130;
  function [0:0] mux_14130(input [0:0] sel);
    case (sel) 0: mux_14130 = 1'h0; 1: mux_14130 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14131;
  wire [0:0] v_14132;
  wire [0:0] v_14133;
  wire [0:0] v_14134;
  function [0:0] mux_14134(input [0:0] sel);
    case (sel) 0: mux_14134 = 1'h0; 1: mux_14134 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14135;
  function [0:0] mux_14135(input [0:0] sel);
    case (sel) 0: mux_14135 = 1'h0; 1: mux_14135 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_14136 = 1'h0;
  wire [0:0] v_14137;
  wire [0:0] v_14138;
  wire [0:0] act_14139;
  wire [0:0] v_14140;
  wire [0:0] v_14141;
  wire [0:0] v_14142;
  wire [0:0] vin0_consume_en_14143;
  wire [0:0] vout_canPeek_14143;
  wire [7:0] vout_peek_14143;
  wire [0:0] v_14144;
  wire [0:0] v_14145;
  function [0:0] mux_14145(input [0:0] sel);
    case (sel) 0: mux_14145 = 1'h0; 1: mux_14145 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14146;
  wire [0:0] v_14147;
  wire [0:0] v_14148;
  wire [0:0] v_14149;
  wire [0:0] v_14150;
  function [0:0] mux_14150(input [0:0] sel);
    case (sel) 0: mux_14150 = 1'h0; 1: mux_14150 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14151;
  wire [0:0] vin0_consume_en_14152;
  wire [0:0] vout_canPeek_14152;
  wire [7:0] vout_peek_14152;
  wire [0:0] v_14153;
  wire [0:0] v_14154;
  function [0:0] mux_14154(input [0:0] sel);
    case (sel) 0: mux_14154 = 1'h0; 1: mux_14154 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14155;
  function [0:0] mux_14155(input [0:0] sel);
    case (sel) 0: mux_14155 = 1'h0; 1: mux_14155 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14156;
  wire [0:0] v_14157;
  wire [0:0] v_14158;
  wire [0:0] v_14159;
  wire [0:0] v_14160;
  wire [0:0] v_14161;
  wire [0:0] v_14162;
  function [0:0] mux_14162(input [0:0] sel);
    case (sel) 0: mux_14162 = 1'h0; 1: mux_14162 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14163;
  function [0:0] mux_14163(input [0:0] sel);
    case (sel) 0: mux_14163 = 1'h0; 1: mux_14163 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14164;
  wire [0:0] v_14165;
  wire [0:0] v_14166;
  wire [0:0] v_14167;
  function [0:0] mux_14167(input [0:0] sel);
    case (sel) 0: mux_14167 = 1'h0; 1: mux_14167 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14168;
  function [0:0] mux_14168(input [0:0] sel);
    case (sel) 0: mux_14168 = 1'h0; 1: mux_14168 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14169;
  wire [0:0] v_14170;
  wire [0:0] v_14171;
  wire [0:0] v_14172;
  wire [0:0] v_14173;
  wire [0:0] v_14174;
  function [0:0] mux_14174(input [0:0] sel);
    case (sel) 0: mux_14174 = 1'h0; 1: mux_14174 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14175;
  function [0:0] mux_14175(input [0:0] sel);
    case (sel) 0: mux_14175 = 1'h0; 1: mux_14175 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14176;
  wire [0:0] v_14177;
  wire [0:0] v_14178;
  wire [0:0] v_14179;
  function [0:0] mux_14179(input [0:0] sel);
    case (sel) 0: mux_14179 = 1'h0; 1: mux_14179 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14180;
  function [0:0] mux_14180(input [0:0] sel);
    case (sel) 0: mux_14180 = 1'h0; 1: mux_14180 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14181;
  wire [0:0] v_14182;
  wire [0:0] v_14183;
  wire [0:0] v_14184;
  wire [0:0] v_14185;
  wire [0:0] v_14186;
  function [0:0] mux_14186(input [0:0] sel);
    case (sel) 0: mux_14186 = 1'h0; 1: mux_14186 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14187;
  function [0:0] mux_14187(input [0:0] sel);
    case (sel) 0: mux_14187 = 1'h0; 1: mux_14187 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14188;
  wire [0:0] v_14189;
  wire [0:0] v_14190;
  wire [0:0] v_14191;
  function [0:0] mux_14191(input [0:0] sel);
    case (sel) 0: mux_14191 = 1'h0; 1: mux_14191 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14192;
  function [0:0] mux_14192(input [0:0] sel);
    case (sel) 0: mux_14192 = 1'h0; 1: mux_14192 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14193;
  wire [0:0] v_14194;
  wire [0:0] v_14195;
  wire [0:0] v_14196;
  wire [0:0] v_14197;
  wire [0:0] v_14198;
  function [0:0] mux_14198(input [0:0] sel);
    case (sel) 0: mux_14198 = 1'h0; 1: mux_14198 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14199;
  function [0:0] mux_14199(input [0:0] sel);
    case (sel) 0: mux_14199 = 1'h0; 1: mux_14199 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14200;
  wire [0:0] v_14201;
  wire [0:0] v_14202;
  wire [0:0] v_14203;
  function [0:0] mux_14203(input [0:0] sel);
    case (sel) 0: mux_14203 = 1'h0; 1: mux_14203 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14204;
  function [0:0] mux_14204(input [0:0] sel);
    case (sel) 0: mux_14204 = 1'h0; 1: mux_14204 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14205;
  wire [0:0] v_14206;
  wire [0:0] v_14207;
  wire [0:0] v_14208;
  wire [0:0] v_14209;
  wire [0:0] v_14210;
  function [0:0] mux_14210(input [0:0] sel);
    case (sel) 0: mux_14210 = 1'h0; 1: mux_14210 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14211;
  wire [0:0] v_14212;
  wire [0:0] v_14213;
  wire [0:0] v_14214;
  wire [0:0] v_14215;
  function [0:0] mux_14215(input [0:0] sel);
    case (sel) 0: mux_14215 = 1'h0; 1: mux_14215 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14216;
  wire [0:0] v_14217;
  wire [0:0] v_14218;
  wire [0:0] v_14219;
  function [0:0] mux_14219(input [0:0] sel);
    case (sel) 0: mux_14219 = 1'h0; 1: mux_14219 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14220;
  function [0:0] mux_14220(input [0:0] sel);
    case (sel) 0: mux_14220 = 1'h0; 1: mux_14220 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_14221 = 1'h0;
  wire [0:0] v_14222;
  wire [0:0] v_14223;
  wire [0:0] act_14224;
  wire [0:0] v_14225;
  wire [0:0] v_14226;
  wire [0:0] v_14227;
  reg [0:0] v_14228 = 1'h0;
  wire [0:0] v_14229;
  wire [0:0] v_14230;
  wire [0:0] act_14231;
  wire [0:0] v_14232;
  wire [0:0] v_14233;
  wire [0:0] v_14234;
  reg [0:0] v_14235 = 1'h0;
  wire [0:0] v_14236;
  wire [0:0] v_14237;
  wire [0:0] act_14238;
  wire [0:0] v_14239;
  wire [0:0] v_14240;
  wire [0:0] v_14241;
  reg [0:0] v_14242 = 1'h0;
  wire [0:0] v_14243;
  wire [0:0] v_14244;
  wire [0:0] act_14245;
  wire [0:0] v_14246;
  wire [0:0] v_14247;
  wire [0:0] v_14248;
  reg [0:0] v_14249 = 1'h0;
  wire [0:0] v_14250;
  wire [0:0] v_14251;
  wire [0:0] act_14252;
  wire [0:0] v_14253;
  wire [0:0] v_14254;
  wire [0:0] v_14255;
  wire [0:0] vin0_consume_en_14256;
  wire [0:0] vout_canPeek_14256;
  wire [7:0] vout_peek_14256;
  wire [0:0] v_14257;
  wire [0:0] v_14258;
  function [0:0] mux_14258(input [0:0] sel);
    case (sel) 0: mux_14258 = 1'h0; 1: mux_14258 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14259;
  wire [0:0] v_14260;
  wire [0:0] v_14261;
  wire [0:0] v_14262;
  wire [0:0] v_14263;
  function [0:0] mux_14263(input [0:0] sel);
    case (sel) 0: mux_14263 = 1'h0; 1: mux_14263 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14264;
  wire [0:0] vin0_consume_en_14265;
  wire [0:0] vout_canPeek_14265;
  wire [7:0] vout_peek_14265;
  wire [0:0] v_14266;
  wire [0:0] v_14267;
  function [0:0] mux_14267(input [0:0] sel);
    case (sel) 0: mux_14267 = 1'h0; 1: mux_14267 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14268;
  function [0:0] mux_14268(input [0:0] sel);
    case (sel) 0: mux_14268 = 1'h0; 1: mux_14268 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14269;
  wire [0:0] v_14270;
  wire [0:0] v_14271;
  wire [0:0] v_14272;
  wire [0:0] v_14273;
  wire [0:0] v_14274;
  wire [0:0] v_14275;
  function [0:0] mux_14275(input [0:0] sel);
    case (sel) 0: mux_14275 = 1'h0; 1: mux_14275 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14276;
  wire [0:0] v_14277;
  wire [0:0] v_14278;
  wire [0:0] v_14279;
  wire [0:0] v_14280;
  function [0:0] mux_14280(input [0:0] sel);
    case (sel) 0: mux_14280 = 1'h0; 1: mux_14280 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14281;
  wire [0:0] v_14282;
  wire [0:0] v_14283;
  wire [0:0] v_14284;
  function [0:0] mux_14284(input [0:0] sel);
    case (sel) 0: mux_14284 = 1'h0; 1: mux_14284 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14285;
  function [0:0] mux_14285(input [0:0] sel);
    case (sel) 0: mux_14285 = 1'h0; 1: mux_14285 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_14286 = 1'h0;
  wire [0:0] v_14287;
  wire [0:0] v_14288;
  wire [0:0] act_14289;
  wire [0:0] v_14290;
  wire [0:0] v_14291;
  wire [0:0] v_14292;
  wire [0:0] vin0_consume_en_14293;
  wire [0:0] vout_canPeek_14293;
  wire [7:0] vout_peek_14293;
  wire [0:0] v_14294;
  wire [0:0] v_14295;
  function [0:0] mux_14295(input [0:0] sel);
    case (sel) 0: mux_14295 = 1'h0; 1: mux_14295 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14296;
  wire [0:0] v_14297;
  wire [0:0] v_14298;
  wire [0:0] v_14299;
  wire [0:0] v_14300;
  function [0:0] mux_14300(input [0:0] sel);
    case (sel) 0: mux_14300 = 1'h0; 1: mux_14300 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14301;
  wire [0:0] vin0_consume_en_14302;
  wire [0:0] vout_canPeek_14302;
  wire [7:0] vout_peek_14302;
  wire [0:0] v_14303;
  wire [0:0] v_14304;
  function [0:0] mux_14304(input [0:0] sel);
    case (sel) 0: mux_14304 = 1'h0; 1: mux_14304 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14305;
  function [0:0] mux_14305(input [0:0] sel);
    case (sel) 0: mux_14305 = 1'h0; 1: mux_14305 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14306;
  wire [0:0] v_14307;
  wire [0:0] v_14308;
  wire [0:0] v_14309;
  wire [0:0] v_14310;
  wire [0:0] v_14311;
  wire [0:0] v_14312;
  function [0:0] mux_14312(input [0:0] sel);
    case (sel) 0: mux_14312 = 1'h0; 1: mux_14312 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14313;
  function [0:0] mux_14313(input [0:0] sel);
    case (sel) 0: mux_14313 = 1'h0; 1: mux_14313 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14314;
  wire [0:0] v_14315;
  wire [0:0] v_14316;
  wire [0:0] v_14317;
  function [0:0] mux_14317(input [0:0] sel);
    case (sel) 0: mux_14317 = 1'h0; 1: mux_14317 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14318;
  function [0:0] mux_14318(input [0:0] sel);
    case (sel) 0: mux_14318 = 1'h0; 1: mux_14318 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14319;
  wire [0:0] v_14320;
  wire [0:0] v_14321;
  wire [0:0] v_14322;
  wire [0:0] v_14323;
  wire [0:0] v_14324;
  function [0:0] mux_14324(input [0:0] sel);
    case (sel) 0: mux_14324 = 1'h0; 1: mux_14324 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14325;
  wire [0:0] v_14326;
  wire [0:0] v_14327;
  wire [0:0] v_14328;
  wire [0:0] v_14329;
  function [0:0] mux_14329(input [0:0] sel);
    case (sel) 0: mux_14329 = 1'h0; 1: mux_14329 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14330;
  wire [0:0] v_14331;
  wire [0:0] v_14332;
  wire [0:0] v_14333;
  function [0:0] mux_14333(input [0:0] sel);
    case (sel) 0: mux_14333 = 1'h0; 1: mux_14333 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14334;
  function [0:0] mux_14334(input [0:0] sel);
    case (sel) 0: mux_14334 = 1'h0; 1: mux_14334 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_14335 = 1'h0;
  wire [0:0] v_14336;
  wire [0:0] v_14337;
  wire [0:0] act_14338;
  wire [0:0] v_14339;
  wire [0:0] v_14340;
  wire [0:0] v_14341;
  reg [0:0] v_14342 = 1'h0;
  wire [0:0] v_14343;
  wire [0:0] v_14344;
  wire [0:0] act_14345;
  wire [0:0] v_14346;
  wire [0:0] v_14347;
  wire [0:0] v_14348;
  wire [0:0] vin0_consume_en_14349;
  wire [0:0] vout_canPeek_14349;
  wire [7:0] vout_peek_14349;
  wire [0:0] v_14350;
  wire [0:0] v_14351;
  function [0:0] mux_14351(input [0:0] sel);
    case (sel) 0: mux_14351 = 1'h0; 1: mux_14351 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14352;
  wire [0:0] v_14353;
  wire [0:0] v_14354;
  wire [0:0] v_14355;
  wire [0:0] v_14356;
  function [0:0] mux_14356(input [0:0] sel);
    case (sel) 0: mux_14356 = 1'h0; 1: mux_14356 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14357;
  wire [0:0] vin0_consume_en_14358;
  wire [0:0] vout_canPeek_14358;
  wire [7:0] vout_peek_14358;
  wire [0:0] v_14359;
  wire [0:0] v_14360;
  function [0:0] mux_14360(input [0:0] sel);
    case (sel) 0: mux_14360 = 1'h0; 1: mux_14360 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14361;
  function [0:0] mux_14361(input [0:0] sel);
    case (sel) 0: mux_14361 = 1'h0; 1: mux_14361 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14362;
  wire [0:0] v_14363;
  wire [0:0] v_14364;
  wire [0:0] v_14365;
  wire [0:0] v_14366;
  wire [0:0] v_14367;
  wire [0:0] v_14368;
  function [0:0] mux_14368(input [0:0] sel);
    case (sel) 0: mux_14368 = 1'h0; 1: mux_14368 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14369;
  wire [0:0] v_14370;
  wire [0:0] v_14371;
  wire [0:0] v_14372;
  wire [0:0] v_14373;
  function [0:0] mux_14373(input [0:0] sel);
    case (sel) 0: mux_14373 = 1'h0; 1: mux_14373 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14374;
  wire [0:0] v_14375;
  wire [0:0] v_14376;
  wire [0:0] v_14377;
  function [0:0] mux_14377(input [0:0] sel);
    case (sel) 0: mux_14377 = 1'h0; 1: mux_14377 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14378;
  function [0:0] mux_14378(input [0:0] sel);
    case (sel) 0: mux_14378 = 1'h0; 1: mux_14378 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_14379 = 1'h0;
  wire [0:0] v_14380;
  wire [0:0] v_14381;
  wire [0:0] act_14382;
  wire [0:0] v_14383;
  wire [0:0] v_14384;
  wire [0:0] v_14385;
  wire [0:0] vin0_consume_en_14386;
  wire [0:0] vout_canPeek_14386;
  wire [7:0] vout_peek_14386;
  wire [0:0] v_14387;
  wire [0:0] v_14388;
  function [0:0] mux_14388(input [0:0] sel);
    case (sel) 0: mux_14388 = 1'h0; 1: mux_14388 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14389;
  wire [0:0] v_14390;
  wire [0:0] v_14391;
  wire [0:0] v_14392;
  wire [0:0] v_14393;
  function [0:0] mux_14393(input [0:0] sel);
    case (sel) 0: mux_14393 = 1'h0; 1: mux_14393 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14394;
  wire [0:0] vin0_consume_en_14395;
  wire [0:0] vout_canPeek_14395;
  wire [7:0] vout_peek_14395;
  wire [0:0] v_14396;
  wire [0:0] v_14397;
  function [0:0] mux_14397(input [0:0] sel);
    case (sel) 0: mux_14397 = 1'h0; 1: mux_14397 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14398;
  function [0:0] mux_14398(input [0:0] sel);
    case (sel) 0: mux_14398 = 1'h0; 1: mux_14398 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14399;
  wire [0:0] v_14400;
  wire [0:0] v_14401;
  wire [0:0] v_14402;
  wire [0:0] v_14403;
  wire [0:0] v_14404;
  wire [0:0] v_14405;
  function [0:0] mux_14405(input [0:0] sel);
    case (sel) 0: mux_14405 = 1'h0; 1: mux_14405 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14406;
  function [0:0] mux_14406(input [0:0] sel);
    case (sel) 0: mux_14406 = 1'h0; 1: mux_14406 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14407;
  wire [0:0] v_14408;
  wire [0:0] v_14409;
  wire [0:0] v_14410;
  function [0:0] mux_14410(input [0:0] sel);
    case (sel) 0: mux_14410 = 1'h0; 1: mux_14410 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14411;
  function [0:0] mux_14411(input [0:0] sel);
    case (sel) 0: mux_14411 = 1'h0; 1: mux_14411 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14412;
  wire [0:0] v_14413;
  wire [0:0] v_14414;
  wire [0:0] v_14415;
  wire [0:0] v_14416;
  wire [0:0] v_14417;
  function [0:0] mux_14417(input [0:0] sel);
    case (sel) 0: mux_14417 = 1'h0; 1: mux_14417 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14418;
  function [0:0] mux_14418(input [0:0] sel);
    case (sel) 0: mux_14418 = 1'h0; 1: mux_14418 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14419;
  wire [0:0] v_14420;
  wire [0:0] v_14421;
  wire [0:0] v_14422;
  function [0:0] mux_14422(input [0:0] sel);
    case (sel) 0: mux_14422 = 1'h0; 1: mux_14422 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14423;
  function [0:0] mux_14423(input [0:0] sel);
    case (sel) 0: mux_14423 = 1'h0; 1: mux_14423 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14424;
  wire [0:0] v_14425;
  wire [0:0] v_14426;
  wire [0:0] v_14427;
  wire [0:0] v_14428;
  wire [0:0] v_14429;
  function [0:0] mux_14429(input [0:0] sel);
    case (sel) 0: mux_14429 = 1'h0; 1: mux_14429 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14430;
  wire [0:0] v_14431;
  wire [0:0] v_14432;
  wire [0:0] v_14433;
  wire [0:0] v_14434;
  function [0:0] mux_14434(input [0:0] sel);
    case (sel) 0: mux_14434 = 1'h0; 1: mux_14434 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14435;
  wire [0:0] v_14436;
  wire [0:0] v_14437;
  wire [0:0] v_14438;
  function [0:0] mux_14438(input [0:0] sel);
    case (sel) 0: mux_14438 = 1'h0; 1: mux_14438 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14439;
  function [0:0] mux_14439(input [0:0] sel);
    case (sel) 0: mux_14439 = 1'h0; 1: mux_14439 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_14440 = 1'h0;
  wire [0:0] v_14441;
  wire [0:0] v_14442;
  wire [0:0] act_14443;
  wire [0:0] v_14444;
  wire [0:0] v_14445;
  wire [0:0] v_14446;
  reg [0:0] v_14447 = 1'h0;
  wire [0:0] v_14448;
  wire [0:0] v_14449;
  wire [0:0] act_14450;
  wire [0:0] v_14451;
  wire [0:0] v_14452;
  wire [0:0] v_14453;
  reg [0:0] v_14454 = 1'h0;
  wire [0:0] v_14455;
  wire [0:0] v_14456;
  wire [0:0] act_14457;
  wire [0:0] v_14458;
  wire [0:0] v_14459;
  wire [0:0] v_14460;
  wire [0:0] vin0_consume_en_14461;
  wire [0:0] vout_canPeek_14461;
  wire [7:0] vout_peek_14461;
  wire [0:0] v_14462;
  wire [0:0] v_14463;
  function [0:0] mux_14463(input [0:0] sel);
    case (sel) 0: mux_14463 = 1'h0; 1: mux_14463 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14464;
  wire [0:0] v_14465;
  wire [0:0] v_14466;
  wire [0:0] v_14467;
  wire [0:0] v_14468;
  function [0:0] mux_14468(input [0:0] sel);
    case (sel) 0: mux_14468 = 1'h0; 1: mux_14468 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14469;
  wire [0:0] vin0_consume_en_14470;
  wire [0:0] vout_canPeek_14470;
  wire [7:0] vout_peek_14470;
  wire [0:0] v_14471;
  wire [0:0] v_14472;
  function [0:0] mux_14472(input [0:0] sel);
    case (sel) 0: mux_14472 = 1'h0; 1: mux_14472 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14473;
  function [0:0] mux_14473(input [0:0] sel);
    case (sel) 0: mux_14473 = 1'h0; 1: mux_14473 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14474;
  wire [0:0] v_14475;
  wire [0:0] v_14476;
  wire [0:0] v_14477;
  wire [0:0] v_14478;
  wire [0:0] v_14479;
  wire [0:0] v_14480;
  function [0:0] mux_14480(input [0:0] sel);
    case (sel) 0: mux_14480 = 1'h0; 1: mux_14480 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14481;
  wire [0:0] v_14482;
  wire [0:0] v_14483;
  wire [0:0] v_14484;
  wire [0:0] v_14485;
  function [0:0] mux_14485(input [0:0] sel);
    case (sel) 0: mux_14485 = 1'h0; 1: mux_14485 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14486;
  wire [0:0] v_14487;
  wire [0:0] v_14488;
  wire [0:0] v_14489;
  function [0:0] mux_14489(input [0:0] sel);
    case (sel) 0: mux_14489 = 1'h0; 1: mux_14489 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14490;
  function [0:0] mux_14490(input [0:0] sel);
    case (sel) 0: mux_14490 = 1'h0; 1: mux_14490 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_14491 = 1'h0;
  wire [0:0] v_14492;
  wire [0:0] v_14493;
  wire [0:0] act_14494;
  wire [0:0] v_14495;
  wire [0:0] v_14496;
  wire [0:0] v_14497;
  wire [0:0] vin0_consume_en_14498;
  wire [0:0] vout_canPeek_14498;
  wire [7:0] vout_peek_14498;
  wire [0:0] v_14499;
  wire [0:0] v_14500;
  function [0:0] mux_14500(input [0:0] sel);
    case (sel) 0: mux_14500 = 1'h0; 1: mux_14500 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14501;
  wire [0:0] v_14502;
  wire [0:0] v_14503;
  wire [0:0] v_14504;
  wire [0:0] v_14505;
  function [0:0] mux_14505(input [0:0] sel);
    case (sel) 0: mux_14505 = 1'h0; 1: mux_14505 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14506;
  wire [0:0] vin0_consume_en_14507;
  wire [0:0] vout_canPeek_14507;
  wire [7:0] vout_peek_14507;
  wire [0:0] v_14508;
  wire [0:0] v_14509;
  function [0:0] mux_14509(input [0:0] sel);
    case (sel) 0: mux_14509 = 1'h0; 1: mux_14509 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14510;
  function [0:0] mux_14510(input [0:0] sel);
    case (sel) 0: mux_14510 = 1'h0; 1: mux_14510 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14511;
  wire [0:0] v_14512;
  wire [0:0] v_14513;
  wire [0:0] v_14514;
  wire [0:0] v_14515;
  wire [0:0] v_14516;
  wire [0:0] v_14517;
  function [0:0] mux_14517(input [0:0] sel);
    case (sel) 0: mux_14517 = 1'h0; 1: mux_14517 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14518;
  function [0:0] mux_14518(input [0:0] sel);
    case (sel) 0: mux_14518 = 1'h0; 1: mux_14518 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14519;
  wire [0:0] v_14520;
  wire [0:0] v_14521;
  wire [0:0] v_14522;
  function [0:0] mux_14522(input [0:0] sel);
    case (sel) 0: mux_14522 = 1'h0; 1: mux_14522 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14523;
  function [0:0] mux_14523(input [0:0] sel);
    case (sel) 0: mux_14523 = 1'h0; 1: mux_14523 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14524;
  wire [0:0] v_14525;
  wire [0:0] v_14526;
  wire [0:0] v_14527;
  wire [0:0] v_14528;
  wire [0:0] v_14529;
  function [0:0] mux_14529(input [0:0] sel);
    case (sel) 0: mux_14529 = 1'h0; 1: mux_14529 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14530;
  wire [0:0] v_14531;
  wire [0:0] v_14532;
  wire [0:0] v_14533;
  wire [0:0] v_14534;
  function [0:0] mux_14534(input [0:0] sel);
    case (sel) 0: mux_14534 = 1'h0; 1: mux_14534 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14535;
  wire [0:0] v_14536;
  wire [0:0] v_14537;
  wire [0:0] v_14538;
  function [0:0] mux_14538(input [0:0] sel);
    case (sel) 0: mux_14538 = 1'h0; 1: mux_14538 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14539;
  function [0:0] mux_14539(input [0:0] sel);
    case (sel) 0: mux_14539 = 1'h0; 1: mux_14539 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_14540 = 1'h0;
  wire [0:0] v_14541;
  wire [0:0] v_14542;
  wire [0:0] act_14543;
  wire [0:0] v_14544;
  wire [0:0] v_14545;
  wire [0:0] v_14546;
  reg [0:0] v_14547 = 1'h0;
  wire [0:0] v_14548;
  wire [0:0] v_14549;
  wire [0:0] act_14550;
  wire [0:0] v_14551;
  wire [0:0] v_14552;
  wire [0:0] v_14553;
  wire [0:0] vin0_consume_en_14554;
  wire [0:0] vout_canPeek_14554;
  wire [7:0] vout_peek_14554;
  wire [0:0] v_14555;
  wire [0:0] v_14556;
  function [0:0] mux_14556(input [0:0] sel);
    case (sel) 0: mux_14556 = 1'h0; 1: mux_14556 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14557;
  wire [0:0] v_14558;
  wire [0:0] v_14559;
  wire [0:0] v_14560;
  wire [0:0] v_14561;
  function [0:0] mux_14561(input [0:0] sel);
    case (sel) 0: mux_14561 = 1'h0; 1: mux_14561 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14562;
  wire [0:0] vin0_consume_en_14563;
  wire [0:0] vout_canPeek_14563;
  wire [7:0] vout_peek_14563;
  wire [0:0] v_14564;
  wire [0:0] v_14565;
  function [0:0] mux_14565(input [0:0] sel);
    case (sel) 0: mux_14565 = 1'h0; 1: mux_14565 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14566;
  function [0:0] mux_14566(input [0:0] sel);
    case (sel) 0: mux_14566 = 1'h0; 1: mux_14566 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14567;
  wire [0:0] v_14568;
  wire [0:0] v_14569;
  wire [0:0] v_14570;
  wire [0:0] v_14571;
  wire [0:0] v_14572;
  wire [0:0] v_14573;
  function [0:0] mux_14573(input [0:0] sel);
    case (sel) 0: mux_14573 = 1'h0; 1: mux_14573 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14574;
  wire [0:0] v_14575;
  wire [0:0] v_14576;
  wire [0:0] v_14577;
  wire [0:0] v_14578;
  function [0:0] mux_14578(input [0:0] sel);
    case (sel) 0: mux_14578 = 1'h0; 1: mux_14578 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14579;
  wire [0:0] v_14580;
  wire [0:0] v_14581;
  wire [0:0] v_14582;
  function [0:0] mux_14582(input [0:0] sel);
    case (sel) 0: mux_14582 = 1'h0; 1: mux_14582 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14583;
  function [0:0] mux_14583(input [0:0] sel);
    case (sel) 0: mux_14583 = 1'h0; 1: mux_14583 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_14584 = 1'h0;
  wire [0:0] v_14585;
  wire [0:0] v_14586;
  wire [0:0] act_14587;
  wire [0:0] v_14588;
  wire [0:0] v_14589;
  wire [0:0] v_14590;
  wire [0:0] vin0_consume_en_14591;
  wire [0:0] vout_canPeek_14591;
  wire [7:0] vout_peek_14591;
  wire [0:0] v_14592;
  wire [0:0] v_14593;
  function [0:0] mux_14593(input [0:0] sel);
    case (sel) 0: mux_14593 = 1'h0; 1: mux_14593 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14594;
  wire [0:0] v_14595;
  wire [0:0] v_14596;
  wire [0:0] v_14597;
  wire [0:0] v_14598;
  function [0:0] mux_14598(input [0:0] sel);
    case (sel) 0: mux_14598 = 1'h0; 1: mux_14598 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14599;
  wire [0:0] vin0_consume_en_14600;
  wire [0:0] vout_canPeek_14600;
  wire [7:0] vout_peek_14600;
  wire [0:0] v_14601;
  wire [0:0] v_14602;
  function [0:0] mux_14602(input [0:0] sel);
    case (sel) 0: mux_14602 = 1'h0; 1: mux_14602 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14603;
  function [0:0] mux_14603(input [0:0] sel);
    case (sel) 0: mux_14603 = 1'h0; 1: mux_14603 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14604;
  wire [0:0] v_14605;
  wire [0:0] v_14606;
  wire [0:0] v_14607;
  wire [0:0] v_14608;
  wire [0:0] v_14609;
  wire [0:0] v_14610;
  function [0:0] mux_14610(input [0:0] sel);
    case (sel) 0: mux_14610 = 1'h0; 1: mux_14610 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14611;
  function [0:0] mux_14611(input [0:0] sel);
    case (sel) 0: mux_14611 = 1'h0; 1: mux_14611 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14612;
  wire [0:0] v_14613;
  wire [0:0] v_14614;
  wire [0:0] v_14615;
  function [0:0] mux_14615(input [0:0] sel);
    case (sel) 0: mux_14615 = 1'h0; 1: mux_14615 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14616;
  function [0:0] mux_14616(input [0:0] sel);
    case (sel) 0: mux_14616 = 1'h0; 1: mux_14616 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14617;
  wire [0:0] v_14618;
  wire [0:0] v_14619;
  wire [0:0] v_14620;
  wire [0:0] v_14621;
  wire [0:0] v_14622;
  function [0:0] mux_14622(input [0:0] sel);
    case (sel) 0: mux_14622 = 1'h0; 1: mux_14622 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14623;
  function [0:0] mux_14623(input [0:0] sel);
    case (sel) 0: mux_14623 = 1'h0; 1: mux_14623 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14624;
  wire [0:0] v_14625;
  wire [0:0] v_14626;
  wire [0:0] v_14627;
  function [0:0] mux_14627(input [0:0] sel);
    case (sel) 0: mux_14627 = 1'h0; 1: mux_14627 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14628;
  function [0:0] mux_14628(input [0:0] sel);
    case (sel) 0: mux_14628 = 1'h0; 1: mux_14628 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14629;
  wire [0:0] v_14630;
  wire [0:0] v_14631;
  wire [0:0] v_14632;
  wire [0:0] v_14633;
  wire [0:0] v_14634;
  function [0:0] mux_14634(input [0:0] sel);
    case (sel) 0: mux_14634 = 1'h0; 1: mux_14634 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14635;
  function [0:0] mux_14635(input [0:0] sel);
    case (sel) 0: mux_14635 = 1'h0; 1: mux_14635 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14636;
  wire [0:0] v_14637;
  wire [0:0] v_14638;
  wire [0:0] v_14639;
  function [0:0] mux_14639(input [0:0] sel);
    case (sel) 0: mux_14639 = 1'h0; 1: mux_14639 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14640;
  function [0:0] mux_14640(input [0:0] sel);
    case (sel) 0: mux_14640 = 1'h0; 1: mux_14640 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14641;
  wire [0:0] v_14642;
  wire [0:0] v_14643;
  wire [0:0] v_14644;
  wire [0:0] v_14645;
  wire [0:0] v_14646;
  function [0:0] mux_14646(input [0:0] sel);
    case (sel) 0: mux_14646 = 1'h0; 1: mux_14646 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14647;
  wire [0:0] v_14648;
  wire [0:0] v_14649;
  wire [0:0] v_14650;
  wire [0:0] v_14651;
  function [0:0] mux_14651(input [0:0] sel);
    case (sel) 0: mux_14651 = 1'h0; 1: mux_14651 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14652;
  wire [0:0] v_14653;
  wire [0:0] v_14654;
  wire [0:0] v_14655;
  function [0:0] mux_14655(input [0:0] sel);
    case (sel) 0: mux_14655 = 1'h0; 1: mux_14655 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14656;
  function [0:0] mux_14656(input [0:0] sel);
    case (sel) 0: mux_14656 = 1'h0; 1: mux_14656 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_14657 = 1'h0;
  wire [0:0] v_14658;
  wire [0:0] v_14659;
  wire [0:0] act_14660;
  wire [0:0] v_14661;
  wire [0:0] v_14662;
  wire [0:0] v_14663;
  reg [0:0] v_14664 = 1'h0;
  wire [0:0] v_14665;
  wire [0:0] v_14666;
  wire [0:0] act_14667;
  wire [0:0] v_14668;
  wire [0:0] v_14669;
  wire [0:0] v_14670;
  reg [0:0] v_14671 = 1'h0;
  wire [0:0] v_14672;
  wire [0:0] v_14673;
  wire [0:0] act_14674;
  wire [0:0] v_14675;
  wire [0:0] v_14676;
  wire [0:0] v_14677;
  reg [0:0] v_14678 = 1'h0;
  wire [0:0] v_14679;
  wire [0:0] v_14680;
  wire [0:0] act_14681;
  wire [0:0] v_14682;
  wire [0:0] v_14683;
  wire [0:0] v_14684;
  wire [0:0] vin0_consume_en_14685;
  wire [0:0] vout_canPeek_14685;
  wire [7:0] vout_peek_14685;
  wire [0:0] v_14686;
  wire [0:0] v_14687;
  function [0:0] mux_14687(input [0:0] sel);
    case (sel) 0: mux_14687 = 1'h0; 1: mux_14687 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14688;
  wire [0:0] v_14689;
  wire [0:0] v_14690;
  wire [0:0] v_14691;
  wire [0:0] v_14692;
  function [0:0] mux_14692(input [0:0] sel);
    case (sel) 0: mux_14692 = 1'h0; 1: mux_14692 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14693;
  wire [0:0] vin0_consume_en_14694;
  wire [0:0] vout_canPeek_14694;
  wire [7:0] vout_peek_14694;
  wire [0:0] v_14695;
  wire [0:0] v_14696;
  function [0:0] mux_14696(input [0:0] sel);
    case (sel) 0: mux_14696 = 1'h0; 1: mux_14696 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14697;
  function [0:0] mux_14697(input [0:0] sel);
    case (sel) 0: mux_14697 = 1'h0; 1: mux_14697 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14698;
  wire [0:0] v_14699;
  wire [0:0] v_14700;
  wire [0:0] v_14701;
  wire [0:0] v_14702;
  wire [0:0] v_14703;
  wire [0:0] v_14704;
  function [0:0] mux_14704(input [0:0] sel);
    case (sel) 0: mux_14704 = 1'h0; 1: mux_14704 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14705;
  wire [0:0] v_14706;
  wire [0:0] v_14707;
  wire [0:0] v_14708;
  wire [0:0] v_14709;
  function [0:0] mux_14709(input [0:0] sel);
    case (sel) 0: mux_14709 = 1'h0; 1: mux_14709 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14710;
  wire [0:0] v_14711;
  wire [0:0] v_14712;
  wire [0:0] v_14713;
  function [0:0] mux_14713(input [0:0] sel);
    case (sel) 0: mux_14713 = 1'h0; 1: mux_14713 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14714;
  function [0:0] mux_14714(input [0:0] sel);
    case (sel) 0: mux_14714 = 1'h0; 1: mux_14714 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_14715 = 1'h0;
  wire [0:0] v_14716;
  wire [0:0] v_14717;
  wire [0:0] act_14718;
  wire [0:0] v_14719;
  wire [0:0] v_14720;
  wire [0:0] v_14721;
  wire [0:0] vin0_consume_en_14722;
  wire [0:0] vout_canPeek_14722;
  wire [7:0] vout_peek_14722;
  wire [0:0] v_14723;
  wire [0:0] v_14724;
  function [0:0] mux_14724(input [0:0] sel);
    case (sel) 0: mux_14724 = 1'h0; 1: mux_14724 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14725;
  wire [0:0] v_14726;
  wire [0:0] v_14727;
  wire [0:0] v_14728;
  wire [0:0] v_14729;
  function [0:0] mux_14729(input [0:0] sel);
    case (sel) 0: mux_14729 = 1'h0; 1: mux_14729 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14730;
  wire [0:0] vin0_consume_en_14731;
  wire [0:0] vout_canPeek_14731;
  wire [7:0] vout_peek_14731;
  wire [0:0] v_14732;
  wire [0:0] v_14733;
  function [0:0] mux_14733(input [0:0] sel);
    case (sel) 0: mux_14733 = 1'h0; 1: mux_14733 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14734;
  function [0:0] mux_14734(input [0:0] sel);
    case (sel) 0: mux_14734 = 1'h0; 1: mux_14734 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14735;
  wire [0:0] v_14736;
  wire [0:0] v_14737;
  wire [0:0] v_14738;
  wire [0:0] v_14739;
  wire [0:0] v_14740;
  wire [0:0] v_14741;
  function [0:0] mux_14741(input [0:0] sel);
    case (sel) 0: mux_14741 = 1'h0; 1: mux_14741 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14742;
  function [0:0] mux_14742(input [0:0] sel);
    case (sel) 0: mux_14742 = 1'h0; 1: mux_14742 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14743;
  wire [0:0] v_14744;
  wire [0:0] v_14745;
  wire [0:0] v_14746;
  function [0:0] mux_14746(input [0:0] sel);
    case (sel) 0: mux_14746 = 1'h0; 1: mux_14746 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14747;
  function [0:0] mux_14747(input [0:0] sel);
    case (sel) 0: mux_14747 = 1'h0; 1: mux_14747 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14748;
  wire [0:0] v_14749;
  wire [0:0] v_14750;
  wire [0:0] v_14751;
  wire [0:0] v_14752;
  wire [0:0] v_14753;
  function [0:0] mux_14753(input [0:0] sel);
    case (sel) 0: mux_14753 = 1'h0; 1: mux_14753 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14754;
  wire [0:0] v_14755;
  wire [0:0] v_14756;
  wire [0:0] v_14757;
  wire [0:0] v_14758;
  function [0:0] mux_14758(input [0:0] sel);
    case (sel) 0: mux_14758 = 1'h0; 1: mux_14758 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14759;
  wire [0:0] v_14760;
  wire [0:0] v_14761;
  wire [0:0] v_14762;
  function [0:0] mux_14762(input [0:0] sel);
    case (sel) 0: mux_14762 = 1'h0; 1: mux_14762 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14763;
  function [0:0] mux_14763(input [0:0] sel);
    case (sel) 0: mux_14763 = 1'h0; 1: mux_14763 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_14764 = 1'h0;
  wire [0:0] v_14765;
  wire [0:0] v_14766;
  wire [0:0] act_14767;
  wire [0:0] v_14768;
  wire [0:0] v_14769;
  wire [0:0] v_14770;
  reg [0:0] v_14771 = 1'h0;
  wire [0:0] v_14772;
  wire [0:0] v_14773;
  wire [0:0] act_14774;
  wire [0:0] v_14775;
  wire [0:0] v_14776;
  wire [0:0] v_14777;
  wire [0:0] vin0_consume_en_14778;
  wire [0:0] vout_canPeek_14778;
  wire [7:0] vout_peek_14778;
  wire [0:0] v_14779;
  wire [0:0] v_14780;
  function [0:0] mux_14780(input [0:0] sel);
    case (sel) 0: mux_14780 = 1'h0; 1: mux_14780 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14781;
  wire [0:0] v_14782;
  wire [0:0] v_14783;
  wire [0:0] v_14784;
  wire [0:0] v_14785;
  function [0:0] mux_14785(input [0:0] sel);
    case (sel) 0: mux_14785 = 1'h0; 1: mux_14785 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14786;
  wire [0:0] vin0_consume_en_14787;
  wire [0:0] vout_canPeek_14787;
  wire [7:0] vout_peek_14787;
  wire [0:0] v_14788;
  wire [0:0] v_14789;
  function [0:0] mux_14789(input [0:0] sel);
    case (sel) 0: mux_14789 = 1'h0; 1: mux_14789 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14790;
  function [0:0] mux_14790(input [0:0] sel);
    case (sel) 0: mux_14790 = 1'h0; 1: mux_14790 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14791;
  wire [0:0] v_14792;
  wire [0:0] v_14793;
  wire [0:0] v_14794;
  wire [0:0] v_14795;
  wire [0:0] v_14796;
  wire [0:0] v_14797;
  function [0:0] mux_14797(input [0:0] sel);
    case (sel) 0: mux_14797 = 1'h0; 1: mux_14797 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14798;
  wire [0:0] v_14799;
  wire [0:0] v_14800;
  wire [0:0] v_14801;
  wire [0:0] v_14802;
  function [0:0] mux_14802(input [0:0] sel);
    case (sel) 0: mux_14802 = 1'h0; 1: mux_14802 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14803;
  wire [0:0] v_14804;
  wire [0:0] v_14805;
  wire [0:0] v_14806;
  function [0:0] mux_14806(input [0:0] sel);
    case (sel) 0: mux_14806 = 1'h0; 1: mux_14806 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14807;
  function [0:0] mux_14807(input [0:0] sel);
    case (sel) 0: mux_14807 = 1'h0; 1: mux_14807 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_14808 = 1'h0;
  wire [0:0] v_14809;
  wire [0:0] v_14810;
  wire [0:0] act_14811;
  wire [0:0] v_14812;
  wire [0:0] v_14813;
  wire [0:0] v_14814;
  wire [0:0] vin0_consume_en_14815;
  wire [0:0] vout_canPeek_14815;
  wire [7:0] vout_peek_14815;
  wire [0:0] v_14816;
  wire [0:0] v_14817;
  function [0:0] mux_14817(input [0:0] sel);
    case (sel) 0: mux_14817 = 1'h0; 1: mux_14817 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14818;
  wire [0:0] v_14819;
  wire [0:0] v_14820;
  wire [0:0] v_14821;
  wire [0:0] v_14822;
  function [0:0] mux_14822(input [0:0] sel);
    case (sel) 0: mux_14822 = 1'h0; 1: mux_14822 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14823;
  wire [0:0] vin0_consume_en_14824;
  wire [0:0] vout_canPeek_14824;
  wire [7:0] vout_peek_14824;
  wire [0:0] v_14825;
  wire [0:0] v_14826;
  function [0:0] mux_14826(input [0:0] sel);
    case (sel) 0: mux_14826 = 1'h0; 1: mux_14826 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14827;
  function [0:0] mux_14827(input [0:0] sel);
    case (sel) 0: mux_14827 = 1'h0; 1: mux_14827 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14828;
  wire [0:0] v_14829;
  wire [0:0] v_14830;
  wire [0:0] v_14831;
  wire [0:0] v_14832;
  wire [0:0] v_14833;
  wire [0:0] v_14834;
  function [0:0] mux_14834(input [0:0] sel);
    case (sel) 0: mux_14834 = 1'h0; 1: mux_14834 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14835;
  function [0:0] mux_14835(input [0:0] sel);
    case (sel) 0: mux_14835 = 1'h0; 1: mux_14835 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14836;
  wire [0:0] v_14837;
  wire [0:0] v_14838;
  wire [0:0] v_14839;
  function [0:0] mux_14839(input [0:0] sel);
    case (sel) 0: mux_14839 = 1'h0; 1: mux_14839 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14840;
  function [0:0] mux_14840(input [0:0] sel);
    case (sel) 0: mux_14840 = 1'h0; 1: mux_14840 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14841;
  wire [0:0] v_14842;
  wire [0:0] v_14843;
  wire [0:0] v_14844;
  wire [0:0] v_14845;
  wire [0:0] v_14846;
  function [0:0] mux_14846(input [0:0] sel);
    case (sel) 0: mux_14846 = 1'h0; 1: mux_14846 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14847;
  function [0:0] mux_14847(input [0:0] sel);
    case (sel) 0: mux_14847 = 1'h0; 1: mux_14847 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14848;
  wire [0:0] v_14849;
  wire [0:0] v_14850;
  wire [0:0] v_14851;
  function [0:0] mux_14851(input [0:0] sel);
    case (sel) 0: mux_14851 = 1'h0; 1: mux_14851 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14852;
  function [0:0] mux_14852(input [0:0] sel);
    case (sel) 0: mux_14852 = 1'h0; 1: mux_14852 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14853;
  wire [0:0] v_14854;
  wire [0:0] v_14855;
  wire [0:0] v_14856;
  wire [0:0] v_14857;
  wire [0:0] v_14858;
  function [0:0] mux_14858(input [0:0] sel);
    case (sel) 0: mux_14858 = 1'h0; 1: mux_14858 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14859;
  wire [0:0] v_14860;
  wire [0:0] v_14861;
  wire [0:0] v_14862;
  wire [0:0] v_14863;
  function [0:0] mux_14863(input [0:0] sel);
    case (sel) 0: mux_14863 = 1'h0; 1: mux_14863 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14864;
  wire [0:0] v_14865;
  wire [0:0] v_14866;
  wire [0:0] v_14867;
  function [0:0] mux_14867(input [0:0] sel);
    case (sel) 0: mux_14867 = 1'h0; 1: mux_14867 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14868;
  function [0:0] mux_14868(input [0:0] sel);
    case (sel) 0: mux_14868 = 1'h0; 1: mux_14868 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_14869 = 1'h0;
  wire [0:0] v_14870;
  wire [0:0] v_14871;
  wire [0:0] act_14872;
  wire [0:0] v_14873;
  wire [0:0] v_14874;
  wire [0:0] v_14875;
  reg [0:0] v_14876 = 1'h0;
  wire [0:0] v_14877;
  wire [0:0] v_14878;
  wire [0:0] act_14879;
  wire [0:0] v_14880;
  wire [0:0] v_14881;
  wire [0:0] v_14882;
  reg [0:0] v_14883 = 1'h0;
  wire [0:0] v_14884;
  wire [0:0] v_14885;
  wire [0:0] act_14886;
  wire [0:0] v_14887;
  wire [0:0] v_14888;
  wire [0:0] v_14889;
  wire [0:0] vin0_consume_en_14890;
  wire [0:0] vout_canPeek_14890;
  wire [7:0] vout_peek_14890;
  wire [0:0] v_14891;
  wire [0:0] v_14892;
  function [0:0] mux_14892(input [0:0] sel);
    case (sel) 0: mux_14892 = 1'h0; 1: mux_14892 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14893;
  wire [0:0] v_14894;
  wire [0:0] v_14895;
  wire [0:0] v_14896;
  wire [0:0] v_14897;
  function [0:0] mux_14897(input [0:0] sel);
    case (sel) 0: mux_14897 = 1'h0; 1: mux_14897 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14898;
  wire [0:0] vin0_consume_en_14899;
  wire [0:0] vout_canPeek_14899;
  wire [7:0] vout_peek_14899;
  wire [0:0] v_14900;
  wire [0:0] v_14901;
  function [0:0] mux_14901(input [0:0] sel);
    case (sel) 0: mux_14901 = 1'h0; 1: mux_14901 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14902;
  function [0:0] mux_14902(input [0:0] sel);
    case (sel) 0: mux_14902 = 1'h0; 1: mux_14902 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14903;
  wire [0:0] v_14904;
  wire [0:0] v_14905;
  wire [0:0] v_14906;
  wire [0:0] v_14907;
  wire [0:0] v_14908;
  wire [0:0] v_14909;
  function [0:0] mux_14909(input [0:0] sel);
    case (sel) 0: mux_14909 = 1'h0; 1: mux_14909 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14910;
  wire [0:0] v_14911;
  wire [0:0] v_14912;
  wire [0:0] v_14913;
  wire [0:0] v_14914;
  function [0:0] mux_14914(input [0:0] sel);
    case (sel) 0: mux_14914 = 1'h0; 1: mux_14914 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14915;
  wire [0:0] v_14916;
  wire [0:0] v_14917;
  wire [0:0] v_14918;
  function [0:0] mux_14918(input [0:0] sel);
    case (sel) 0: mux_14918 = 1'h0; 1: mux_14918 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14919;
  function [0:0] mux_14919(input [0:0] sel);
    case (sel) 0: mux_14919 = 1'h0; 1: mux_14919 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_14920 = 1'h0;
  wire [0:0] v_14921;
  wire [0:0] v_14922;
  wire [0:0] act_14923;
  wire [0:0] v_14924;
  wire [0:0] v_14925;
  wire [0:0] v_14926;
  wire [0:0] vin0_consume_en_14927;
  wire [0:0] vout_canPeek_14927;
  wire [7:0] vout_peek_14927;
  wire [0:0] v_14928;
  wire [0:0] v_14929;
  function [0:0] mux_14929(input [0:0] sel);
    case (sel) 0: mux_14929 = 1'h0; 1: mux_14929 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14930;
  wire [0:0] v_14931;
  wire [0:0] v_14932;
  wire [0:0] v_14933;
  wire [0:0] v_14934;
  function [0:0] mux_14934(input [0:0] sel);
    case (sel) 0: mux_14934 = 1'h0; 1: mux_14934 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14935;
  wire [0:0] vin0_consume_en_14936;
  wire [0:0] vout_canPeek_14936;
  wire [7:0] vout_peek_14936;
  wire [0:0] v_14937;
  wire [0:0] v_14938;
  function [0:0] mux_14938(input [0:0] sel);
    case (sel) 0: mux_14938 = 1'h0; 1: mux_14938 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14939;
  function [0:0] mux_14939(input [0:0] sel);
    case (sel) 0: mux_14939 = 1'h0; 1: mux_14939 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14940;
  wire [0:0] v_14941;
  wire [0:0] v_14942;
  wire [0:0] v_14943;
  wire [0:0] v_14944;
  wire [0:0] v_14945;
  wire [0:0] v_14946;
  function [0:0] mux_14946(input [0:0] sel);
    case (sel) 0: mux_14946 = 1'h0; 1: mux_14946 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14947;
  function [0:0] mux_14947(input [0:0] sel);
    case (sel) 0: mux_14947 = 1'h0; 1: mux_14947 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14948;
  wire [0:0] v_14949;
  wire [0:0] v_14950;
  wire [0:0] v_14951;
  function [0:0] mux_14951(input [0:0] sel);
    case (sel) 0: mux_14951 = 1'h0; 1: mux_14951 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14952;
  function [0:0] mux_14952(input [0:0] sel);
    case (sel) 0: mux_14952 = 1'h0; 1: mux_14952 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14953;
  wire [0:0] v_14954;
  wire [0:0] v_14955;
  wire [0:0] v_14956;
  wire [0:0] v_14957;
  wire [0:0] v_14958;
  function [0:0] mux_14958(input [0:0] sel);
    case (sel) 0: mux_14958 = 1'h0; 1: mux_14958 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14959;
  wire [0:0] v_14960;
  wire [0:0] v_14961;
  wire [0:0] v_14962;
  wire [0:0] v_14963;
  function [0:0] mux_14963(input [0:0] sel);
    case (sel) 0: mux_14963 = 1'h0; 1: mux_14963 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14964;
  wire [0:0] v_14965;
  wire [0:0] v_14966;
  wire [0:0] v_14967;
  function [0:0] mux_14967(input [0:0] sel);
    case (sel) 0: mux_14967 = 1'h0; 1: mux_14967 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14968;
  function [0:0] mux_14968(input [0:0] sel);
    case (sel) 0: mux_14968 = 1'h0; 1: mux_14968 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_14969 = 1'h0;
  wire [0:0] v_14970;
  wire [0:0] v_14971;
  wire [0:0] act_14972;
  wire [0:0] v_14973;
  wire [0:0] v_14974;
  wire [0:0] v_14975;
  reg [0:0] v_14976 = 1'h0;
  wire [0:0] v_14977;
  wire [0:0] v_14978;
  wire [0:0] act_14979;
  wire [0:0] v_14980;
  wire [0:0] v_14981;
  wire [0:0] v_14982;
  wire [0:0] vin0_consume_en_14983;
  wire [0:0] vout_canPeek_14983;
  wire [7:0] vout_peek_14983;
  wire [0:0] v_14984;
  wire [0:0] v_14985;
  function [0:0] mux_14985(input [0:0] sel);
    case (sel) 0: mux_14985 = 1'h0; 1: mux_14985 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14986;
  wire [0:0] v_14987;
  wire [0:0] v_14988;
  wire [0:0] v_14989;
  wire [0:0] v_14990;
  function [0:0] mux_14990(input [0:0] sel);
    case (sel) 0: mux_14990 = 1'h0; 1: mux_14990 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14991;
  wire [0:0] vin0_consume_en_14992;
  wire [0:0] vout_canPeek_14992;
  wire [7:0] vout_peek_14992;
  wire [0:0] v_14993;
  wire [0:0] v_14994;
  function [0:0] mux_14994(input [0:0] sel);
    case (sel) 0: mux_14994 = 1'h0; 1: mux_14994 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_14995;
  function [0:0] mux_14995(input [0:0] sel);
    case (sel) 0: mux_14995 = 1'h0; 1: mux_14995 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_14996;
  wire [0:0] v_14997;
  wire [0:0] v_14998;
  wire [0:0] v_14999;
  wire [0:0] v_15000;
  wire [0:0] v_15001;
  wire [0:0] v_15002;
  function [0:0] mux_15002(input [0:0] sel);
    case (sel) 0: mux_15002 = 1'h0; 1: mux_15002 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15003;
  wire [0:0] v_15004;
  wire [0:0] v_15005;
  wire [0:0] v_15006;
  wire [0:0] v_15007;
  function [0:0] mux_15007(input [0:0] sel);
    case (sel) 0: mux_15007 = 1'h0; 1: mux_15007 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15008;
  wire [0:0] v_15009;
  wire [0:0] v_15010;
  wire [0:0] v_15011;
  function [0:0] mux_15011(input [0:0] sel);
    case (sel) 0: mux_15011 = 1'h0; 1: mux_15011 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15012;
  function [0:0] mux_15012(input [0:0] sel);
    case (sel) 0: mux_15012 = 1'h0; 1: mux_15012 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_15013 = 1'h0;
  wire [0:0] v_15014;
  wire [0:0] v_15015;
  wire [0:0] act_15016;
  wire [0:0] v_15017;
  wire [0:0] v_15018;
  wire [0:0] v_15019;
  wire [0:0] vin0_consume_en_15020;
  wire [0:0] vout_canPeek_15020;
  wire [7:0] vout_peek_15020;
  wire [0:0] v_15021;
  wire [0:0] v_15022;
  function [0:0] mux_15022(input [0:0] sel);
    case (sel) 0: mux_15022 = 1'h0; 1: mux_15022 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15023;
  wire [0:0] v_15024;
  wire [0:0] v_15025;
  wire [0:0] v_15026;
  wire [0:0] v_15027;
  function [0:0] mux_15027(input [0:0] sel);
    case (sel) 0: mux_15027 = 1'h0; 1: mux_15027 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15028;
  wire [0:0] vin0_consume_en_15029;
  wire [0:0] vout_canPeek_15029;
  wire [7:0] vout_peek_15029;
  wire [0:0] v_15030;
  wire [0:0] v_15031;
  function [0:0] mux_15031(input [0:0] sel);
    case (sel) 0: mux_15031 = 1'h0; 1: mux_15031 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15032;
  function [0:0] mux_15032(input [0:0] sel);
    case (sel) 0: mux_15032 = 1'h0; 1: mux_15032 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15033;
  wire [0:0] v_15034;
  wire [0:0] v_15035;
  wire [0:0] v_15036;
  wire [0:0] v_15037;
  wire [0:0] v_15038;
  wire [0:0] v_15039;
  function [0:0] mux_15039(input [0:0] sel);
    case (sel) 0: mux_15039 = 1'h0; 1: mux_15039 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15040;
  function [0:0] mux_15040(input [0:0] sel);
    case (sel) 0: mux_15040 = 1'h0; 1: mux_15040 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15041;
  wire [0:0] v_15042;
  wire [0:0] v_15043;
  wire [0:0] v_15044;
  function [0:0] mux_15044(input [0:0] sel);
    case (sel) 0: mux_15044 = 1'h0; 1: mux_15044 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15045;
  function [0:0] mux_15045(input [0:0] sel);
    case (sel) 0: mux_15045 = 1'h0; 1: mux_15045 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15046;
  wire [0:0] v_15047;
  wire [0:0] v_15048;
  wire [0:0] v_15049;
  wire [0:0] v_15050;
  wire [0:0] v_15051;
  function [0:0] mux_15051(input [0:0] sel);
    case (sel) 0: mux_15051 = 1'h0; 1: mux_15051 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15052;
  function [0:0] mux_15052(input [0:0] sel);
    case (sel) 0: mux_15052 = 1'h0; 1: mux_15052 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15053;
  wire [0:0] v_15054;
  wire [0:0] v_15055;
  wire [0:0] v_15056;
  function [0:0] mux_15056(input [0:0] sel);
    case (sel) 0: mux_15056 = 1'h0; 1: mux_15056 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15057;
  function [0:0] mux_15057(input [0:0] sel);
    case (sel) 0: mux_15057 = 1'h0; 1: mux_15057 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15058;
  wire [0:0] v_15059;
  wire [0:0] v_15060;
  wire [0:0] v_15061;
  wire [0:0] v_15062;
  wire [0:0] v_15063;
  function [0:0] mux_15063(input [0:0] sel);
    case (sel) 0: mux_15063 = 1'h0; 1: mux_15063 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15064;
  function [0:0] mux_15064(input [0:0] sel);
    case (sel) 0: mux_15064 = 1'h0; 1: mux_15064 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15065;
  wire [0:0] v_15066;
  wire [0:0] v_15067;
  wire [0:0] v_15068;
  function [0:0] mux_15068(input [0:0] sel);
    case (sel) 0: mux_15068 = 1'h0; 1: mux_15068 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15069;
  function [0:0] mux_15069(input [0:0] sel);
    case (sel) 0: mux_15069 = 1'h0; 1: mux_15069 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15070;
  wire [0:0] v_15071;
  wire [0:0] v_15072;
  wire [0:0] v_15073;
  wire [0:0] v_15074;
  wire [0:0] v_15075;
  function [0:0] mux_15075(input [0:0] sel);
    case (sel) 0: mux_15075 = 1'h0; 1: mux_15075 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15076;
  function [0:0] mux_15076(input [0:0] sel);
    case (sel) 0: mux_15076 = 1'h0; 1: mux_15076 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15077;
  wire [0:0] v_15078;
  wire [0:0] v_15079;
  wire [0:0] v_15080;
  function [0:0] mux_15080(input [0:0] sel);
    case (sel) 0: mux_15080 = 1'h0; 1: mux_15080 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15081;
  function [0:0] mux_15081(input [0:0] sel);
    case (sel) 0: mux_15081 = 1'h0; 1: mux_15081 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15082;
  wire [0:0] v_15083;
  wire [0:0] v_15084;
  wire [0:0] v_15085;
  wire [0:0] v_15086;
  wire [0:0] v_15087;
  function [0:0] mux_15087(input [0:0] sel);
    case (sel) 0: mux_15087 = 1'h0; 1: mux_15087 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15088;
  function [0:0] mux_15088(input [0:0] sel);
    case (sel) 0: mux_15088 = 1'h0; 1: mux_15088 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15089;
  wire [0:0] v_15090;
  wire [0:0] v_15091;
  wire [0:0] v_15092;
  function [0:0] mux_15092(input [0:0] sel);
    case (sel) 0: mux_15092 = 1'h0; 1: mux_15092 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15093;
  function [0:0] mux_15093(input [0:0] sel);
    case (sel) 0: mux_15093 = 1'h0; 1: mux_15093 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15094;
  wire [0:0] v_15095;
  wire [0:0] v_15096;
  wire [0:0] v_15097;
  wire [0:0] v_15098;
  wire [0:0] v_15099;
  function [0:0] mux_15099(input [0:0] sel);
    case (sel) 0: mux_15099 = 1'h0; 1: mux_15099 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15100;
  function [0:0] mux_15100(input [0:0] sel);
    case (sel) 0: mux_15100 = 1'h0; 1: mux_15100 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15101;
  wire [0:0] v_15102;
  wire [0:0] v_15103;
  wire [0:0] v_15104;
  function [0:0] mux_15104(input [0:0] sel);
    case (sel) 0: mux_15104 = 1'h0; 1: mux_15104 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15105;
  function [0:0] mux_15105(input [0:0] sel);
    case (sel) 0: mux_15105 = 1'h0; 1: mux_15105 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15106;
  wire [0:0] v_15107;
  wire [0:0] v_15108;
  wire [0:0] v_15109;
  wire [0:0] v_15110;
  wire [0:0] v_15111;
  function [0:0] mux_15111(input [0:0] sel);
    case (sel) 0: mux_15111 = 1'h0; 1: mux_15111 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15112;
  function [0:0] mux_15112(input [0:0] sel);
    case (sel) 0: mux_15112 = 1'h0; 1: mux_15112 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15113;
  wire [0:0] v_15114;
  wire [0:0] v_15115;
  wire [0:0] v_15116;
  function [0:0] mux_15116(input [0:0] sel);
    case (sel) 0: mux_15116 = 1'h0; 1: mux_15116 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15117;
  function [0:0] mux_15117(input [0:0] sel);
    case (sel) 0: mux_15117 = 1'h0; 1: mux_15117 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15118;
  wire [0:0] v_15119;
  wire [0:0] v_15120;
  wire [0:0] v_15121;
  wire [0:0] v_15122;
  wire [0:0] v_15123;
  function [0:0] mux_15123(input [0:0] sel);
    case (sel) 0: mux_15123 = 1'h0; 1: mux_15123 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15124;
  wire [0:0] v_15125;
  wire [0:0] v_15126;
  wire [0:0] v_15127;
  wire [0:0] v_15128;
  function [0:0] mux_15128(input [0:0] sel);
    case (sel) 0: mux_15128 = 1'h0; 1: mux_15128 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15129;
  wire [0:0] v_15130;
  wire [0:0] v_15131;
  wire [0:0] v_15132;
  function [0:0] mux_15132(input [0:0] sel);
    case (sel) 0: mux_15132 = 1'h0; 1: mux_15132 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15133;
  function [0:0] mux_15133(input [0:0] sel);
    case (sel) 0: mux_15133 = 1'h0; 1: mux_15133 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_15134 = 1'h0;
  wire [0:0] v_15135;
  wire [0:0] v_15136;
  wire [0:0] act_15137;
  wire [0:0] v_15138;
  wire [0:0] v_15139;
  wire [0:0] v_15140;
  reg [0:0] v_15141 = 1'h0;
  wire [0:0] v_15142;
  wire [0:0] v_15143;
  wire [0:0] act_15144;
  wire [0:0] v_15145;
  wire [0:0] v_15146;
  wire [0:0] v_15147;
  reg [0:0] v_15148 = 1'h0;
  wire [0:0] v_15149;
  wire [0:0] v_15150;
  wire [0:0] act_15151;
  wire [0:0] v_15152;
  wire [0:0] v_15153;
  wire [0:0] v_15154;
  reg [0:0] v_15155 = 1'h0;
  wire [0:0] v_15156;
  wire [0:0] v_15157;
  wire [0:0] act_15158;
  wire [0:0] v_15159;
  wire [0:0] v_15160;
  wire [0:0] v_15161;
  reg [0:0] v_15162 = 1'h0;
  wire [0:0] v_15163;
  wire [0:0] v_15164;
  wire [0:0] act_15165;
  wire [0:0] v_15166;
  wire [0:0] v_15167;
  wire [0:0] v_15168;
  reg [0:0] v_15169 = 1'h0;
  wire [0:0] v_15170;
  wire [0:0] v_15171;
  wire [0:0] act_15172;
  wire [0:0] v_15173;
  wire [0:0] v_15174;
  wire [0:0] v_15175;
  reg [0:0] v_15176 = 1'h0;
  wire [0:0] v_15177;
  wire [0:0] v_15178;
  wire [0:0] act_15179;
  wire [0:0] v_15180;
  wire [0:0] v_15181;
  wire [0:0] v_15182;
  reg [0:0] v_15183 = 1'h0;
  wire [0:0] v_15184;
  wire [0:0] v_15185;
  wire [0:0] act_15186;
  wire [0:0] v_15187;
  wire [0:0] v_15188;
  wire [0:0] v_15189;
  wire [0:0] vin0_consume_en_15190;
  wire [0:0] vout_canPeek_15190;
  wire [7:0] vout_peek_15190;
  wire [0:0] v_15191;
  wire [0:0] v_15192;
  function [0:0] mux_15192(input [0:0] sel);
    case (sel) 0: mux_15192 = 1'h0; 1: mux_15192 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15193;
  wire [0:0] v_15194;
  wire [0:0] v_15195;
  wire [0:0] v_15196;
  wire [0:0] v_15197;
  function [0:0] mux_15197(input [0:0] sel);
    case (sel) 0: mux_15197 = 1'h0; 1: mux_15197 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15198;
  wire [0:0] vin0_consume_en_15199;
  wire [0:0] vout_canPeek_15199;
  wire [7:0] vout_peek_15199;
  wire [0:0] v_15200;
  wire [0:0] v_15201;
  function [0:0] mux_15201(input [0:0] sel);
    case (sel) 0: mux_15201 = 1'h0; 1: mux_15201 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15202;
  function [0:0] mux_15202(input [0:0] sel);
    case (sel) 0: mux_15202 = 1'h0; 1: mux_15202 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15203;
  wire [0:0] v_15204;
  wire [0:0] v_15205;
  wire [0:0] v_15206;
  wire [0:0] v_15207;
  wire [0:0] v_15208;
  wire [0:0] v_15209;
  function [0:0] mux_15209(input [0:0] sel);
    case (sel) 0: mux_15209 = 1'h0; 1: mux_15209 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15210;
  wire [0:0] v_15211;
  wire [0:0] v_15212;
  wire [0:0] v_15213;
  wire [0:0] v_15214;
  function [0:0] mux_15214(input [0:0] sel);
    case (sel) 0: mux_15214 = 1'h0; 1: mux_15214 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15215;
  wire [0:0] v_15216;
  wire [0:0] v_15217;
  wire [0:0] v_15218;
  function [0:0] mux_15218(input [0:0] sel);
    case (sel) 0: mux_15218 = 1'h0; 1: mux_15218 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15219;
  function [0:0] mux_15219(input [0:0] sel);
    case (sel) 0: mux_15219 = 1'h0; 1: mux_15219 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_15220 = 1'h0;
  wire [0:0] v_15221;
  wire [0:0] v_15222;
  wire [0:0] act_15223;
  wire [0:0] v_15224;
  wire [0:0] v_15225;
  wire [0:0] v_15226;
  wire [0:0] vin0_consume_en_15227;
  wire [0:0] vout_canPeek_15227;
  wire [7:0] vout_peek_15227;
  wire [0:0] v_15228;
  wire [0:0] v_15229;
  function [0:0] mux_15229(input [0:0] sel);
    case (sel) 0: mux_15229 = 1'h0; 1: mux_15229 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15230;
  wire [0:0] v_15231;
  wire [0:0] v_15232;
  wire [0:0] v_15233;
  wire [0:0] v_15234;
  function [0:0] mux_15234(input [0:0] sel);
    case (sel) 0: mux_15234 = 1'h0; 1: mux_15234 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15235;
  wire [0:0] vin0_consume_en_15236;
  wire [0:0] vout_canPeek_15236;
  wire [7:0] vout_peek_15236;
  wire [0:0] v_15237;
  wire [0:0] v_15238;
  function [0:0] mux_15238(input [0:0] sel);
    case (sel) 0: mux_15238 = 1'h0; 1: mux_15238 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15239;
  function [0:0] mux_15239(input [0:0] sel);
    case (sel) 0: mux_15239 = 1'h0; 1: mux_15239 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15240;
  wire [0:0] v_15241;
  wire [0:0] v_15242;
  wire [0:0] v_15243;
  wire [0:0] v_15244;
  wire [0:0] v_15245;
  wire [0:0] v_15246;
  function [0:0] mux_15246(input [0:0] sel);
    case (sel) 0: mux_15246 = 1'h0; 1: mux_15246 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15247;
  function [0:0] mux_15247(input [0:0] sel);
    case (sel) 0: mux_15247 = 1'h0; 1: mux_15247 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15248;
  wire [0:0] v_15249;
  wire [0:0] v_15250;
  wire [0:0] v_15251;
  function [0:0] mux_15251(input [0:0] sel);
    case (sel) 0: mux_15251 = 1'h0; 1: mux_15251 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15252;
  function [0:0] mux_15252(input [0:0] sel);
    case (sel) 0: mux_15252 = 1'h0; 1: mux_15252 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15253;
  wire [0:0] v_15254;
  wire [0:0] v_15255;
  wire [0:0] v_15256;
  wire [0:0] v_15257;
  wire [0:0] v_15258;
  function [0:0] mux_15258(input [0:0] sel);
    case (sel) 0: mux_15258 = 1'h0; 1: mux_15258 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15259;
  wire [0:0] v_15260;
  wire [0:0] v_15261;
  wire [0:0] v_15262;
  wire [0:0] v_15263;
  function [0:0] mux_15263(input [0:0] sel);
    case (sel) 0: mux_15263 = 1'h0; 1: mux_15263 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15264;
  wire [0:0] v_15265;
  wire [0:0] v_15266;
  wire [0:0] v_15267;
  function [0:0] mux_15267(input [0:0] sel);
    case (sel) 0: mux_15267 = 1'h0; 1: mux_15267 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15268;
  function [0:0] mux_15268(input [0:0] sel);
    case (sel) 0: mux_15268 = 1'h0; 1: mux_15268 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_15269 = 1'h0;
  wire [0:0] v_15270;
  wire [0:0] v_15271;
  wire [0:0] act_15272;
  wire [0:0] v_15273;
  wire [0:0] v_15274;
  wire [0:0] v_15275;
  reg [0:0] v_15276 = 1'h0;
  wire [0:0] v_15277;
  wire [0:0] v_15278;
  wire [0:0] act_15279;
  wire [0:0] v_15280;
  wire [0:0] v_15281;
  wire [0:0] v_15282;
  wire [0:0] vin0_consume_en_15283;
  wire [0:0] vout_canPeek_15283;
  wire [7:0] vout_peek_15283;
  wire [0:0] v_15284;
  wire [0:0] v_15285;
  function [0:0] mux_15285(input [0:0] sel);
    case (sel) 0: mux_15285 = 1'h0; 1: mux_15285 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15286;
  wire [0:0] v_15287;
  wire [0:0] v_15288;
  wire [0:0] v_15289;
  wire [0:0] v_15290;
  function [0:0] mux_15290(input [0:0] sel);
    case (sel) 0: mux_15290 = 1'h0; 1: mux_15290 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15291;
  wire [0:0] vin0_consume_en_15292;
  wire [0:0] vout_canPeek_15292;
  wire [7:0] vout_peek_15292;
  wire [0:0] v_15293;
  wire [0:0] v_15294;
  function [0:0] mux_15294(input [0:0] sel);
    case (sel) 0: mux_15294 = 1'h0; 1: mux_15294 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15295;
  function [0:0] mux_15295(input [0:0] sel);
    case (sel) 0: mux_15295 = 1'h0; 1: mux_15295 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15296;
  wire [0:0] v_15297;
  wire [0:0] v_15298;
  wire [0:0] v_15299;
  wire [0:0] v_15300;
  wire [0:0] v_15301;
  wire [0:0] v_15302;
  function [0:0] mux_15302(input [0:0] sel);
    case (sel) 0: mux_15302 = 1'h0; 1: mux_15302 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15303;
  wire [0:0] v_15304;
  wire [0:0] v_15305;
  wire [0:0] v_15306;
  wire [0:0] v_15307;
  function [0:0] mux_15307(input [0:0] sel);
    case (sel) 0: mux_15307 = 1'h0; 1: mux_15307 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15308;
  wire [0:0] v_15309;
  wire [0:0] v_15310;
  wire [0:0] v_15311;
  function [0:0] mux_15311(input [0:0] sel);
    case (sel) 0: mux_15311 = 1'h0; 1: mux_15311 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15312;
  function [0:0] mux_15312(input [0:0] sel);
    case (sel) 0: mux_15312 = 1'h0; 1: mux_15312 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_15313 = 1'h0;
  wire [0:0] v_15314;
  wire [0:0] v_15315;
  wire [0:0] act_15316;
  wire [0:0] v_15317;
  wire [0:0] v_15318;
  wire [0:0] v_15319;
  wire [0:0] vin0_consume_en_15320;
  wire [0:0] vout_canPeek_15320;
  wire [7:0] vout_peek_15320;
  wire [0:0] v_15321;
  wire [0:0] v_15322;
  function [0:0] mux_15322(input [0:0] sel);
    case (sel) 0: mux_15322 = 1'h0; 1: mux_15322 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15323;
  wire [0:0] v_15324;
  wire [0:0] v_15325;
  wire [0:0] v_15326;
  wire [0:0] v_15327;
  function [0:0] mux_15327(input [0:0] sel);
    case (sel) 0: mux_15327 = 1'h0; 1: mux_15327 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15328;
  wire [0:0] vin0_consume_en_15329;
  wire [0:0] vout_canPeek_15329;
  wire [7:0] vout_peek_15329;
  wire [0:0] v_15330;
  wire [0:0] v_15331;
  function [0:0] mux_15331(input [0:0] sel);
    case (sel) 0: mux_15331 = 1'h0; 1: mux_15331 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15332;
  function [0:0] mux_15332(input [0:0] sel);
    case (sel) 0: mux_15332 = 1'h0; 1: mux_15332 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15333;
  wire [0:0] v_15334;
  wire [0:0] v_15335;
  wire [0:0] v_15336;
  wire [0:0] v_15337;
  wire [0:0] v_15338;
  wire [0:0] v_15339;
  function [0:0] mux_15339(input [0:0] sel);
    case (sel) 0: mux_15339 = 1'h0; 1: mux_15339 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15340;
  function [0:0] mux_15340(input [0:0] sel);
    case (sel) 0: mux_15340 = 1'h0; 1: mux_15340 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15341;
  wire [0:0] v_15342;
  wire [0:0] v_15343;
  wire [0:0] v_15344;
  function [0:0] mux_15344(input [0:0] sel);
    case (sel) 0: mux_15344 = 1'h0; 1: mux_15344 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15345;
  function [0:0] mux_15345(input [0:0] sel);
    case (sel) 0: mux_15345 = 1'h0; 1: mux_15345 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15346;
  wire [0:0] v_15347;
  wire [0:0] v_15348;
  wire [0:0] v_15349;
  wire [0:0] v_15350;
  wire [0:0] v_15351;
  function [0:0] mux_15351(input [0:0] sel);
    case (sel) 0: mux_15351 = 1'h0; 1: mux_15351 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15352;
  function [0:0] mux_15352(input [0:0] sel);
    case (sel) 0: mux_15352 = 1'h0; 1: mux_15352 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15353;
  wire [0:0] v_15354;
  wire [0:0] v_15355;
  wire [0:0] v_15356;
  function [0:0] mux_15356(input [0:0] sel);
    case (sel) 0: mux_15356 = 1'h0; 1: mux_15356 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15357;
  function [0:0] mux_15357(input [0:0] sel);
    case (sel) 0: mux_15357 = 1'h0; 1: mux_15357 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15358;
  wire [0:0] v_15359;
  wire [0:0] v_15360;
  wire [0:0] v_15361;
  wire [0:0] v_15362;
  wire [0:0] v_15363;
  function [0:0] mux_15363(input [0:0] sel);
    case (sel) 0: mux_15363 = 1'h0; 1: mux_15363 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15364;
  wire [0:0] v_15365;
  wire [0:0] v_15366;
  wire [0:0] v_15367;
  wire [0:0] v_15368;
  function [0:0] mux_15368(input [0:0] sel);
    case (sel) 0: mux_15368 = 1'h0; 1: mux_15368 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15369;
  wire [0:0] v_15370;
  wire [0:0] v_15371;
  wire [0:0] v_15372;
  function [0:0] mux_15372(input [0:0] sel);
    case (sel) 0: mux_15372 = 1'h0; 1: mux_15372 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15373;
  function [0:0] mux_15373(input [0:0] sel);
    case (sel) 0: mux_15373 = 1'h0; 1: mux_15373 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_15374 = 1'h0;
  wire [0:0] v_15375;
  wire [0:0] v_15376;
  wire [0:0] act_15377;
  wire [0:0] v_15378;
  wire [0:0] v_15379;
  wire [0:0] v_15380;
  reg [0:0] v_15381 = 1'h0;
  wire [0:0] v_15382;
  wire [0:0] v_15383;
  wire [0:0] act_15384;
  wire [0:0] v_15385;
  wire [0:0] v_15386;
  wire [0:0] v_15387;
  reg [0:0] v_15388 = 1'h0;
  wire [0:0] v_15389;
  wire [0:0] v_15390;
  wire [0:0] act_15391;
  wire [0:0] v_15392;
  wire [0:0] v_15393;
  wire [0:0] v_15394;
  wire [0:0] vin0_consume_en_15395;
  wire [0:0] vout_canPeek_15395;
  wire [7:0] vout_peek_15395;
  wire [0:0] v_15396;
  wire [0:0] v_15397;
  function [0:0] mux_15397(input [0:0] sel);
    case (sel) 0: mux_15397 = 1'h0; 1: mux_15397 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15398;
  wire [0:0] v_15399;
  wire [0:0] v_15400;
  wire [0:0] v_15401;
  wire [0:0] v_15402;
  function [0:0] mux_15402(input [0:0] sel);
    case (sel) 0: mux_15402 = 1'h0; 1: mux_15402 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15403;
  wire [0:0] vin0_consume_en_15404;
  wire [0:0] vout_canPeek_15404;
  wire [7:0] vout_peek_15404;
  wire [0:0] v_15405;
  wire [0:0] v_15406;
  function [0:0] mux_15406(input [0:0] sel);
    case (sel) 0: mux_15406 = 1'h0; 1: mux_15406 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15407;
  function [0:0] mux_15407(input [0:0] sel);
    case (sel) 0: mux_15407 = 1'h0; 1: mux_15407 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15408;
  wire [0:0] v_15409;
  wire [0:0] v_15410;
  wire [0:0] v_15411;
  wire [0:0] v_15412;
  wire [0:0] v_15413;
  wire [0:0] v_15414;
  function [0:0] mux_15414(input [0:0] sel);
    case (sel) 0: mux_15414 = 1'h0; 1: mux_15414 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15415;
  wire [0:0] v_15416;
  wire [0:0] v_15417;
  wire [0:0] v_15418;
  wire [0:0] v_15419;
  function [0:0] mux_15419(input [0:0] sel);
    case (sel) 0: mux_15419 = 1'h0; 1: mux_15419 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15420;
  wire [0:0] v_15421;
  wire [0:0] v_15422;
  wire [0:0] v_15423;
  function [0:0] mux_15423(input [0:0] sel);
    case (sel) 0: mux_15423 = 1'h0; 1: mux_15423 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15424;
  function [0:0] mux_15424(input [0:0] sel);
    case (sel) 0: mux_15424 = 1'h0; 1: mux_15424 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_15425 = 1'h0;
  wire [0:0] v_15426;
  wire [0:0] v_15427;
  wire [0:0] act_15428;
  wire [0:0] v_15429;
  wire [0:0] v_15430;
  wire [0:0] v_15431;
  wire [0:0] vin0_consume_en_15432;
  wire [0:0] vout_canPeek_15432;
  wire [7:0] vout_peek_15432;
  wire [0:0] v_15433;
  wire [0:0] v_15434;
  function [0:0] mux_15434(input [0:0] sel);
    case (sel) 0: mux_15434 = 1'h0; 1: mux_15434 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15435;
  wire [0:0] v_15436;
  wire [0:0] v_15437;
  wire [0:0] v_15438;
  wire [0:0] v_15439;
  function [0:0] mux_15439(input [0:0] sel);
    case (sel) 0: mux_15439 = 1'h0; 1: mux_15439 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15440;
  wire [0:0] vin0_consume_en_15441;
  wire [0:0] vout_canPeek_15441;
  wire [7:0] vout_peek_15441;
  wire [0:0] v_15442;
  wire [0:0] v_15443;
  function [0:0] mux_15443(input [0:0] sel);
    case (sel) 0: mux_15443 = 1'h0; 1: mux_15443 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15444;
  function [0:0] mux_15444(input [0:0] sel);
    case (sel) 0: mux_15444 = 1'h0; 1: mux_15444 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15445;
  wire [0:0] v_15446;
  wire [0:0] v_15447;
  wire [0:0] v_15448;
  wire [0:0] v_15449;
  wire [0:0] v_15450;
  wire [0:0] v_15451;
  function [0:0] mux_15451(input [0:0] sel);
    case (sel) 0: mux_15451 = 1'h0; 1: mux_15451 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15452;
  function [0:0] mux_15452(input [0:0] sel);
    case (sel) 0: mux_15452 = 1'h0; 1: mux_15452 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15453;
  wire [0:0] v_15454;
  wire [0:0] v_15455;
  wire [0:0] v_15456;
  function [0:0] mux_15456(input [0:0] sel);
    case (sel) 0: mux_15456 = 1'h0; 1: mux_15456 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15457;
  function [0:0] mux_15457(input [0:0] sel);
    case (sel) 0: mux_15457 = 1'h0; 1: mux_15457 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15458;
  wire [0:0] v_15459;
  wire [0:0] v_15460;
  wire [0:0] v_15461;
  wire [0:0] v_15462;
  wire [0:0] v_15463;
  function [0:0] mux_15463(input [0:0] sel);
    case (sel) 0: mux_15463 = 1'h0; 1: mux_15463 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15464;
  wire [0:0] v_15465;
  wire [0:0] v_15466;
  wire [0:0] v_15467;
  wire [0:0] v_15468;
  function [0:0] mux_15468(input [0:0] sel);
    case (sel) 0: mux_15468 = 1'h0; 1: mux_15468 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15469;
  wire [0:0] v_15470;
  wire [0:0] v_15471;
  wire [0:0] v_15472;
  function [0:0] mux_15472(input [0:0] sel);
    case (sel) 0: mux_15472 = 1'h0; 1: mux_15472 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15473;
  function [0:0] mux_15473(input [0:0] sel);
    case (sel) 0: mux_15473 = 1'h0; 1: mux_15473 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_15474 = 1'h0;
  wire [0:0] v_15475;
  wire [0:0] v_15476;
  wire [0:0] act_15477;
  wire [0:0] v_15478;
  wire [0:0] v_15479;
  wire [0:0] v_15480;
  reg [0:0] v_15481 = 1'h0;
  wire [0:0] v_15482;
  wire [0:0] v_15483;
  wire [0:0] act_15484;
  wire [0:0] v_15485;
  wire [0:0] v_15486;
  wire [0:0] v_15487;
  wire [0:0] vin0_consume_en_15488;
  wire [0:0] vout_canPeek_15488;
  wire [7:0] vout_peek_15488;
  wire [0:0] v_15489;
  wire [0:0] v_15490;
  function [0:0] mux_15490(input [0:0] sel);
    case (sel) 0: mux_15490 = 1'h0; 1: mux_15490 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15491;
  wire [0:0] v_15492;
  wire [0:0] v_15493;
  wire [0:0] v_15494;
  wire [0:0] v_15495;
  function [0:0] mux_15495(input [0:0] sel);
    case (sel) 0: mux_15495 = 1'h0; 1: mux_15495 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15496;
  wire [0:0] vin0_consume_en_15497;
  wire [0:0] vout_canPeek_15497;
  wire [7:0] vout_peek_15497;
  wire [0:0] v_15498;
  wire [0:0] v_15499;
  function [0:0] mux_15499(input [0:0] sel);
    case (sel) 0: mux_15499 = 1'h0; 1: mux_15499 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15500;
  function [0:0] mux_15500(input [0:0] sel);
    case (sel) 0: mux_15500 = 1'h0; 1: mux_15500 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15501;
  wire [0:0] v_15502;
  wire [0:0] v_15503;
  wire [0:0] v_15504;
  wire [0:0] v_15505;
  wire [0:0] v_15506;
  wire [0:0] v_15507;
  function [0:0] mux_15507(input [0:0] sel);
    case (sel) 0: mux_15507 = 1'h0; 1: mux_15507 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15508;
  wire [0:0] v_15509;
  wire [0:0] v_15510;
  wire [0:0] v_15511;
  wire [0:0] v_15512;
  function [0:0] mux_15512(input [0:0] sel);
    case (sel) 0: mux_15512 = 1'h0; 1: mux_15512 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15513;
  wire [0:0] v_15514;
  wire [0:0] v_15515;
  wire [0:0] v_15516;
  function [0:0] mux_15516(input [0:0] sel);
    case (sel) 0: mux_15516 = 1'h0; 1: mux_15516 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15517;
  function [0:0] mux_15517(input [0:0] sel);
    case (sel) 0: mux_15517 = 1'h0; 1: mux_15517 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_15518 = 1'h0;
  wire [0:0] v_15519;
  wire [0:0] v_15520;
  wire [0:0] act_15521;
  wire [0:0] v_15522;
  wire [0:0] v_15523;
  wire [0:0] v_15524;
  wire [0:0] vin0_consume_en_15525;
  wire [0:0] vout_canPeek_15525;
  wire [7:0] vout_peek_15525;
  wire [0:0] v_15526;
  wire [0:0] v_15527;
  function [0:0] mux_15527(input [0:0] sel);
    case (sel) 0: mux_15527 = 1'h0; 1: mux_15527 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15528;
  wire [0:0] v_15529;
  wire [0:0] v_15530;
  wire [0:0] v_15531;
  wire [0:0] v_15532;
  function [0:0] mux_15532(input [0:0] sel);
    case (sel) 0: mux_15532 = 1'h0; 1: mux_15532 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15533;
  wire [0:0] vin0_consume_en_15534;
  wire [0:0] vout_canPeek_15534;
  wire [7:0] vout_peek_15534;
  wire [0:0] v_15535;
  wire [0:0] v_15536;
  function [0:0] mux_15536(input [0:0] sel);
    case (sel) 0: mux_15536 = 1'h0; 1: mux_15536 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15537;
  function [0:0] mux_15537(input [0:0] sel);
    case (sel) 0: mux_15537 = 1'h0; 1: mux_15537 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15538;
  wire [0:0] v_15539;
  wire [0:0] v_15540;
  wire [0:0] v_15541;
  wire [0:0] v_15542;
  wire [0:0] v_15543;
  wire [0:0] v_15544;
  function [0:0] mux_15544(input [0:0] sel);
    case (sel) 0: mux_15544 = 1'h0; 1: mux_15544 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15545;
  function [0:0] mux_15545(input [0:0] sel);
    case (sel) 0: mux_15545 = 1'h0; 1: mux_15545 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15546;
  wire [0:0] v_15547;
  wire [0:0] v_15548;
  wire [0:0] v_15549;
  function [0:0] mux_15549(input [0:0] sel);
    case (sel) 0: mux_15549 = 1'h0; 1: mux_15549 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15550;
  function [0:0] mux_15550(input [0:0] sel);
    case (sel) 0: mux_15550 = 1'h0; 1: mux_15550 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15551;
  wire [0:0] v_15552;
  wire [0:0] v_15553;
  wire [0:0] v_15554;
  wire [0:0] v_15555;
  wire [0:0] v_15556;
  function [0:0] mux_15556(input [0:0] sel);
    case (sel) 0: mux_15556 = 1'h0; 1: mux_15556 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15557;
  function [0:0] mux_15557(input [0:0] sel);
    case (sel) 0: mux_15557 = 1'h0; 1: mux_15557 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15558;
  wire [0:0] v_15559;
  wire [0:0] v_15560;
  wire [0:0] v_15561;
  function [0:0] mux_15561(input [0:0] sel);
    case (sel) 0: mux_15561 = 1'h0; 1: mux_15561 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15562;
  function [0:0] mux_15562(input [0:0] sel);
    case (sel) 0: mux_15562 = 1'h0; 1: mux_15562 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15563;
  wire [0:0] v_15564;
  wire [0:0] v_15565;
  wire [0:0] v_15566;
  wire [0:0] v_15567;
  wire [0:0] v_15568;
  function [0:0] mux_15568(input [0:0] sel);
    case (sel) 0: mux_15568 = 1'h0; 1: mux_15568 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15569;
  function [0:0] mux_15569(input [0:0] sel);
    case (sel) 0: mux_15569 = 1'h0; 1: mux_15569 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15570;
  wire [0:0] v_15571;
  wire [0:0] v_15572;
  wire [0:0] v_15573;
  function [0:0] mux_15573(input [0:0] sel);
    case (sel) 0: mux_15573 = 1'h0; 1: mux_15573 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15574;
  function [0:0] mux_15574(input [0:0] sel);
    case (sel) 0: mux_15574 = 1'h0; 1: mux_15574 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15575;
  wire [0:0] v_15576;
  wire [0:0] v_15577;
  wire [0:0] v_15578;
  wire [0:0] v_15579;
  wire [0:0] v_15580;
  function [0:0] mux_15580(input [0:0] sel);
    case (sel) 0: mux_15580 = 1'h0; 1: mux_15580 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15581;
  wire [0:0] v_15582;
  wire [0:0] v_15583;
  wire [0:0] v_15584;
  wire [0:0] v_15585;
  function [0:0] mux_15585(input [0:0] sel);
    case (sel) 0: mux_15585 = 1'h0; 1: mux_15585 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15586;
  wire [0:0] v_15587;
  wire [0:0] v_15588;
  wire [0:0] v_15589;
  function [0:0] mux_15589(input [0:0] sel);
    case (sel) 0: mux_15589 = 1'h0; 1: mux_15589 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15590;
  function [0:0] mux_15590(input [0:0] sel);
    case (sel) 0: mux_15590 = 1'h0; 1: mux_15590 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_15591 = 1'h0;
  wire [0:0] v_15592;
  wire [0:0] v_15593;
  wire [0:0] act_15594;
  wire [0:0] v_15595;
  wire [0:0] v_15596;
  wire [0:0] v_15597;
  reg [0:0] v_15598 = 1'h0;
  wire [0:0] v_15599;
  wire [0:0] v_15600;
  wire [0:0] act_15601;
  wire [0:0] v_15602;
  wire [0:0] v_15603;
  wire [0:0] v_15604;
  reg [0:0] v_15605 = 1'h0;
  wire [0:0] v_15606;
  wire [0:0] v_15607;
  wire [0:0] act_15608;
  wire [0:0] v_15609;
  wire [0:0] v_15610;
  wire [0:0] v_15611;
  reg [0:0] v_15612 = 1'h0;
  wire [0:0] v_15613;
  wire [0:0] v_15614;
  wire [0:0] act_15615;
  wire [0:0] v_15616;
  wire [0:0] v_15617;
  wire [0:0] v_15618;
  wire [0:0] vin0_consume_en_15619;
  wire [0:0] vout_canPeek_15619;
  wire [7:0] vout_peek_15619;
  wire [0:0] v_15620;
  wire [0:0] v_15621;
  function [0:0] mux_15621(input [0:0] sel);
    case (sel) 0: mux_15621 = 1'h0; 1: mux_15621 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15622;
  wire [0:0] v_15623;
  wire [0:0] v_15624;
  wire [0:0] v_15625;
  wire [0:0] v_15626;
  function [0:0] mux_15626(input [0:0] sel);
    case (sel) 0: mux_15626 = 1'h0; 1: mux_15626 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15627;
  wire [0:0] vin0_consume_en_15628;
  wire [0:0] vout_canPeek_15628;
  wire [7:0] vout_peek_15628;
  wire [0:0] v_15629;
  wire [0:0] v_15630;
  function [0:0] mux_15630(input [0:0] sel);
    case (sel) 0: mux_15630 = 1'h0; 1: mux_15630 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15631;
  function [0:0] mux_15631(input [0:0] sel);
    case (sel) 0: mux_15631 = 1'h0; 1: mux_15631 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15632;
  wire [0:0] v_15633;
  wire [0:0] v_15634;
  wire [0:0] v_15635;
  wire [0:0] v_15636;
  wire [0:0] v_15637;
  wire [0:0] v_15638;
  function [0:0] mux_15638(input [0:0] sel);
    case (sel) 0: mux_15638 = 1'h0; 1: mux_15638 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15639;
  wire [0:0] v_15640;
  wire [0:0] v_15641;
  wire [0:0] v_15642;
  wire [0:0] v_15643;
  function [0:0] mux_15643(input [0:0] sel);
    case (sel) 0: mux_15643 = 1'h0; 1: mux_15643 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15644;
  wire [0:0] v_15645;
  wire [0:0] v_15646;
  wire [0:0] v_15647;
  function [0:0] mux_15647(input [0:0] sel);
    case (sel) 0: mux_15647 = 1'h0; 1: mux_15647 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15648;
  function [0:0] mux_15648(input [0:0] sel);
    case (sel) 0: mux_15648 = 1'h0; 1: mux_15648 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_15649 = 1'h0;
  wire [0:0] v_15650;
  wire [0:0] v_15651;
  wire [0:0] act_15652;
  wire [0:0] v_15653;
  wire [0:0] v_15654;
  wire [0:0] v_15655;
  wire [0:0] vin0_consume_en_15656;
  wire [0:0] vout_canPeek_15656;
  wire [7:0] vout_peek_15656;
  wire [0:0] v_15657;
  wire [0:0] v_15658;
  function [0:0] mux_15658(input [0:0] sel);
    case (sel) 0: mux_15658 = 1'h0; 1: mux_15658 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15659;
  wire [0:0] v_15660;
  wire [0:0] v_15661;
  wire [0:0] v_15662;
  wire [0:0] v_15663;
  function [0:0] mux_15663(input [0:0] sel);
    case (sel) 0: mux_15663 = 1'h0; 1: mux_15663 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15664;
  wire [0:0] vin0_consume_en_15665;
  wire [0:0] vout_canPeek_15665;
  wire [7:0] vout_peek_15665;
  wire [0:0] v_15666;
  wire [0:0] v_15667;
  function [0:0] mux_15667(input [0:0] sel);
    case (sel) 0: mux_15667 = 1'h0; 1: mux_15667 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15668;
  function [0:0] mux_15668(input [0:0] sel);
    case (sel) 0: mux_15668 = 1'h0; 1: mux_15668 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15669;
  wire [0:0] v_15670;
  wire [0:0] v_15671;
  wire [0:0] v_15672;
  wire [0:0] v_15673;
  wire [0:0] v_15674;
  wire [0:0] v_15675;
  function [0:0] mux_15675(input [0:0] sel);
    case (sel) 0: mux_15675 = 1'h0; 1: mux_15675 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15676;
  function [0:0] mux_15676(input [0:0] sel);
    case (sel) 0: mux_15676 = 1'h0; 1: mux_15676 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15677;
  wire [0:0] v_15678;
  wire [0:0] v_15679;
  wire [0:0] v_15680;
  function [0:0] mux_15680(input [0:0] sel);
    case (sel) 0: mux_15680 = 1'h0; 1: mux_15680 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15681;
  function [0:0] mux_15681(input [0:0] sel);
    case (sel) 0: mux_15681 = 1'h0; 1: mux_15681 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15682;
  wire [0:0] v_15683;
  wire [0:0] v_15684;
  wire [0:0] v_15685;
  wire [0:0] v_15686;
  wire [0:0] v_15687;
  function [0:0] mux_15687(input [0:0] sel);
    case (sel) 0: mux_15687 = 1'h0; 1: mux_15687 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15688;
  wire [0:0] v_15689;
  wire [0:0] v_15690;
  wire [0:0] v_15691;
  wire [0:0] v_15692;
  function [0:0] mux_15692(input [0:0] sel);
    case (sel) 0: mux_15692 = 1'h0; 1: mux_15692 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15693;
  wire [0:0] v_15694;
  wire [0:0] v_15695;
  wire [0:0] v_15696;
  function [0:0] mux_15696(input [0:0] sel);
    case (sel) 0: mux_15696 = 1'h0; 1: mux_15696 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15697;
  function [0:0] mux_15697(input [0:0] sel);
    case (sel) 0: mux_15697 = 1'h0; 1: mux_15697 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_15698 = 1'h0;
  wire [0:0] v_15699;
  wire [0:0] v_15700;
  wire [0:0] act_15701;
  wire [0:0] v_15702;
  wire [0:0] v_15703;
  wire [0:0] v_15704;
  reg [0:0] v_15705 = 1'h0;
  wire [0:0] v_15706;
  wire [0:0] v_15707;
  wire [0:0] act_15708;
  wire [0:0] v_15709;
  wire [0:0] v_15710;
  wire [0:0] v_15711;
  wire [0:0] vin0_consume_en_15712;
  wire [0:0] vout_canPeek_15712;
  wire [7:0] vout_peek_15712;
  wire [0:0] v_15713;
  wire [0:0] v_15714;
  function [0:0] mux_15714(input [0:0] sel);
    case (sel) 0: mux_15714 = 1'h0; 1: mux_15714 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15715;
  wire [0:0] v_15716;
  wire [0:0] v_15717;
  wire [0:0] v_15718;
  wire [0:0] v_15719;
  function [0:0] mux_15719(input [0:0] sel);
    case (sel) 0: mux_15719 = 1'h0; 1: mux_15719 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15720;
  wire [0:0] vin0_consume_en_15721;
  wire [0:0] vout_canPeek_15721;
  wire [7:0] vout_peek_15721;
  wire [0:0] v_15722;
  wire [0:0] v_15723;
  function [0:0] mux_15723(input [0:0] sel);
    case (sel) 0: mux_15723 = 1'h0; 1: mux_15723 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15724;
  function [0:0] mux_15724(input [0:0] sel);
    case (sel) 0: mux_15724 = 1'h0; 1: mux_15724 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15725;
  wire [0:0] v_15726;
  wire [0:0] v_15727;
  wire [0:0] v_15728;
  wire [0:0] v_15729;
  wire [0:0] v_15730;
  wire [0:0] v_15731;
  function [0:0] mux_15731(input [0:0] sel);
    case (sel) 0: mux_15731 = 1'h0; 1: mux_15731 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15732;
  wire [0:0] v_15733;
  wire [0:0] v_15734;
  wire [0:0] v_15735;
  wire [0:0] v_15736;
  function [0:0] mux_15736(input [0:0] sel);
    case (sel) 0: mux_15736 = 1'h0; 1: mux_15736 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15737;
  wire [0:0] v_15738;
  wire [0:0] v_15739;
  wire [0:0] v_15740;
  function [0:0] mux_15740(input [0:0] sel);
    case (sel) 0: mux_15740 = 1'h0; 1: mux_15740 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15741;
  function [0:0] mux_15741(input [0:0] sel);
    case (sel) 0: mux_15741 = 1'h0; 1: mux_15741 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_15742 = 1'h0;
  wire [0:0] v_15743;
  wire [0:0] v_15744;
  wire [0:0] act_15745;
  wire [0:0] v_15746;
  wire [0:0] v_15747;
  wire [0:0] v_15748;
  wire [0:0] vin0_consume_en_15749;
  wire [0:0] vout_canPeek_15749;
  wire [7:0] vout_peek_15749;
  wire [0:0] v_15750;
  wire [0:0] v_15751;
  function [0:0] mux_15751(input [0:0] sel);
    case (sel) 0: mux_15751 = 1'h0; 1: mux_15751 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15752;
  wire [0:0] v_15753;
  wire [0:0] v_15754;
  wire [0:0] v_15755;
  wire [0:0] v_15756;
  function [0:0] mux_15756(input [0:0] sel);
    case (sel) 0: mux_15756 = 1'h0; 1: mux_15756 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15757;
  wire [0:0] vin0_consume_en_15758;
  wire [0:0] vout_canPeek_15758;
  wire [7:0] vout_peek_15758;
  wire [0:0] v_15759;
  wire [0:0] v_15760;
  function [0:0] mux_15760(input [0:0] sel);
    case (sel) 0: mux_15760 = 1'h0; 1: mux_15760 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15761;
  function [0:0] mux_15761(input [0:0] sel);
    case (sel) 0: mux_15761 = 1'h0; 1: mux_15761 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15762;
  wire [0:0] v_15763;
  wire [0:0] v_15764;
  wire [0:0] v_15765;
  wire [0:0] v_15766;
  wire [0:0] v_15767;
  wire [0:0] v_15768;
  function [0:0] mux_15768(input [0:0] sel);
    case (sel) 0: mux_15768 = 1'h0; 1: mux_15768 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15769;
  function [0:0] mux_15769(input [0:0] sel);
    case (sel) 0: mux_15769 = 1'h0; 1: mux_15769 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15770;
  wire [0:0] v_15771;
  wire [0:0] v_15772;
  wire [0:0] v_15773;
  function [0:0] mux_15773(input [0:0] sel);
    case (sel) 0: mux_15773 = 1'h0; 1: mux_15773 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15774;
  function [0:0] mux_15774(input [0:0] sel);
    case (sel) 0: mux_15774 = 1'h0; 1: mux_15774 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15775;
  wire [0:0] v_15776;
  wire [0:0] v_15777;
  wire [0:0] v_15778;
  wire [0:0] v_15779;
  wire [0:0] v_15780;
  function [0:0] mux_15780(input [0:0] sel);
    case (sel) 0: mux_15780 = 1'h0; 1: mux_15780 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15781;
  function [0:0] mux_15781(input [0:0] sel);
    case (sel) 0: mux_15781 = 1'h0; 1: mux_15781 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15782;
  wire [0:0] v_15783;
  wire [0:0] v_15784;
  wire [0:0] v_15785;
  function [0:0] mux_15785(input [0:0] sel);
    case (sel) 0: mux_15785 = 1'h0; 1: mux_15785 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15786;
  function [0:0] mux_15786(input [0:0] sel);
    case (sel) 0: mux_15786 = 1'h0; 1: mux_15786 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15787;
  wire [0:0] v_15788;
  wire [0:0] v_15789;
  wire [0:0] v_15790;
  wire [0:0] v_15791;
  wire [0:0] v_15792;
  function [0:0] mux_15792(input [0:0] sel);
    case (sel) 0: mux_15792 = 1'h0; 1: mux_15792 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15793;
  wire [0:0] v_15794;
  wire [0:0] v_15795;
  wire [0:0] v_15796;
  wire [0:0] v_15797;
  function [0:0] mux_15797(input [0:0] sel);
    case (sel) 0: mux_15797 = 1'h0; 1: mux_15797 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15798;
  wire [0:0] v_15799;
  wire [0:0] v_15800;
  wire [0:0] v_15801;
  function [0:0] mux_15801(input [0:0] sel);
    case (sel) 0: mux_15801 = 1'h0; 1: mux_15801 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15802;
  function [0:0] mux_15802(input [0:0] sel);
    case (sel) 0: mux_15802 = 1'h0; 1: mux_15802 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_15803 = 1'h0;
  wire [0:0] v_15804;
  wire [0:0] v_15805;
  wire [0:0] act_15806;
  wire [0:0] v_15807;
  wire [0:0] v_15808;
  wire [0:0] v_15809;
  reg [0:0] v_15810 = 1'h0;
  wire [0:0] v_15811;
  wire [0:0] v_15812;
  wire [0:0] act_15813;
  wire [0:0] v_15814;
  wire [0:0] v_15815;
  wire [0:0] v_15816;
  reg [0:0] v_15817 = 1'h0;
  wire [0:0] v_15818;
  wire [0:0] v_15819;
  wire [0:0] act_15820;
  wire [0:0] v_15821;
  wire [0:0] v_15822;
  wire [0:0] v_15823;
  wire [0:0] vin0_consume_en_15824;
  wire [0:0] vout_canPeek_15824;
  wire [7:0] vout_peek_15824;
  wire [0:0] v_15825;
  wire [0:0] v_15826;
  function [0:0] mux_15826(input [0:0] sel);
    case (sel) 0: mux_15826 = 1'h0; 1: mux_15826 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15827;
  wire [0:0] v_15828;
  wire [0:0] v_15829;
  wire [0:0] v_15830;
  wire [0:0] v_15831;
  function [0:0] mux_15831(input [0:0] sel);
    case (sel) 0: mux_15831 = 1'h0; 1: mux_15831 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15832;
  wire [0:0] vin0_consume_en_15833;
  wire [0:0] vout_canPeek_15833;
  wire [7:0] vout_peek_15833;
  wire [0:0] v_15834;
  wire [0:0] v_15835;
  function [0:0] mux_15835(input [0:0] sel);
    case (sel) 0: mux_15835 = 1'h0; 1: mux_15835 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15836;
  function [0:0] mux_15836(input [0:0] sel);
    case (sel) 0: mux_15836 = 1'h0; 1: mux_15836 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15837;
  wire [0:0] v_15838;
  wire [0:0] v_15839;
  wire [0:0] v_15840;
  wire [0:0] v_15841;
  wire [0:0] v_15842;
  wire [0:0] v_15843;
  function [0:0] mux_15843(input [0:0] sel);
    case (sel) 0: mux_15843 = 1'h0; 1: mux_15843 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15844;
  wire [0:0] v_15845;
  wire [0:0] v_15846;
  wire [0:0] v_15847;
  wire [0:0] v_15848;
  function [0:0] mux_15848(input [0:0] sel);
    case (sel) 0: mux_15848 = 1'h0; 1: mux_15848 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15849;
  wire [0:0] v_15850;
  wire [0:0] v_15851;
  wire [0:0] v_15852;
  function [0:0] mux_15852(input [0:0] sel);
    case (sel) 0: mux_15852 = 1'h0; 1: mux_15852 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15853;
  function [0:0] mux_15853(input [0:0] sel);
    case (sel) 0: mux_15853 = 1'h0; 1: mux_15853 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_15854 = 1'h0;
  wire [0:0] v_15855;
  wire [0:0] v_15856;
  wire [0:0] act_15857;
  wire [0:0] v_15858;
  wire [0:0] v_15859;
  wire [0:0] v_15860;
  wire [0:0] vin0_consume_en_15861;
  wire [0:0] vout_canPeek_15861;
  wire [7:0] vout_peek_15861;
  wire [0:0] v_15862;
  wire [0:0] v_15863;
  function [0:0] mux_15863(input [0:0] sel);
    case (sel) 0: mux_15863 = 1'h0; 1: mux_15863 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15864;
  wire [0:0] v_15865;
  wire [0:0] v_15866;
  wire [0:0] v_15867;
  wire [0:0] v_15868;
  function [0:0] mux_15868(input [0:0] sel);
    case (sel) 0: mux_15868 = 1'h0; 1: mux_15868 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15869;
  wire [0:0] vin0_consume_en_15870;
  wire [0:0] vout_canPeek_15870;
  wire [7:0] vout_peek_15870;
  wire [0:0] v_15871;
  wire [0:0] v_15872;
  function [0:0] mux_15872(input [0:0] sel);
    case (sel) 0: mux_15872 = 1'h0; 1: mux_15872 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15873;
  function [0:0] mux_15873(input [0:0] sel);
    case (sel) 0: mux_15873 = 1'h0; 1: mux_15873 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15874;
  wire [0:0] v_15875;
  wire [0:0] v_15876;
  wire [0:0] v_15877;
  wire [0:0] v_15878;
  wire [0:0] v_15879;
  wire [0:0] v_15880;
  function [0:0] mux_15880(input [0:0] sel);
    case (sel) 0: mux_15880 = 1'h0; 1: mux_15880 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15881;
  function [0:0] mux_15881(input [0:0] sel);
    case (sel) 0: mux_15881 = 1'h0; 1: mux_15881 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15882;
  wire [0:0] v_15883;
  wire [0:0] v_15884;
  wire [0:0] v_15885;
  function [0:0] mux_15885(input [0:0] sel);
    case (sel) 0: mux_15885 = 1'h0; 1: mux_15885 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15886;
  function [0:0] mux_15886(input [0:0] sel);
    case (sel) 0: mux_15886 = 1'h0; 1: mux_15886 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15887;
  wire [0:0] v_15888;
  wire [0:0] v_15889;
  wire [0:0] v_15890;
  wire [0:0] v_15891;
  wire [0:0] v_15892;
  function [0:0] mux_15892(input [0:0] sel);
    case (sel) 0: mux_15892 = 1'h0; 1: mux_15892 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15893;
  wire [0:0] v_15894;
  wire [0:0] v_15895;
  wire [0:0] v_15896;
  wire [0:0] v_15897;
  function [0:0] mux_15897(input [0:0] sel);
    case (sel) 0: mux_15897 = 1'h0; 1: mux_15897 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15898;
  wire [0:0] v_15899;
  wire [0:0] v_15900;
  wire [0:0] v_15901;
  function [0:0] mux_15901(input [0:0] sel);
    case (sel) 0: mux_15901 = 1'h0; 1: mux_15901 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15902;
  function [0:0] mux_15902(input [0:0] sel);
    case (sel) 0: mux_15902 = 1'h0; 1: mux_15902 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_15903 = 1'h0;
  wire [0:0] v_15904;
  wire [0:0] v_15905;
  wire [0:0] act_15906;
  wire [0:0] v_15907;
  wire [0:0] v_15908;
  wire [0:0] v_15909;
  reg [0:0] v_15910 = 1'h0;
  wire [0:0] v_15911;
  wire [0:0] v_15912;
  wire [0:0] act_15913;
  wire [0:0] v_15914;
  wire [0:0] v_15915;
  wire [0:0] v_15916;
  wire [0:0] vin0_consume_en_15917;
  wire [0:0] vout_canPeek_15917;
  wire [7:0] vout_peek_15917;
  wire [0:0] v_15918;
  wire [0:0] v_15919;
  function [0:0] mux_15919(input [0:0] sel);
    case (sel) 0: mux_15919 = 1'h0; 1: mux_15919 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15920;
  wire [0:0] v_15921;
  wire [0:0] v_15922;
  wire [0:0] v_15923;
  wire [0:0] v_15924;
  function [0:0] mux_15924(input [0:0] sel);
    case (sel) 0: mux_15924 = 1'h0; 1: mux_15924 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15925;
  wire [0:0] vin0_consume_en_15926;
  wire [0:0] vout_canPeek_15926;
  wire [7:0] vout_peek_15926;
  wire [0:0] v_15927;
  wire [0:0] v_15928;
  function [0:0] mux_15928(input [0:0] sel);
    case (sel) 0: mux_15928 = 1'h0; 1: mux_15928 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15929;
  function [0:0] mux_15929(input [0:0] sel);
    case (sel) 0: mux_15929 = 1'h0; 1: mux_15929 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15930;
  wire [0:0] v_15931;
  wire [0:0] v_15932;
  wire [0:0] v_15933;
  wire [0:0] v_15934;
  wire [0:0] v_15935;
  wire [0:0] v_15936;
  function [0:0] mux_15936(input [0:0] sel);
    case (sel) 0: mux_15936 = 1'h0; 1: mux_15936 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15937;
  wire [0:0] v_15938;
  wire [0:0] v_15939;
  wire [0:0] v_15940;
  wire [0:0] v_15941;
  function [0:0] mux_15941(input [0:0] sel);
    case (sel) 0: mux_15941 = 1'h0; 1: mux_15941 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15942;
  wire [0:0] v_15943;
  wire [0:0] v_15944;
  wire [0:0] v_15945;
  function [0:0] mux_15945(input [0:0] sel);
    case (sel) 0: mux_15945 = 1'h0; 1: mux_15945 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15946;
  function [0:0] mux_15946(input [0:0] sel);
    case (sel) 0: mux_15946 = 1'h0; 1: mux_15946 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_15947 = 1'h0;
  wire [0:0] v_15948;
  wire [0:0] v_15949;
  wire [0:0] act_15950;
  wire [0:0] v_15951;
  wire [0:0] v_15952;
  wire [0:0] v_15953;
  wire [0:0] vin0_consume_en_15954;
  wire [0:0] vout_canPeek_15954;
  wire [7:0] vout_peek_15954;
  wire [0:0] v_15955;
  wire [0:0] v_15956;
  function [0:0] mux_15956(input [0:0] sel);
    case (sel) 0: mux_15956 = 1'h0; 1: mux_15956 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15957;
  wire [0:0] v_15958;
  wire [0:0] v_15959;
  wire [0:0] v_15960;
  wire [0:0] v_15961;
  function [0:0] mux_15961(input [0:0] sel);
    case (sel) 0: mux_15961 = 1'h0; 1: mux_15961 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15962;
  wire [0:0] vin0_consume_en_15963;
  wire [0:0] vout_canPeek_15963;
  wire [7:0] vout_peek_15963;
  wire [0:0] v_15964;
  wire [0:0] v_15965;
  function [0:0] mux_15965(input [0:0] sel);
    case (sel) 0: mux_15965 = 1'h0; 1: mux_15965 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15966;
  function [0:0] mux_15966(input [0:0] sel);
    case (sel) 0: mux_15966 = 1'h0; 1: mux_15966 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15967;
  wire [0:0] v_15968;
  wire [0:0] v_15969;
  wire [0:0] v_15970;
  wire [0:0] v_15971;
  wire [0:0] v_15972;
  wire [0:0] v_15973;
  function [0:0] mux_15973(input [0:0] sel);
    case (sel) 0: mux_15973 = 1'h0; 1: mux_15973 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15974;
  function [0:0] mux_15974(input [0:0] sel);
    case (sel) 0: mux_15974 = 1'h0; 1: mux_15974 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15975;
  wire [0:0] v_15976;
  wire [0:0] v_15977;
  wire [0:0] v_15978;
  function [0:0] mux_15978(input [0:0] sel);
    case (sel) 0: mux_15978 = 1'h0; 1: mux_15978 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15979;
  function [0:0] mux_15979(input [0:0] sel);
    case (sel) 0: mux_15979 = 1'h0; 1: mux_15979 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15980;
  wire [0:0] v_15981;
  wire [0:0] v_15982;
  wire [0:0] v_15983;
  wire [0:0] v_15984;
  wire [0:0] v_15985;
  function [0:0] mux_15985(input [0:0] sel);
    case (sel) 0: mux_15985 = 1'h0; 1: mux_15985 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15986;
  function [0:0] mux_15986(input [0:0] sel);
    case (sel) 0: mux_15986 = 1'h0; 1: mux_15986 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15987;
  wire [0:0] v_15988;
  wire [0:0] v_15989;
  wire [0:0] v_15990;
  function [0:0] mux_15990(input [0:0] sel);
    case (sel) 0: mux_15990 = 1'h0; 1: mux_15990 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15991;
  function [0:0] mux_15991(input [0:0] sel);
    case (sel) 0: mux_15991 = 1'h0; 1: mux_15991 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15992;
  wire [0:0] v_15993;
  wire [0:0] v_15994;
  wire [0:0] v_15995;
  wire [0:0] v_15996;
  wire [0:0] v_15997;
  function [0:0] mux_15997(input [0:0] sel);
    case (sel) 0: mux_15997 = 1'h0; 1: mux_15997 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_15998;
  function [0:0] mux_15998(input [0:0] sel);
    case (sel) 0: mux_15998 = 1'h0; 1: mux_15998 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_15999;
  wire [0:0] v_16000;
  wire [0:0] v_16001;
  wire [0:0] v_16002;
  function [0:0] mux_16002(input [0:0] sel);
    case (sel) 0: mux_16002 = 1'h0; 1: mux_16002 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16003;
  function [0:0] mux_16003(input [0:0] sel);
    case (sel) 0: mux_16003 = 1'h0; 1: mux_16003 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16004;
  wire [0:0] v_16005;
  wire [0:0] v_16006;
  wire [0:0] v_16007;
  wire [0:0] v_16008;
  wire [0:0] v_16009;
  function [0:0] mux_16009(input [0:0] sel);
    case (sel) 0: mux_16009 = 1'h0; 1: mux_16009 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16010;
  function [0:0] mux_16010(input [0:0] sel);
    case (sel) 0: mux_16010 = 1'h0; 1: mux_16010 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16011;
  wire [0:0] v_16012;
  wire [0:0] v_16013;
  wire [0:0] v_16014;
  function [0:0] mux_16014(input [0:0] sel);
    case (sel) 0: mux_16014 = 1'h0; 1: mux_16014 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16015;
  function [0:0] mux_16015(input [0:0] sel);
    case (sel) 0: mux_16015 = 1'h0; 1: mux_16015 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16016;
  wire [0:0] v_16017;
  wire [0:0] v_16018;
  wire [0:0] v_16019;
  wire [0:0] v_16020;
  wire [0:0] v_16021;
  function [0:0] mux_16021(input [0:0] sel);
    case (sel) 0: mux_16021 = 1'h0; 1: mux_16021 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16022;
  wire [0:0] v_16023;
  wire [0:0] v_16024;
  wire [0:0] v_16025;
  wire [0:0] v_16026;
  function [0:0] mux_16026(input [0:0] sel);
    case (sel) 0: mux_16026 = 1'h0; 1: mux_16026 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16027;
  wire [0:0] v_16028;
  wire [0:0] v_16029;
  wire [0:0] v_16030;
  function [0:0] mux_16030(input [0:0] sel);
    case (sel) 0: mux_16030 = 1'h0; 1: mux_16030 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16031;
  function [0:0] mux_16031(input [0:0] sel);
    case (sel) 0: mux_16031 = 1'h0; 1: mux_16031 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_16032 = 1'h0;
  wire [0:0] v_16033;
  wire [0:0] v_16034;
  wire [0:0] act_16035;
  wire [0:0] v_16036;
  wire [0:0] v_16037;
  wire [0:0] v_16038;
  reg [0:0] v_16039 = 1'h0;
  wire [0:0] v_16040;
  wire [0:0] v_16041;
  wire [0:0] act_16042;
  wire [0:0] v_16043;
  wire [0:0] v_16044;
  wire [0:0] v_16045;
  reg [0:0] v_16046 = 1'h0;
  wire [0:0] v_16047;
  wire [0:0] v_16048;
  wire [0:0] act_16049;
  wire [0:0] v_16050;
  wire [0:0] v_16051;
  wire [0:0] v_16052;
  reg [0:0] v_16053 = 1'h0;
  wire [0:0] v_16054;
  wire [0:0] v_16055;
  wire [0:0] act_16056;
  wire [0:0] v_16057;
  wire [0:0] v_16058;
  wire [0:0] v_16059;
  reg [0:0] v_16060 = 1'h0;
  wire [0:0] v_16061;
  wire [0:0] v_16062;
  wire [0:0] act_16063;
  wire [0:0] v_16064;
  wire [0:0] v_16065;
  wire [0:0] v_16066;
  wire [0:0] vin0_consume_en_16067;
  wire [0:0] vout_canPeek_16067;
  wire [7:0] vout_peek_16067;
  wire [0:0] v_16068;
  wire [0:0] v_16069;
  function [0:0] mux_16069(input [0:0] sel);
    case (sel) 0: mux_16069 = 1'h0; 1: mux_16069 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16070;
  wire [0:0] v_16071;
  wire [0:0] v_16072;
  wire [0:0] v_16073;
  wire [0:0] v_16074;
  function [0:0] mux_16074(input [0:0] sel);
    case (sel) 0: mux_16074 = 1'h0; 1: mux_16074 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16075;
  wire [0:0] vin0_consume_en_16076;
  wire [0:0] vout_canPeek_16076;
  wire [7:0] vout_peek_16076;
  wire [0:0] v_16077;
  wire [0:0] v_16078;
  function [0:0] mux_16078(input [0:0] sel);
    case (sel) 0: mux_16078 = 1'h0; 1: mux_16078 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16079;
  function [0:0] mux_16079(input [0:0] sel);
    case (sel) 0: mux_16079 = 1'h0; 1: mux_16079 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16080;
  wire [0:0] v_16081;
  wire [0:0] v_16082;
  wire [0:0] v_16083;
  wire [0:0] v_16084;
  wire [0:0] v_16085;
  wire [0:0] v_16086;
  function [0:0] mux_16086(input [0:0] sel);
    case (sel) 0: mux_16086 = 1'h0; 1: mux_16086 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16087;
  wire [0:0] v_16088;
  wire [0:0] v_16089;
  wire [0:0] v_16090;
  wire [0:0] v_16091;
  function [0:0] mux_16091(input [0:0] sel);
    case (sel) 0: mux_16091 = 1'h0; 1: mux_16091 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16092;
  wire [0:0] v_16093;
  wire [0:0] v_16094;
  wire [0:0] v_16095;
  function [0:0] mux_16095(input [0:0] sel);
    case (sel) 0: mux_16095 = 1'h0; 1: mux_16095 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16096;
  function [0:0] mux_16096(input [0:0] sel);
    case (sel) 0: mux_16096 = 1'h0; 1: mux_16096 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_16097 = 1'h0;
  wire [0:0] v_16098;
  wire [0:0] v_16099;
  wire [0:0] act_16100;
  wire [0:0] v_16101;
  wire [0:0] v_16102;
  wire [0:0] v_16103;
  wire [0:0] vin0_consume_en_16104;
  wire [0:0] vout_canPeek_16104;
  wire [7:0] vout_peek_16104;
  wire [0:0] v_16105;
  wire [0:0] v_16106;
  function [0:0] mux_16106(input [0:0] sel);
    case (sel) 0: mux_16106 = 1'h0; 1: mux_16106 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16107;
  wire [0:0] v_16108;
  wire [0:0] v_16109;
  wire [0:0] v_16110;
  wire [0:0] v_16111;
  function [0:0] mux_16111(input [0:0] sel);
    case (sel) 0: mux_16111 = 1'h0; 1: mux_16111 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16112;
  wire [0:0] vin0_consume_en_16113;
  wire [0:0] vout_canPeek_16113;
  wire [7:0] vout_peek_16113;
  wire [0:0] v_16114;
  wire [0:0] v_16115;
  function [0:0] mux_16115(input [0:0] sel);
    case (sel) 0: mux_16115 = 1'h0; 1: mux_16115 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16116;
  function [0:0] mux_16116(input [0:0] sel);
    case (sel) 0: mux_16116 = 1'h0; 1: mux_16116 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16117;
  wire [0:0] v_16118;
  wire [0:0] v_16119;
  wire [0:0] v_16120;
  wire [0:0] v_16121;
  wire [0:0] v_16122;
  wire [0:0] v_16123;
  function [0:0] mux_16123(input [0:0] sel);
    case (sel) 0: mux_16123 = 1'h0; 1: mux_16123 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16124;
  function [0:0] mux_16124(input [0:0] sel);
    case (sel) 0: mux_16124 = 1'h0; 1: mux_16124 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16125;
  wire [0:0] v_16126;
  wire [0:0] v_16127;
  wire [0:0] v_16128;
  function [0:0] mux_16128(input [0:0] sel);
    case (sel) 0: mux_16128 = 1'h0; 1: mux_16128 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16129;
  function [0:0] mux_16129(input [0:0] sel);
    case (sel) 0: mux_16129 = 1'h0; 1: mux_16129 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16130;
  wire [0:0] v_16131;
  wire [0:0] v_16132;
  wire [0:0] v_16133;
  wire [0:0] v_16134;
  wire [0:0] v_16135;
  function [0:0] mux_16135(input [0:0] sel);
    case (sel) 0: mux_16135 = 1'h0; 1: mux_16135 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16136;
  wire [0:0] v_16137;
  wire [0:0] v_16138;
  wire [0:0] v_16139;
  wire [0:0] v_16140;
  function [0:0] mux_16140(input [0:0] sel);
    case (sel) 0: mux_16140 = 1'h0; 1: mux_16140 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16141;
  wire [0:0] v_16142;
  wire [0:0] v_16143;
  wire [0:0] v_16144;
  function [0:0] mux_16144(input [0:0] sel);
    case (sel) 0: mux_16144 = 1'h0; 1: mux_16144 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16145;
  function [0:0] mux_16145(input [0:0] sel);
    case (sel) 0: mux_16145 = 1'h0; 1: mux_16145 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_16146 = 1'h0;
  wire [0:0] v_16147;
  wire [0:0] v_16148;
  wire [0:0] act_16149;
  wire [0:0] v_16150;
  wire [0:0] v_16151;
  wire [0:0] v_16152;
  reg [0:0] v_16153 = 1'h0;
  wire [0:0] v_16154;
  wire [0:0] v_16155;
  wire [0:0] act_16156;
  wire [0:0] v_16157;
  wire [0:0] v_16158;
  wire [0:0] v_16159;
  wire [0:0] vin0_consume_en_16160;
  wire [0:0] vout_canPeek_16160;
  wire [7:0] vout_peek_16160;
  wire [0:0] v_16161;
  wire [0:0] v_16162;
  function [0:0] mux_16162(input [0:0] sel);
    case (sel) 0: mux_16162 = 1'h0; 1: mux_16162 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16163;
  wire [0:0] v_16164;
  wire [0:0] v_16165;
  wire [0:0] v_16166;
  wire [0:0] v_16167;
  function [0:0] mux_16167(input [0:0] sel);
    case (sel) 0: mux_16167 = 1'h0; 1: mux_16167 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16168;
  wire [0:0] vin0_consume_en_16169;
  wire [0:0] vout_canPeek_16169;
  wire [7:0] vout_peek_16169;
  wire [0:0] v_16170;
  wire [0:0] v_16171;
  function [0:0] mux_16171(input [0:0] sel);
    case (sel) 0: mux_16171 = 1'h0; 1: mux_16171 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16172;
  function [0:0] mux_16172(input [0:0] sel);
    case (sel) 0: mux_16172 = 1'h0; 1: mux_16172 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16173;
  wire [0:0] v_16174;
  wire [0:0] v_16175;
  wire [0:0] v_16176;
  wire [0:0] v_16177;
  wire [0:0] v_16178;
  wire [0:0] v_16179;
  function [0:0] mux_16179(input [0:0] sel);
    case (sel) 0: mux_16179 = 1'h0; 1: mux_16179 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16180;
  wire [0:0] v_16181;
  wire [0:0] v_16182;
  wire [0:0] v_16183;
  wire [0:0] v_16184;
  function [0:0] mux_16184(input [0:0] sel);
    case (sel) 0: mux_16184 = 1'h0; 1: mux_16184 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16185;
  wire [0:0] v_16186;
  wire [0:0] v_16187;
  wire [0:0] v_16188;
  function [0:0] mux_16188(input [0:0] sel);
    case (sel) 0: mux_16188 = 1'h0; 1: mux_16188 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16189;
  function [0:0] mux_16189(input [0:0] sel);
    case (sel) 0: mux_16189 = 1'h0; 1: mux_16189 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_16190 = 1'h0;
  wire [0:0] v_16191;
  wire [0:0] v_16192;
  wire [0:0] act_16193;
  wire [0:0] v_16194;
  wire [0:0] v_16195;
  wire [0:0] v_16196;
  wire [0:0] vin0_consume_en_16197;
  wire [0:0] vout_canPeek_16197;
  wire [7:0] vout_peek_16197;
  wire [0:0] v_16198;
  wire [0:0] v_16199;
  function [0:0] mux_16199(input [0:0] sel);
    case (sel) 0: mux_16199 = 1'h0; 1: mux_16199 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16200;
  wire [0:0] v_16201;
  wire [0:0] v_16202;
  wire [0:0] v_16203;
  wire [0:0] v_16204;
  function [0:0] mux_16204(input [0:0] sel);
    case (sel) 0: mux_16204 = 1'h0; 1: mux_16204 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16205;
  wire [0:0] vin0_consume_en_16206;
  wire [0:0] vout_canPeek_16206;
  wire [7:0] vout_peek_16206;
  wire [0:0] v_16207;
  wire [0:0] v_16208;
  function [0:0] mux_16208(input [0:0] sel);
    case (sel) 0: mux_16208 = 1'h0; 1: mux_16208 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16209;
  function [0:0] mux_16209(input [0:0] sel);
    case (sel) 0: mux_16209 = 1'h0; 1: mux_16209 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16210;
  wire [0:0] v_16211;
  wire [0:0] v_16212;
  wire [0:0] v_16213;
  wire [0:0] v_16214;
  wire [0:0] v_16215;
  wire [0:0] v_16216;
  function [0:0] mux_16216(input [0:0] sel);
    case (sel) 0: mux_16216 = 1'h0; 1: mux_16216 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16217;
  function [0:0] mux_16217(input [0:0] sel);
    case (sel) 0: mux_16217 = 1'h0; 1: mux_16217 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16218;
  wire [0:0] v_16219;
  wire [0:0] v_16220;
  wire [0:0] v_16221;
  function [0:0] mux_16221(input [0:0] sel);
    case (sel) 0: mux_16221 = 1'h0; 1: mux_16221 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16222;
  function [0:0] mux_16222(input [0:0] sel);
    case (sel) 0: mux_16222 = 1'h0; 1: mux_16222 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16223;
  wire [0:0] v_16224;
  wire [0:0] v_16225;
  wire [0:0] v_16226;
  wire [0:0] v_16227;
  wire [0:0] v_16228;
  function [0:0] mux_16228(input [0:0] sel);
    case (sel) 0: mux_16228 = 1'h0; 1: mux_16228 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16229;
  function [0:0] mux_16229(input [0:0] sel);
    case (sel) 0: mux_16229 = 1'h0; 1: mux_16229 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16230;
  wire [0:0] v_16231;
  wire [0:0] v_16232;
  wire [0:0] v_16233;
  function [0:0] mux_16233(input [0:0] sel);
    case (sel) 0: mux_16233 = 1'h0; 1: mux_16233 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16234;
  function [0:0] mux_16234(input [0:0] sel);
    case (sel) 0: mux_16234 = 1'h0; 1: mux_16234 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16235;
  wire [0:0] v_16236;
  wire [0:0] v_16237;
  wire [0:0] v_16238;
  wire [0:0] v_16239;
  wire [0:0] v_16240;
  function [0:0] mux_16240(input [0:0] sel);
    case (sel) 0: mux_16240 = 1'h0; 1: mux_16240 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16241;
  wire [0:0] v_16242;
  wire [0:0] v_16243;
  wire [0:0] v_16244;
  wire [0:0] v_16245;
  function [0:0] mux_16245(input [0:0] sel);
    case (sel) 0: mux_16245 = 1'h0; 1: mux_16245 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16246;
  wire [0:0] v_16247;
  wire [0:0] v_16248;
  wire [0:0] v_16249;
  function [0:0] mux_16249(input [0:0] sel);
    case (sel) 0: mux_16249 = 1'h0; 1: mux_16249 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16250;
  function [0:0] mux_16250(input [0:0] sel);
    case (sel) 0: mux_16250 = 1'h0; 1: mux_16250 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_16251 = 1'h0;
  wire [0:0] v_16252;
  wire [0:0] v_16253;
  wire [0:0] act_16254;
  wire [0:0] v_16255;
  wire [0:0] v_16256;
  wire [0:0] v_16257;
  reg [0:0] v_16258 = 1'h0;
  wire [0:0] v_16259;
  wire [0:0] v_16260;
  wire [0:0] act_16261;
  wire [0:0] v_16262;
  wire [0:0] v_16263;
  wire [0:0] v_16264;
  reg [0:0] v_16265 = 1'h0;
  wire [0:0] v_16266;
  wire [0:0] v_16267;
  wire [0:0] act_16268;
  wire [0:0] v_16269;
  wire [0:0] v_16270;
  wire [0:0] v_16271;
  wire [0:0] vin0_consume_en_16272;
  wire [0:0] vout_canPeek_16272;
  wire [7:0] vout_peek_16272;
  wire [0:0] v_16273;
  wire [0:0] v_16274;
  function [0:0] mux_16274(input [0:0] sel);
    case (sel) 0: mux_16274 = 1'h0; 1: mux_16274 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16275;
  wire [0:0] v_16276;
  wire [0:0] v_16277;
  wire [0:0] v_16278;
  wire [0:0] v_16279;
  function [0:0] mux_16279(input [0:0] sel);
    case (sel) 0: mux_16279 = 1'h0; 1: mux_16279 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16280;
  wire [0:0] vin0_consume_en_16281;
  wire [0:0] vout_canPeek_16281;
  wire [7:0] vout_peek_16281;
  wire [0:0] v_16282;
  wire [0:0] v_16283;
  function [0:0] mux_16283(input [0:0] sel);
    case (sel) 0: mux_16283 = 1'h0; 1: mux_16283 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16284;
  function [0:0] mux_16284(input [0:0] sel);
    case (sel) 0: mux_16284 = 1'h0; 1: mux_16284 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16285;
  wire [0:0] v_16286;
  wire [0:0] v_16287;
  wire [0:0] v_16288;
  wire [0:0] v_16289;
  wire [0:0] v_16290;
  wire [0:0] v_16291;
  function [0:0] mux_16291(input [0:0] sel);
    case (sel) 0: mux_16291 = 1'h0; 1: mux_16291 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16292;
  wire [0:0] v_16293;
  wire [0:0] v_16294;
  wire [0:0] v_16295;
  wire [0:0] v_16296;
  function [0:0] mux_16296(input [0:0] sel);
    case (sel) 0: mux_16296 = 1'h0; 1: mux_16296 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16297;
  wire [0:0] v_16298;
  wire [0:0] v_16299;
  wire [0:0] v_16300;
  function [0:0] mux_16300(input [0:0] sel);
    case (sel) 0: mux_16300 = 1'h0; 1: mux_16300 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16301;
  function [0:0] mux_16301(input [0:0] sel);
    case (sel) 0: mux_16301 = 1'h0; 1: mux_16301 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_16302 = 1'h0;
  wire [0:0] v_16303;
  wire [0:0] v_16304;
  wire [0:0] act_16305;
  wire [0:0] v_16306;
  wire [0:0] v_16307;
  wire [0:0] v_16308;
  wire [0:0] vin0_consume_en_16309;
  wire [0:0] vout_canPeek_16309;
  wire [7:0] vout_peek_16309;
  wire [0:0] v_16310;
  wire [0:0] v_16311;
  function [0:0] mux_16311(input [0:0] sel);
    case (sel) 0: mux_16311 = 1'h0; 1: mux_16311 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16312;
  wire [0:0] v_16313;
  wire [0:0] v_16314;
  wire [0:0] v_16315;
  wire [0:0] v_16316;
  function [0:0] mux_16316(input [0:0] sel);
    case (sel) 0: mux_16316 = 1'h0; 1: mux_16316 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16317;
  wire [0:0] vin0_consume_en_16318;
  wire [0:0] vout_canPeek_16318;
  wire [7:0] vout_peek_16318;
  wire [0:0] v_16319;
  wire [0:0] v_16320;
  function [0:0] mux_16320(input [0:0] sel);
    case (sel) 0: mux_16320 = 1'h0; 1: mux_16320 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16321;
  function [0:0] mux_16321(input [0:0] sel);
    case (sel) 0: mux_16321 = 1'h0; 1: mux_16321 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16322;
  wire [0:0] v_16323;
  wire [0:0] v_16324;
  wire [0:0] v_16325;
  wire [0:0] v_16326;
  wire [0:0] v_16327;
  wire [0:0] v_16328;
  function [0:0] mux_16328(input [0:0] sel);
    case (sel) 0: mux_16328 = 1'h0; 1: mux_16328 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16329;
  function [0:0] mux_16329(input [0:0] sel);
    case (sel) 0: mux_16329 = 1'h0; 1: mux_16329 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16330;
  wire [0:0] v_16331;
  wire [0:0] v_16332;
  wire [0:0] v_16333;
  function [0:0] mux_16333(input [0:0] sel);
    case (sel) 0: mux_16333 = 1'h0; 1: mux_16333 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16334;
  function [0:0] mux_16334(input [0:0] sel);
    case (sel) 0: mux_16334 = 1'h0; 1: mux_16334 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16335;
  wire [0:0] v_16336;
  wire [0:0] v_16337;
  wire [0:0] v_16338;
  wire [0:0] v_16339;
  wire [0:0] v_16340;
  function [0:0] mux_16340(input [0:0] sel);
    case (sel) 0: mux_16340 = 1'h0; 1: mux_16340 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16341;
  wire [0:0] v_16342;
  wire [0:0] v_16343;
  wire [0:0] v_16344;
  wire [0:0] v_16345;
  function [0:0] mux_16345(input [0:0] sel);
    case (sel) 0: mux_16345 = 1'h0; 1: mux_16345 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16346;
  wire [0:0] v_16347;
  wire [0:0] v_16348;
  wire [0:0] v_16349;
  function [0:0] mux_16349(input [0:0] sel);
    case (sel) 0: mux_16349 = 1'h0; 1: mux_16349 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16350;
  function [0:0] mux_16350(input [0:0] sel);
    case (sel) 0: mux_16350 = 1'h0; 1: mux_16350 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_16351 = 1'h0;
  wire [0:0] v_16352;
  wire [0:0] v_16353;
  wire [0:0] act_16354;
  wire [0:0] v_16355;
  wire [0:0] v_16356;
  wire [0:0] v_16357;
  reg [0:0] v_16358 = 1'h0;
  wire [0:0] v_16359;
  wire [0:0] v_16360;
  wire [0:0] act_16361;
  wire [0:0] v_16362;
  wire [0:0] v_16363;
  wire [0:0] v_16364;
  wire [0:0] vin0_consume_en_16365;
  wire [0:0] vout_canPeek_16365;
  wire [7:0] vout_peek_16365;
  wire [0:0] v_16366;
  wire [0:0] v_16367;
  function [0:0] mux_16367(input [0:0] sel);
    case (sel) 0: mux_16367 = 1'h0; 1: mux_16367 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16368;
  wire [0:0] v_16369;
  wire [0:0] v_16370;
  wire [0:0] v_16371;
  wire [0:0] v_16372;
  function [0:0] mux_16372(input [0:0] sel);
    case (sel) 0: mux_16372 = 1'h0; 1: mux_16372 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16373;
  wire [0:0] vin0_consume_en_16374;
  wire [0:0] vout_canPeek_16374;
  wire [7:0] vout_peek_16374;
  wire [0:0] v_16375;
  wire [0:0] v_16376;
  function [0:0] mux_16376(input [0:0] sel);
    case (sel) 0: mux_16376 = 1'h0; 1: mux_16376 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16377;
  function [0:0] mux_16377(input [0:0] sel);
    case (sel) 0: mux_16377 = 1'h0; 1: mux_16377 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16378;
  wire [0:0] v_16379;
  wire [0:0] v_16380;
  wire [0:0] v_16381;
  wire [0:0] v_16382;
  wire [0:0] v_16383;
  wire [0:0] v_16384;
  function [0:0] mux_16384(input [0:0] sel);
    case (sel) 0: mux_16384 = 1'h0; 1: mux_16384 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16385;
  wire [0:0] v_16386;
  wire [0:0] v_16387;
  wire [0:0] v_16388;
  wire [0:0] v_16389;
  function [0:0] mux_16389(input [0:0] sel);
    case (sel) 0: mux_16389 = 1'h0; 1: mux_16389 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16390;
  wire [0:0] v_16391;
  wire [0:0] v_16392;
  wire [0:0] v_16393;
  function [0:0] mux_16393(input [0:0] sel);
    case (sel) 0: mux_16393 = 1'h0; 1: mux_16393 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16394;
  function [0:0] mux_16394(input [0:0] sel);
    case (sel) 0: mux_16394 = 1'h0; 1: mux_16394 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_16395 = 1'h0;
  wire [0:0] v_16396;
  wire [0:0] v_16397;
  wire [0:0] act_16398;
  wire [0:0] v_16399;
  wire [0:0] v_16400;
  wire [0:0] v_16401;
  wire [0:0] vin0_consume_en_16402;
  wire [0:0] vout_canPeek_16402;
  wire [7:0] vout_peek_16402;
  wire [0:0] v_16403;
  wire [0:0] v_16404;
  function [0:0] mux_16404(input [0:0] sel);
    case (sel) 0: mux_16404 = 1'h0; 1: mux_16404 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16405;
  wire [0:0] v_16406;
  wire [0:0] v_16407;
  wire [0:0] v_16408;
  wire [0:0] v_16409;
  function [0:0] mux_16409(input [0:0] sel);
    case (sel) 0: mux_16409 = 1'h0; 1: mux_16409 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16410;
  wire [0:0] vin0_consume_en_16411;
  wire [0:0] vout_canPeek_16411;
  wire [7:0] vout_peek_16411;
  wire [0:0] v_16412;
  wire [0:0] v_16413;
  function [0:0] mux_16413(input [0:0] sel);
    case (sel) 0: mux_16413 = 1'h0; 1: mux_16413 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16414;
  function [0:0] mux_16414(input [0:0] sel);
    case (sel) 0: mux_16414 = 1'h0; 1: mux_16414 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16415;
  wire [0:0] v_16416;
  wire [0:0] v_16417;
  wire [0:0] v_16418;
  wire [0:0] v_16419;
  wire [0:0] v_16420;
  wire [0:0] v_16421;
  function [0:0] mux_16421(input [0:0] sel);
    case (sel) 0: mux_16421 = 1'h0; 1: mux_16421 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16422;
  function [0:0] mux_16422(input [0:0] sel);
    case (sel) 0: mux_16422 = 1'h0; 1: mux_16422 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16423;
  wire [0:0] v_16424;
  wire [0:0] v_16425;
  wire [0:0] v_16426;
  function [0:0] mux_16426(input [0:0] sel);
    case (sel) 0: mux_16426 = 1'h0; 1: mux_16426 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16427;
  function [0:0] mux_16427(input [0:0] sel);
    case (sel) 0: mux_16427 = 1'h0; 1: mux_16427 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16428;
  wire [0:0] v_16429;
  wire [0:0] v_16430;
  wire [0:0] v_16431;
  wire [0:0] v_16432;
  wire [0:0] v_16433;
  function [0:0] mux_16433(input [0:0] sel);
    case (sel) 0: mux_16433 = 1'h0; 1: mux_16433 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16434;
  function [0:0] mux_16434(input [0:0] sel);
    case (sel) 0: mux_16434 = 1'h0; 1: mux_16434 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16435;
  wire [0:0] v_16436;
  wire [0:0] v_16437;
  wire [0:0] v_16438;
  function [0:0] mux_16438(input [0:0] sel);
    case (sel) 0: mux_16438 = 1'h0; 1: mux_16438 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16439;
  function [0:0] mux_16439(input [0:0] sel);
    case (sel) 0: mux_16439 = 1'h0; 1: mux_16439 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16440;
  wire [0:0] v_16441;
  wire [0:0] v_16442;
  wire [0:0] v_16443;
  wire [0:0] v_16444;
  wire [0:0] v_16445;
  function [0:0] mux_16445(input [0:0] sel);
    case (sel) 0: mux_16445 = 1'h0; 1: mux_16445 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16446;
  function [0:0] mux_16446(input [0:0] sel);
    case (sel) 0: mux_16446 = 1'h0; 1: mux_16446 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16447;
  wire [0:0] v_16448;
  wire [0:0] v_16449;
  wire [0:0] v_16450;
  function [0:0] mux_16450(input [0:0] sel);
    case (sel) 0: mux_16450 = 1'h0; 1: mux_16450 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16451;
  function [0:0] mux_16451(input [0:0] sel);
    case (sel) 0: mux_16451 = 1'h0; 1: mux_16451 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16452;
  wire [0:0] v_16453;
  wire [0:0] v_16454;
  wire [0:0] v_16455;
  wire [0:0] v_16456;
  wire [0:0] v_16457;
  function [0:0] mux_16457(input [0:0] sel);
    case (sel) 0: mux_16457 = 1'h0; 1: mux_16457 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16458;
  wire [0:0] v_16459;
  wire [0:0] v_16460;
  wire [0:0] v_16461;
  wire [0:0] v_16462;
  function [0:0] mux_16462(input [0:0] sel);
    case (sel) 0: mux_16462 = 1'h0; 1: mux_16462 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16463;
  wire [0:0] v_16464;
  wire [0:0] v_16465;
  wire [0:0] v_16466;
  function [0:0] mux_16466(input [0:0] sel);
    case (sel) 0: mux_16466 = 1'h0; 1: mux_16466 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16467;
  function [0:0] mux_16467(input [0:0] sel);
    case (sel) 0: mux_16467 = 1'h0; 1: mux_16467 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_16468 = 1'h0;
  wire [0:0] v_16469;
  wire [0:0] v_16470;
  wire [0:0] act_16471;
  wire [0:0] v_16472;
  wire [0:0] v_16473;
  wire [0:0] v_16474;
  reg [0:0] v_16475 = 1'h0;
  wire [0:0] v_16476;
  wire [0:0] v_16477;
  wire [0:0] act_16478;
  wire [0:0] v_16479;
  wire [0:0] v_16480;
  wire [0:0] v_16481;
  reg [0:0] v_16482 = 1'h0;
  wire [0:0] v_16483;
  wire [0:0] v_16484;
  wire [0:0] act_16485;
  wire [0:0] v_16486;
  wire [0:0] v_16487;
  wire [0:0] v_16488;
  reg [0:0] v_16489 = 1'h0;
  wire [0:0] v_16490;
  wire [0:0] v_16491;
  wire [0:0] act_16492;
  wire [0:0] v_16493;
  wire [0:0] v_16494;
  wire [0:0] v_16495;
  wire [0:0] vin0_consume_en_16496;
  wire [0:0] vout_canPeek_16496;
  wire [7:0] vout_peek_16496;
  wire [0:0] v_16497;
  wire [0:0] v_16498;
  function [0:0] mux_16498(input [0:0] sel);
    case (sel) 0: mux_16498 = 1'h0; 1: mux_16498 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16499;
  wire [0:0] v_16500;
  wire [0:0] v_16501;
  wire [0:0] v_16502;
  wire [0:0] v_16503;
  function [0:0] mux_16503(input [0:0] sel);
    case (sel) 0: mux_16503 = 1'h0; 1: mux_16503 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16504;
  wire [0:0] vin0_consume_en_16505;
  wire [0:0] vout_canPeek_16505;
  wire [7:0] vout_peek_16505;
  wire [0:0] v_16506;
  wire [0:0] v_16507;
  function [0:0] mux_16507(input [0:0] sel);
    case (sel) 0: mux_16507 = 1'h0; 1: mux_16507 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16508;
  function [0:0] mux_16508(input [0:0] sel);
    case (sel) 0: mux_16508 = 1'h0; 1: mux_16508 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16509;
  wire [0:0] v_16510;
  wire [0:0] v_16511;
  wire [0:0] v_16512;
  wire [0:0] v_16513;
  wire [0:0] v_16514;
  wire [0:0] v_16515;
  function [0:0] mux_16515(input [0:0] sel);
    case (sel) 0: mux_16515 = 1'h0; 1: mux_16515 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16516;
  wire [0:0] v_16517;
  wire [0:0] v_16518;
  wire [0:0] v_16519;
  wire [0:0] v_16520;
  function [0:0] mux_16520(input [0:0] sel);
    case (sel) 0: mux_16520 = 1'h0; 1: mux_16520 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16521;
  wire [0:0] v_16522;
  wire [0:0] v_16523;
  wire [0:0] v_16524;
  function [0:0] mux_16524(input [0:0] sel);
    case (sel) 0: mux_16524 = 1'h0; 1: mux_16524 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16525;
  function [0:0] mux_16525(input [0:0] sel);
    case (sel) 0: mux_16525 = 1'h0; 1: mux_16525 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_16526 = 1'h0;
  wire [0:0] v_16527;
  wire [0:0] v_16528;
  wire [0:0] act_16529;
  wire [0:0] v_16530;
  wire [0:0] v_16531;
  wire [0:0] v_16532;
  wire [0:0] vin0_consume_en_16533;
  wire [0:0] vout_canPeek_16533;
  wire [7:0] vout_peek_16533;
  wire [0:0] v_16534;
  wire [0:0] v_16535;
  function [0:0] mux_16535(input [0:0] sel);
    case (sel) 0: mux_16535 = 1'h0; 1: mux_16535 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16536;
  wire [0:0] v_16537;
  wire [0:0] v_16538;
  wire [0:0] v_16539;
  wire [0:0] v_16540;
  function [0:0] mux_16540(input [0:0] sel);
    case (sel) 0: mux_16540 = 1'h0; 1: mux_16540 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16541;
  wire [0:0] vin0_consume_en_16542;
  wire [0:0] vout_canPeek_16542;
  wire [7:0] vout_peek_16542;
  wire [0:0] v_16543;
  wire [0:0] v_16544;
  function [0:0] mux_16544(input [0:0] sel);
    case (sel) 0: mux_16544 = 1'h0; 1: mux_16544 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16545;
  function [0:0] mux_16545(input [0:0] sel);
    case (sel) 0: mux_16545 = 1'h0; 1: mux_16545 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16546;
  wire [0:0] v_16547;
  wire [0:0] v_16548;
  wire [0:0] v_16549;
  wire [0:0] v_16550;
  wire [0:0] v_16551;
  wire [0:0] v_16552;
  function [0:0] mux_16552(input [0:0] sel);
    case (sel) 0: mux_16552 = 1'h0; 1: mux_16552 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16553;
  function [0:0] mux_16553(input [0:0] sel);
    case (sel) 0: mux_16553 = 1'h0; 1: mux_16553 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16554;
  wire [0:0] v_16555;
  wire [0:0] v_16556;
  wire [0:0] v_16557;
  function [0:0] mux_16557(input [0:0] sel);
    case (sel) 0: mux_16557 = 1'h0; 1: mux_16557 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16558;
  function [0:0] mux_16558(input [0:0] sel);
    case (sel) 0: mux_16558 = 1'h0; 1: mux_16558 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16559;
  wire [0:0] v_16560;
  wire [0:0] v_16561;
  wire [0:0] v_16562;
  wire [0:0] v_16563;
  wire [0:0] v_16564;
  function [0:0] mux_16564(input [0:0] sel);
    case (sel) 0: mux_16564 = 1'h0; 1: mux_16564 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16565;
  wire [0:0] v_16566;
  wire [0:0] v_16567;
  wire [0:0] v_16568;
  wire [0:0] v_16569;
  function [0:0] mux_16569(input [0:0] sel);
    case (sel) 0: mux_16569 = 1'h0; 1: mux_16569 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16570;
  wire [0:0] v_16571;
  wire [0:0] v_16572;
  wire [0:0] v_16573;
  function [0:0] mux_16573(input [0:0] sel);
    case (sel) 0: mux_16573 = 1'h0; 1: mux_16573 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16574;
  function [0:0] mux_16574(input [0:0] sel);
    case (sel) 0: mux_16574 = 1'h0; 1: mux_16574 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_16575 = 1'h0;
  wire [0:0] v_16576;
  wire [0:0] v_16577;
  wire [0:0] act_16578;
  wire [0:0] v_16579;
  wire [0:0] v_16580;
  wire [0:0] v_16581;
  reg [0:0] v_16582 = 1'h0;
  wire [0:0] v_16583;
  wire [0:0] v_16584;
  wire [0:0] act_16585;
  wire [0:0] v_16586;
  wire [0:0] v_16587;
  wire [0:0] v_16588;
  wire [0:0] vin0_consume_en_16589;
  wire [0:0] vout_canPeek_16589;
  wire [7:0] vout_peek_16589;
  wire [0:0] v_16590;
  wire [0:0] v_16591;
  function [0:0] mux_16591(input [0:0] sel);
    case (sel) 0: mux_16591 = 1'h0; 1: mux_16591 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16592;
  wire [0:0] v_16593;
  wire [0:0] v_16594;
  wire [0:0] v_16595;
  wire [0:0] v_16596;
  function [0:0] mux_16596(input [0:0] sel);
    case (sel) 0: mux_16596 = 1'h0; 1: mux_16596 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16597;
  wire [0:0] vin0_consume_en_16598;
  wire [0:0] vout_canPeek_16598;
  wire [7:0] vout_peek_16598;
  wire [0:0] v_16599;
  wire [0:0] v_16600;
  function [0:0] mux_16600(input [0:0] sel);
    case (sel) 0: mux_16600 = 1'h0; 1: mux_16600 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16601;
  function [0:0] mux_16601(input [0:0] sel);
    case (sel) 0: mux_16601 = 1'h0; 1: mux_16601 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16602;
  wire [0:0] v_16603;
  wire [0:0] v_16604;
  wire [0:0] v_16605;
  wire [0:0] v_16606;
  wire [0:0] v_16607;
  wire [0:0] v_16608;
  function [0:0] mux_16608(input [0:0] sel);
    case (sel) 0: mux_16608 = 1'h0; 1: mux_16608 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16609;
  wire [0:0] v_16610;
  wire [0:0] v_16611;
  wire [0:0] v_16612;
  wire [0:0] v_16613;
  function [0:0] mux_16613(input [0:0] sel);
    case (sel) 0: mux_16613 = 1'h0; 1: mux_16613 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16614;
  wire [0:0] v_16615;
  wire [0:0] v_16616;
  wire [0:0] v_16617;
  function [0:0] mux_16617(input [0:0] sel);
    case (sel) 0: mux_16617 = 1'h0; 1: mux_16617 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16618;
  function [0:0] mux_16618(input [0:0] sel);
    case (sel) 0: mux_16618 = 1'h0; 1: mux_16618 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_16619 = 1'h0;
  wire [0:0] v_16620;
  wire [0:0] v_16621;
  wire [0:0] act_16622;
  wire [0:0] v_16623;
  wire [0:0] v_16624;
  wire [0:0] v_16625;
  wire [0:0] vin0_consume_en_16626;
  wire [0:0] vout_canPeek_16626;
  wire [7:0] vout_peek_16626;
  wire [0:0] v_16627;
  wire [0:0] v_16628;
  function [0:0] mux_16628(input [0:0] sel);
    case (sel) 0: mux_16628 = 1'h0; 1: mux_16628 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16629;
  wire [0:0] v_16630;
  wire [0:0] v_16631;
  wire [0:0] v_16632;
  wire [0:0] v_16633;
  function [0:0] mux_16633(input [0:0] sel);
    case (sel) 0: mux_16633 = 1'h0; 1: mux_16633 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16634;
  wire [0:0] vin0_consume_en_16635;
  wire [0:0] vout_canPeek_16635;
  wire [7:0] vout_peek_16635;
  wire [0:0] v_16636;
  wire [0:0] v_16637;
  function [0:0] mux_16637(input [0:0] sel);
    case (sel) 0: mux_16637 = 1'h0; 1: mux_16637 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16638;
  function [0:0] mux_16638(input [0:0] sel);
    case (sel) 0: mux_16638 = 1'h0; 1: mux_16638 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16639;
  wire [0:0] v_16640;
  wire [0:0] v_16641;
  wire [0:0] v_16642;
  wire [0:0] v_16643;
  wire [0:0] v_16644;
  wire [0:0] v_16645;
  function [0:0] mux_16645(input [0:0] sel);
    case (sel) 0: mux_16645 = 1'h0; 1: mux_16645 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16646;
  function [0:0] mux_16646(input [0:0] sel);
    case (sel) 0: mux_16646 = 1'h0; 1: mux_16646 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16647;
  wire [0:0] v_16648;
  wire [0:0] v_16649;
  wire [0:0] v_16650;
  function [0:0] mux_16650(input [0:0] sel);
    case (sel) 0: mux_16650 = 1'h0; 1: mux_16650 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16651;
  function [0:0] mux_16651(input [0:0] sel);
    case (sel) 0: mux_16651 = 1'h0; 1: mux_16651 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16652;
  wire [0:0] v_16653;
  wire [0:0] v_16654;
  wire [0:0] v_16655;
  wire [0:0] v_16656;
  wire [0:0] v_16657;
  function [0:0] mux_16657(input [0:0] sel);
    case (sel) 0: mux_16657 = 1'h0; 1: mux_16657 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16658;
  function [0:0] mux_16658(input [0:0] sel);
    case (sel) 0: mux_16658 = 1'h0; 1: mux_16658 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16659;
  wire [0:0] v_16660;
  wire [0:0] v_16661;
  wire [0:0] v_16662;
  function [0:0] mux_16662(input [0:0] sel);
    case (sel) 0: mux_16662 = 1'h0; 1: mux_16662 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16663;
  function [0:0] mux_16663(input [0:0] sel);
    case (sel) 0: mux_16663 = 1'h0; 1: mux_16663 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16664;
  wire [0:0] v_16665;
  wire [0:0] v_16666;
  wire [0:0] v_16667;
  wire [0:0] v_16668;
  wire [0:0] v_16669;
  function [0:0] mux_16669(input [0:0] sel);
    case (sel) 0: mux_16669 = 1'h0; 1: mux_16669 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16670;
  wire [0:0] v_16671;
  wire [0:0] v_16672;
  wire [0:0] v_16673;
  wire [0:0] v_16674;
  function [0:0] mux_16674(input [0:0] sel);
    case (sel) 0: mux_16674 = 1'h0; 1: mux_16674 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16675;
  wire [0:0] v_16676;
  wire [0:0] v_16677;
  wire [0:0] v_16678;
  function [0:0] mux_16678(input [0:0] sel);
    case (sel) 0: mux_16678 = 1'h0; 1: mux_16678 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16679;
  function [0:0] mux_16679(input [0:0] sel);
    case (sel) 0: mux_16679 = 1'h0; 1: mux_16679 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_16680 = 1'h0;
  wire [0:0] v_16681;
  wire [0:0] v_16682;
  wire [0:0] act_16683;
  wire [0:0] v_16684;
  wire [0:0] v_16685;
  wire [0:0] v_16686;
  reg [0:0] v_16687 = 1'h0;
  wire [0:0] v_16688;
  wire [0:0] v_16689;
  wire [0:0] act_16690;
  wire [0:0] v_16691;
  wire [0:0] v_16692;
  wire [0:0] v_16693;
  reg [0:0] v_16694 = 1'h0;
  wire [0:0] v_16695;
  wire [0:0] v_16696;
  wire [0:0] act_16697;
  wire [0:0] v_16698;
  wire [0:0] v_16699;
  wire [0:0] v_16700;
  wire [0:0] vin0_consume_en_16701;
  wire [0:0] vout_canPeek_16701;
  wire [7:0] vout_peek_16701;
  wire [0:0] v_16702;
  wire [0:0] v_16703;
  function [0:0] mux_16703(input [0:0] sel);
    case (sel) 0: mux_16703 = 1'h0; 1: mux_16703 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16704;
  wire [0:0] v_16705;
  wire [0:0] v_16706;
  wire [0:0] v_16707;
  wire [0:0] v_16708;
  function [0:0] mux_16708(input [0:0] sel);
    case (sel) 0: mux_16708 = 1'h0; 1: mux_16708 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16709;
  wire [0:0] vin0_consume_en_16710;
  wire [0:0] vout_canPeek_16710;
  wire [7:0] vout_peek_16710;
  wire [0:0] v_16711;
  wire [0:0] v_16712;
  function [0:0] mux_16712(input [0:0] sel);
    case (sel) 0: mux_16712 = 1'h0; 1: mux_16712 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16713;
  function [0:0] mux_16713(input [0:0] sel);
    case (sel) 0: mux_16713 = 1'h0; 1: mux_16713 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16714;
  wire [0:0] v_16715;
  wire [0:0] v_16716;
  wire [0:0] v_16717;
  wire [0:0] v_16718;
  wire [0:0] v_16719;
  wire [0:0] v_16720;
  function [0:0] mux_16720(input [0:0] sel);
    case (sel) 0: mux_16720 = 1'h0; 1: mux_16720 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16721;
  wire [0:0] v_16722;
  wire [0:0] v_16723;
  wire [0:0] v_16724;
  wire [0:0] v_16725;
  function [0:0] mux_16725(input [0:0] sel);
    case (sel) 0: mux_16725 = 1'h0; 1: mux_16725 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16726;
  wire [0:0] v_16727;
  wire [0:0] v_16728;
  wire [0:0] v_16729;
  function [0:0] mux_16729(input [0:0] sel);
    case (sel) 0: mux_16729 = 1'h0; 1: mux_16729 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16730;
  function [0:0] mux_16730(input [0:0] sel);
    case (sel) 0: mux_16730 = 1'h0; 1: mux_16730 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_16731 = 1'h0;
  wire [0:0] v_16732;
  wire [0:0] v_16733;
  wire [0:0] act_16734;
  wire [0:0] v_16735;
  wire [0:0] v_16736;
  wire [0:0] v_16737;
  wire [0:0] vin0_consume_en_16738;
  wire [0:0] vout_canPeek_16738;
  wire [7:0] vout_peek_16738;
  wire [0:0] v_16739;
  wire [0:0] v_16740;
  function [0:0] mux_16740(input [0:0] sel);
    case (sel) 0: mux_16740 = 1'h0; 1: mux_16740 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16741;
  wire [0:0] v_16742;
  wire [0:0] v_16743;
  wire [0:0] v_16744;
  wire [0:0] v_16745;
  function [0:0] mux_16745(input [0:0] sel);
    case (sel) 0: mux_16745 = 1'h0; 1: mux_16745 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16746;
  wire [0:0] vin0_consume_en_16747;
  wire [0:0] vout_canPeek_16747;
  wire [7:0] vout_peek_16747;
  wire [0:0] v_16748;
  wire [0:0] v_16749;
  function [0:0] mux_16749(input [0:0] sel);
    case (sel) 0: mux_16749 = 1'h0; 1: mux_16749 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16750;
  function [0:0] mux_16750(input [0:0] sel);
    case (sel) 0: mux_16750 = 1'h0; 1: mux_16750 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16751;
  wire [0:0] v_16752;
  wire [0:0] v_16753;
  wire [0:0] v_16754;
  wire [0:0] v_16755;
  wire [0:0] v_16756;
  wire [0:0] v_16757;
  function [0:0] mux_16757(input [0:0] sel);
    case (sel) 0: mux_16757 = 1'h0; 1: mux_16757 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16758;
  function [0:0] mux_16758(input [0:0] sel);
    case (sel) 0: mux_16758 = 1'h0; 1: mux_16758 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16759;
  wire [0:0] v_16760;
  wire [0:0] v_16761;
  wire [0:0] v_16762;
  function [0:0] mux_16762(input [0:0] sel);
    case (sel) 0: mux_16762 = 1'h0; 1: mux_16762 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16763;
  function [0:0] mux_16763(input [0:0] sel);
    case (sel) 0: mux_16763 = 1'h0; 1: mux_16763 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16764;
  wire [0:0] v_16765;
  wire [0:0] v_16766;
  wire [0:0] v_16767;
  wire [0:0] v_16768;
  wire [0:0] v_16769;
  function [0:0] mux_16769(input [0:0] sel);
    case (sel) 0: mux_16769 = 1'h0; 1: mux_16769 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16770;
  wire [0:0] v_16771;
  wire [0:0] v_16772;
  wire [0:0] v_16773;
  wire [0:0] v_16774;
  function [0:0] mux_16774(input [0:0] sel);
    case (sel) 0: mux_16774 = 1'h0; 1: mux_16774 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16775;
  wire [0:0] v_16776;
  wire [0:0] v_16777;
  wire [0:0] v_16778;
  function [0:0] mux_16778(input [0:0] sel);
    case (sel) 0: mux_16778 = 1'h0; 1: mux_16778 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16779;
  function [0:0] mux_16779(input [0:0] sel);
    case (sel) 0: mux_16779 = 1'h0; 1: mux_16779 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_16780 = 1'h0;
  wire [0:0] v_16781;
  wire [0:0] v_16782;
  wire [0:0] act_16783;
  wire [0:0] v_16784;
  wire [0:0] v_16785;
  wire [0:0] v_16786;
  reg [0:0] v_16787 = 1'h0;
  wire [0:0] v_16788;
  wire [0:0] v_16789;
  wire [0:0] act_16790;
  wire [0:0] v_16791;
  wire [0:0] v_16792;
  wire [0:0] v_16793;
  wire [0:0] vin0_consume_en_16794;
  wire [0:0] vout_canPeek_16794;
  wire [7:0] vout_peek_16794;
  wire [0:0] v_16795;
  wire [0:0] v_16796;
  function [0:0] mux_16796(input [0:0] sel);
    case (sel) 0: mux_16796 = 1'h0; 1: mux_16796 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16797;
  wire [0:0] v_16798;
  wire [0:0] v_16799;
  wire [0:0] v_16800;
  wire [0:0] v_16801;
  function [0:0] mux_16801(input [0:0] sel);
    case (sel) 0: mux_16801 = 1'h0; 1: mux_16801 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16802;
  wire [0:0] vin0_consume_en_16803;
  wire [0:0] vout_canPeek_16803;
  wire [7:0] vout_peek_16803;
  wire [0:0] v_16804;
  wire [0:0] v_16805;
  function [0:0] mux_16805(input [0:0] sel);
    case (sel) 0: mux_16805 = 1'h0; 1: mux_16805 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16806;
  function [0:0] mux_16806(input [0:0] sel);
    case (sel) 0: mux_16806 = 1'h0; 1: mux_16806 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16807;
  wire [0:0] v_16808;
  wire [0:0] v_16809;
  wire [0:0] v_16810;
  wire [0:0] v_16811;
  wire [0:0] v_16812;
  wire [0:0] v_16813;
  function [0:0] mux_16813(input [0:0] sel);
    case (sel) 0: mux_16813 = 1'h0; 1: mux_16813 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16814;
  wire [0:0] v_16815;
  wire [0:0] v_16816;
  wire [0:0] v_16817;
  wire [0:0] v_16818;
  function [0:0] mux_16818(input [0:0] sel);
    case (sel) 0: mux_16818 = 1'h0; 1: mux_16818 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16819;
  wire [0:0] v_16820;
  wire [0:0] v_16821;
  wire [0:0] v_16822;
  function [0:0] mux_16822(input [0:0] sel);
    case (sel) 0: mux_16822 = 1'h0; 1: mux_16822 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16823;
  function [0:0] mux_16823(input [0:0] sel);
    case (sel) 0: mux_16823 = 1'h0; 1: mux_16823 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_16824 = 1'h0;
  wire [0:0] v_16825;
  wire [0:0] v_16826;
  wire [0:0] act_16827;
  wire [0:0] v_16828;
  wire [0:0] v_16829;
  wire [0:0] v_16830;
  wire [0:0] vin0_consume_en_16831;
  wire [0:0] vout_canPeek_16831;
  wire [7:0] vout_peek_16831;
  wire [0:0] v_16832;
  wire [0:0] v_16833;
  function [0:0] mux_16833(input [0:0] sel);
    case (sel) 0: mux_16833 = 1'h0; 1: mux_16833 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16834;
  wire [0:0] v_16835;
  wire [0:0] v_16836;
  wire [0:0] v_16837;
  wire [0:0] v_16838;
  function [0:0] mux_16838(input [0:0] sel);
    case (sel) 0: mux_16838 = 1'h0; 1: mux_16838 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16839;
  wire [0:0] vin0_consume_en_16840;
  wire [0:0] vout_canPeek_16840;
  wire [7:0] vout_peek_16840;
  wire [0:0] v_16841;
  wire [0:0] v_16842;
  function [0:0] mux_16842(input [0:0] sel);
    case (sel) 0: mux_16842 = 1'h0; 1: mux_16842 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16843;
  function [0:0] mux_16843(input [0:0] sel);
    case (sel) 0: mux_16843 = 1'h0; 1: mux_16843 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16844;
  wire [0:0] v_16845;
  wire [0:0] v_16846;
  wire [0:0] v_16847;
  wire [0:0] v_16848;
  wire [0:0] v_16849;
  wire [0:0] v_16850;
  function [0:0] mux_16850(input [0:0] sel);
    case (sel) 0: mux_16850 = 1'h0; 1: mux_16850 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16851;
  function [0:0] mux_16851(input [0:0] sel);
    case (sel) 0: mux_16851 = 1'h0; 1: mux_16851 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16852;
  wire [0:0] v_16853;
  wire [0:0] v_16854;
  wire [0:0] v_16855;
  function [0:0] mux_16855(input [0:0] sel);
    case (sel) 0: mux_16855 = 1'h0; 1: mux_16855 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16856;
  function [0:0] mux_16856(input [0:0] sel);
    case (sel) 0: mux_16856 = 1'h0; 1: mux_16856 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16857;
  wire [0:0] v_16858;
  wire [0:0] v_16859;
  wire [0:0] v_16860;
  wire [0:0] v_16861;
  wire [0:0] v_16862;
  function [0:0] mux_16862(input [0:0] sel);
    case (sel) 0: mux_16862 = 1'h0; 1: mux_16862 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16863;
  function [0:0] mux_16863(input [0:0] sel);
    case (sel) 0: mux_16863 = 1'h0; 1: mux_16863 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16864;
  wire [0:0] v_16865;
  wire [0:0] v_16866;
  wire [0:0] v_16867;
  function [0:0] mux_16867(input [0:0] sel);
    case (sel) 0: mux_16867 = 1'h0; 1: mux_16867 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16868;
  function [0:0] mux_16868(input [0:0] sel);
    case (sel) 0: mux_16868 = 1'h0; 1: mux_16868 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16869;
  wire [0:0] v_16870;
  wire [0:0] v_16871;
  wire [0:0] v_16872;
  wire [0:0] v_16873;
  wire [0:0] v_16874;
  function [0:0] mux_16874(input [0:0] sel);
    case (sel) 0: mux_16874 = 1'h0; 1: mux_16874 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16875;
  function [0:0] mux_16875(input [0:0] sel);
    case (sel) 0: mux_16875 = 1'h0; 1: mux_16875 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16876;
  wire [0:0] v_16877;
  wire [0:0] v_16878;
  wire [0:0] v_16879;
  function [0:0] mux_16879(input [0:0] sel);
    case (sel) 0: mux_16879 = 1'h0; 1: mux_16879 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16880;
  function [0:0] mux_16880(input [0:0] sel);
    case (sel) 0: mux_16880 = 1'h0; 1: mux_16880 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16881;
  wire [0:0] v_16882;
  wire [0:0] v_16883;
  wire [0:0] v_16884;
  wire [0:0] v_16885;
  wire [0:0] v_16886;
  function [0:0] mux_16886(input [0:0] sel);
    case (sel) 0: mux_16886 = 1'h0; 1: mux_16886 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16887;
  function [0:0] mux_16887(input [0:0] sel);
    case (sel) 0: mux_16887 = 1'h0; 1: mux_16887 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16888;
  wire [0:0] v_16889;
  wire [0:0] v_16890;
  wire [0:0] v_16891;
  function [0:0] mux_16891(input [0:0] sel);
    case (sel) 0: mux_16891 = 1'h0; 1: mux_16891 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16892;
  function [0:0] mux_16892(input [0:0] sel);
    case (sel) 0: mux_16892 = 1'h0; 1: mux_16892 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16893;
  wire [0:0] v_16894;
  wire [0:0] v_16895;
  wire [0:0] v_16896;
  wire [0:0] v_16897;
  wire [0:0] v_16898;
  function [0:0] mux_16898(input [0:0] sel);
    case (sel) 0: mux_16898 = 1'h0; 1: mux_16898 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16899;
  function [0:0] mux_16899(input [0:0] sel);
    case (sel) 0: mux_16899 = 1'h0; 1: mux_16899 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16900;
  wire [0:0] v_16901;
  wire [0:0] v_16902;
  wire [0:0] v_16903;
  function [0:0] mux_16903(input [0:0] sel);
    case (sel) 0: mux_16903 = 1'h0; 1: mux_16903 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16904;
  function [0:0] mux_16904(input [0:0] sel);
    case (sel) 0: mux_16904 = 1'h0; 1: mux_16904 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16905;
  wire [0:0] v_16906;
  wire [0:0] v_16907;
  wire [0:0] v_16908;
  wire [0:0] v_16909;
  wire [0:0] v_16910;
  function [0:0] mux_16910(input [0:0] sel);
    case (sel) 0: mux_16910 = 1'h0; 1: mux_16910 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16911;
  wire [0:0] v_16912;
  wire [0:0] v_16913;
  wire [0:0] v_16914;
  wire [0:0] v_16915;
  function [0:0] mux_16915(input [0:0] sel);
    case (sel) 0: mux_16915 = 1'h0; 1: mux_16915 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16916;
  wire [0:0] v_16917;
  wire [0:0] v_16918;
  wire [0:0] v_16919;
  function [0:0] mux_16919(input [0:0] sel);
    case (sel) 0: mux_16919 = 1'h0; 1: mux_16919 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16920;
  function [0:0] mux_16920(input [0:0] sel);
    case (sel) 0: mux_16920 = 1'h0; 1: mux_16920 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_16921 = 1'h0;
  wire [0:0] v_16922;
  wire [0:0] v_16923;
  wire [0:0] act_16924;
  wire [0:0] v_16925;
  wire [0:0] v_16926;
  wire [0:0] v_16927;
  reg [0:0] v_16928 = 1'h0;
  wire [0:0] v_16929;
  wire [0:0] v_16930;
  wire [0:0] act_16931;
  wire [0:0] v_16932;
  wire [0:0] v_16933;
  wire [0:0] v_16934;
  reg [0:0] v_16935 = 1'h0;
  wire [0:0] v_16936;
  wire [0:0] v_16937;
  wire [0:0] act_16938;
  wire [0:0] v_16939;
  wire [0:0] v_16940;
  wire [0:0] v_16941;
  reg [0:0] v_16942 = 1'h0;
  wire [0:0] v_16943;
  wire [0:0] v_16944;
  wire [0:0] act_16945;
  wire [0:0] v_16946;
  wire [0:0] v_16947;
  wire [0:0] v_16948;
  reg [0:0] v_16949 = 1'h0;
  wire [0:0] v_16950;
  wire [0:0] v_16951;
  wire [0:0] act_16952;
  wire [0:0] v_16953;
  wire [0:0] v_16954;
  wire [0:0] v_16955;
  reg [0:0] v_16956 = 1'h0;
  wire [0:0] v_16957;
  wire [0:0] v_16958;
  wire [0:0] act_16959;
  wire [0:0] v_16960;
  wire [0:0] v_16961;
  wire [0:0] v_16962;
  wire [0:0] vin0_consume_en_16963;
  wire [0:0] vout_canPeek_16963;
  wire [7:0] vout_peek_16963;
  wire [0:0] v_16964;
  wire [0:0] v_16965;
  function [0:0] mux_16965(input [0:0] sel);
    case (sel) 0: mux_16965 = 1'h0; 1: mux_16965 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16966;
  wire [0:0] v_16967;
  wire [0:0] v_16968;
  wire [0:0] v_16969;
  wire [0:0] v_16970;
  function [0:0] mux_16970(input [0:0] sel);
    case (sel) 0: mux_16970 = 1'h0; 1: mux_16970 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16971;
  wire [0:0] vin0_consume_en_16972;
  wire [0:0] vout_canPeek_16972;
  wire [7:0] vout_peek_16972;
  wire [0:0] v_16973;
  wire [0:0] v_16974;
  function [0:0] mux_16974(input [0:0] sel);
    case (sel) 0: mux_16974 = 1'h0; 1: mux_16974 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16975;
  function [0:0] mux_16975(input [0:0] sel);
    case (sel) 0: mux_16975 = 1'h0; 1: mux_16975 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16976;
  wire [0:0] v_16977;
  wire [0:0] v_16978;
  wire [0:0] v_16979;
  wire [0:0] v_16980;
  wire [0:0] v_16981;
  wire [0:0] v_16982;
  function [0:0] mux_16982(input [0:0] sel);
    case (sel) 0: mux_16982 = 1'h0; 1: mux_16982 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16983;
  wire [0:0] v_16984;
  wire [0:0] v_16985;
  wire [0:0] v_16986;
  wire [0:0] v_16987;
  function [0:0] mux_16987(input [0:0] sel);
    case (sel) 0: mux_16987 = 1'h0; 1: mux_16987 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_16988;
  wire [0:0] v_16989;
  wire [0:0] v_16990;
  wire [0:0] v_16991;
  function [0:0] mux_16991(input [0:0] sel);
    case (sel) 0: mux_16991 = 1'h0; 1: mux_16991 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16992;
  function [0:0] mux_16992(input [0:0] sel);
    case (sel) 0: mux_16992 = 1'h0; 1: mux_16992 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_16993 = 1'h0;
  wire [0:0] v_16994;
  wire [0:0] v_16995;
  wire [0:0] act_16996;
  wire [0:0] v_16997;
  wire [0:0] v_16998;
  wire [0:0] v_16999;
  wire [0:0] vin0_consume_en_17000;
  wire [0:0] vout_canPeek_17000;
  wire [7:0] vout_peek_17000;
  wire [0:0] v_17001;
  wire [0:0] v_17002;
  function [0:0] mux_17002(input [0:0] sel);
    case (sel) 0: mux_17002 = 1'h0; 1: mux_17002 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17003;
  wire [0:0] v_17004;
  wire [0:0] v_17005;
  wire [0:0] v_17006;
  wire [0:0] v_17007;
  function [0:0] mux_17007(input [0:0] sel);
    case (sel) 0: mux_17007 = 1'h0; 1: mux_17007 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17008;
  wire [0:0] vin0_consume_en_17009;
  wire [0:0] vout_canPeek_17009;
  wire [7:0] vout_peek_17009;
  wire [0:0] v_17010;
  wire [0:0] v_17011;
  function [0:0] mux_17011(input [0:0] sel);
    case (sel) 0: mux_17011 = 1'h0; 1: mux_17011 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17012;
  function [0:0] mux_17012(input [0:0] sel);
    case (sel) 0: mux_17012 = 1'h0; 1: mux_17012 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17013;
  wire [0:0] v_17014;
  wire [0:0] v_17015;
  wire [0:0] v_17016;
  wire [0:0] v_17017;
  wire [0:0] v_17018;
  wire [0:0] v_17019;
  function [0:0] mux_17019(input [0:0] sel);
    case (sel) 0: mux_17019 = 1'h0; 1: mux_17019 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17020;
  function [0:0] mux_17020(input [0:0] sel);
    case (sel) 0: mux_17020 = 1'h0; 1: mux_17020 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17021;
  wire [0:0] v_17022;
  wire [0:0] v_17023;
  wire [0:0] v_17024;
  function [0:0] mux_17024(input [0:0] sel);
    case (sel) 0: mux_17024 = 1'h0; 1: mux_17024 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17025;
  function [0:0] mux_17025(input [0:0] sel);
    case (sel) 0: mux_17025 = 1'h0; 1: mux_17025 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17026;
  wire [0:0] v_17027;
  wire [0:0] v_17028;
  wire [0:0] v_17029;
  wire [0:0] v_17030;
  wire [0:0] v_17031;
  function [0:0] mux_17031(input [0:0] sel);
    case (sel) 0: mux_17031 = 1'h0; 1: mux_17031 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17032;
  wire [0:0] v_17033;
  wire [0:0] v_17034;
  wire [0:0] v_17035;
  wire [0:0] v_17036;
  function [0:0] mux_17036(input [0:0] sel);
    case (sel) 0: mux_17036 = 1'h0; 1: mux_17036 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17037;
  wire [0:0] v_17038;
  wire [0:0] v_17039;
  wire [0:0] v_17040;
  function [0:0] mux_17040(input [0:0] sel);
    case (sel) 0: mux_17040 = 1'h0; 1: mux_17040 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17041;
  function [0:0] mux_17041(input [0:0] sel);
    case (sel) 0: mux_17041 = 1'h0; 1: mux_17041 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_17042 = 1'h0;
  wire [0:0] v_17043;
  wire [0:0] v_17044;
  wire [0:0] act_17045;
  wire [0:0] v_17046;
  wire [0:0] v_17047;
  wire [0:0] v_17048;
  reg [0:0] v_17049 = 1'h0;
  wire [0:0] v_17050;
  wire [0:0] v_17051;
  wire [0:0] act_17052;
  wire [0:0] v_17053;
  wire [0:0] v_17054;
  wire [0:0] v_17055;
  wire [0:0] vin0_consume_en_17056;
  wire [0:0] vout_canPeek_17056;
  wire [7:0] vout_peek_17056;
  wire [0:0] v_17057;
  wire [0:0] v_17058;
  function [0:0] mux_17058(input [0:0] sel);
    case (sel) 0: mux_17058 = 1'h0; 1: mux_17058 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17059;
  wire [0:0] v_17060;
  wire [0:0] v_17061;
  wire [0:0] v_17062;
  wire [0:0] v_17063;
  function [0:0] mux_17063(input [0:0] sel);
    case (sel) 0: mux_17063 = 1'h0; 1: mux_17063 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17064;
  wire [0:0] vin0_consume_en_17065;
  wire [0:0] vout_canPeek_17065;
  wire [7:0] vout_peek_17065;
  wire [0:0] v_17066;
  wire [0:0] v_17067;
  function [0:0] mux_17067(input [0:0] sel);
    case (sel) 0: mux_17067 = 1'h0; 1: mux_17067 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17068;
  function [0:0] mux_17068(input [0:0] sel);
    case (sel) 0: mux_17068 = 1'h0; 1: mux_17068 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17069;
  wire [0:0] v_17070;
  wire [0:0] v_17071;
  wire [0:0] v_17072;
  wire [0:0] v_17073;
  wire [0:0] v_17074;
  wire [0:0] v_17075;
  function [0:0] mux_17075(input [0:0] sel);
    case (sel) 0: mux_17075 = 1'h0; 1: mux_17075 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17076;
  wire [0:0] v_17077;
  wire [0:0] v_17078;
  wire [0:0] v_17079;
  wire [0:0] v_17080;
  function [0:0] mux_17080(input [0:0] sel);
    case (sel) 0: mux_17080 = 1'h0; 1: mux_17080 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17081;
  wire [0:0] v_17082;
  wire [0:0] v_17083;
  wire [0:0] v_17084;
  function [0:0] mux_17084(input [0:0] sel);
    case (sel) 0: mux_17084 = 1'h0; 1: mux_17084 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17085;
  function [0:0] mux_17085(input [0:0] sel);
    case (sel) 0: mux_17085 = 1'h0; 1: mux_17085 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_17086 = 1'h0;
  wire [0:0] v_17087;
  wire [0:0] v_17088;
  wire [0:0] act_17089;
  wire [0:0] v_17090;
  wire [0:0] v_17091;
  wire [0:0] v_17092;
  wire [0:0] vin0_consume_en_17093;
  wire [0:0] vout_canPeek_17093;
  wire [7:0] vout_peek_17093;
  wire [0:0] v_17094;
  wire [0:0] v_17095;
  function [0:0] mux_17095(input [0:0] sel);
    case (sel) 0: mux_17095 = 1'h0; 1: mux_17095 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17096;
  wire [0:0] v_17097;
  wire [0:0] v_17098;
  wire [0:0] v_17099;
  wire [0:0] v_17100;
  function [0:0] mux_17100(input [0:0] sel);
    case (sel) 0: mux_17100 = 1'h0; 1: mux_17100 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17101;
  wire [0:0] vin0_consume_en_17102;
  wire [0:0] vout_canPeek_17102;
  wire [7:0] vout_peek_17102;
  wire [0:0] v_17103;
  wire [0:0] v_17104;
  function [0:0] mux_17104(input [0:0] sel);
    case (sel) 0: mux_17104 = 1'h0; 1: mux_17104 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17105;
  function [0:0] mux_17105(input [0:0] sel);
    case (sel) 0: mux_17105 = 1'h0; 1: mux_17105 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17106;
  wire [0:0] v_17107;
  wire [0:0] v_17108;
  wire [0:0] v_17109;
  wire [0:0] v_17110;
  wire [0:0] v_17111;
  wire [0:0] v_17112;
  function [0:0] mux_17112(input [0:0] sel);
    case (sel) 0: mux_17112 = 1'h0; 1: mux_17112 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17113;
  function [0:0] mux_17113(input [0:0] sel);
    case (sel) 0: mux_17113 = 1'h0; 1: mux_17113 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17114;
  wire [0:0] v_17115;
  wire [0:0] v_17116;
  wire [0:0] v_17117;
  function [0:0] mux_17117(input [0:0] sel);
    case (sel) 0: mux_17117 = 1'h0; 1: mux_17117 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17118;
  function [0:0] mux_17118(input [0:0] sel);
    case (sel) 0: mux_17118 = 1'h0; 1: mux_17118 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17119;
  wire [0:0] v_17120;
  wire [0:0] v_17121;
  wire [0:0] v_17122;
  wire [0:0] v_17123;
  wire [0:0] v_17124;
  function [0:0] mux_17124(input [0:0] sel);
    case (sel) 0: mux_17124 = 1'h0; 1: mux_17124 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17125;
  function [0:0] mux_17125(input [0:0] sel);
    case (sel) 0: mux_17125 = 1'h0; 1: mux_17125 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17126;
  wire [0:0] v_17127;
  wire [0:0] v_17128;
  wire [0:0] v_17129;
  function [0:0] mux_17129(input [0:0] sel);
    case (sel) 0: mux_17129 = 1'h0; 1: mux_17129 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17130;
  function [0:0] mux_17130(input [0:0] sel);
    case (sel) 0: mux_17130 = 1'h0; 1: mux_17130 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17131;
  wire [0:0] v_17132;
  wire [0:0] v_17133;
  wire [0:0] v_17134;
  wire [0:0] v_17135;
  wire [0:0] v_17136;
  function [0:0] mux_17136(input [0:0] sel);
    case (sel) 0: mux_17136 = 1'h0; 1: mux_17136 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17137;
  wire [0:0] v_17138;
  wire [0:0] v_17139;
  wire [0:0] v_17140;
  wire [0:0] v_17141;
  function [0:0] mux_17141(input [0:0] sel);
    case (sel) 0: mux_17141 = 1'h0; 1: mux_17141 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17142;
  wire [0:0] v_17143;
  wire [0:0] v_17144;
  wire [0:0] v_17145;
  function [0:0] mux_17145(input [0:0] sel);
    case (sel) 0: mux_17145 = 1'h0; 1: mux_17145 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17146;
  function [0:0] mux_17146(input [0:0] sel);
    case (sel) 0: mux_17146 = 1'h0; 1: mux_17146 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_17147 = 1'h0;
  wire [0:0] v_17148;
  wire [0:0] v_17149;
  wire [0:0] act_17150;
  wire [0:0] v_17151;
  wire [0:0] v_17152;
  wire [0:0] v_17153;
  reg [0:0] v_17154 = 1'h0;
  wire [0:0] v_17155;
  wire [0:0] v_17156;
  wire [0:0] act_17157;
  wire [0:0] v_17158;
  wire [0:0] v_17159;
  wire [0:0] v_17160;
  reg [0:0] v_17161 = 1'h0;
  wire [0:0] v_17162;
  wire [0:0] v_17163;
  wire [0:0] act_17164;
  wire [0:0] v_17165;
  wire [0:0] v_17166;
  wire [0:0] v_17167;
  wire [0:0] vin0_consume_en_17168;
  wire [0:0] vout_canPeek_17168;
  wire [7:0] vout_peek_17168;
  wire [0:0] v_17169;
  wire [0:0] v_17170;
  function [0:0] mux_17170(input [0:0] sel);
    case (sel) 0: mux_17170 = 1'h0; 1: mux_17170 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17171;
  wire [0:0] v_17172;
  wire [0:0] v_17173;
  wire [0:0] v_17174;
  wire [0:0] v_17175;
  function [0:0] mux_17175(input [0:0] sel);
    case (sel) 0: mux_17175 = 1'h0; 1: mux_17175 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17176;
  wire [0:0] vin0_consume_en_17177;
  wire [0:0] vout_canPeek_17177;
  wire [7:0] vout_peek_17177;
  wire [0:0] v_17178;
  wire [0:0] v_17179;
  function [0:0] mux_17179(input [0:0] sel);
    case (sel) 0: mux_17179 = 1'h0; 1: mux_17179 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17180;
  function [0:0] mux_17180(input [0:0] sel);
    case (sel) 0: mux_17180 = 1'h0; 1: mux_17180 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17181;
  wire [0:0] v_17182;
  wire [0:0] v_17183;
  wire [0:0] v_17184;
  wire [0:0] v_17185;
  wire [0:0] v_17186;
  wire [0:0] v_17187;
  function [0:0] mux_17187(input [0:0] sel);
    case (sel) 0: mux_17187 = 1'h0; 1: mux_17187 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17188;
  wire [0:0] v_17189;
  wire [0:0] v_17190;
  wire [0:0] v_17191;
  wire [0:0] v_17192;
  function [0:0] mux_17192(input [0:0] sel);
    case (sel) 0: mux_17192 = 1'h0; 1: mux_17192 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17193;
  wire [0:0] v_17194;
  wire [0:0] v_17195;
  wire [0:0] v_17196;
  function [0:0] mux_17196(input [0:0] sel);
    case (sel) 0: mux_17196 = 1'h0; 1: mux_17196 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17197;
  function [0:0] mux_17197(input [0:0] sel);
    case (sel) 0: mux_17197 = 1'h0; 1: mux_17197 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_17198 = 1'h0;
  wire [0:0] v_17199;
  wire [0:0] v_17200;
  wire [0:0] act_17201;
  wire [0:0] v_17202;
  wire [0:0] v_17203;
  wire [0:0] v_17204;
  wire [0:0] vin0_consume_en_17205;
  wire [0:0] vout_canPeek_17205;
  wire [7:0] vout_peek_17205;
  wire [0:0] v_17206;
  wire [0:0] v_17207;
  function [0:0] mux_17207(input [0:0] sel);
    case (sel) 0: mux_17207 = 1'h0; 1: mux_17207 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17208;
  wire [0:0] v_17209;
  wire [0:0] v_17210;
  wire [0:0] v_17211;
  wire [0:0] v_17212;
  function [0:0] mux_17212(input [0:0] sel);
    case (sel) 0: mux_17212 = 1'h0; 1: mux_17212 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17213;
  wire [0:0] vin0_consume_en_17214;
  wire [0:0] vout_canPeek_17214;
  wire [7:0] vout_peek_17214;
  wire [0:0] v_17215;
  wire [0:0] v_17216;
  function [0:0] mux_17216(input [0:0] sel);
    case (sel) 0: mux_17216 = 1'h0; 1: mux_17216 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17217;
  function [0:0] mux_17217(input [0:0] sel);
    case (sel) 0: mux_17217 = 1'h0; 1: mux_17217 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17218;
  wire [0:0] v_17219;
  wire [0:0] v_17220;
  wire [0:0] v_17221;
  wire [0:0] v_17222;
  wire [0:0] v_17223;
  wire [0:0] v_17224;
  function [0:0] mux_17224(input [0:0] sel);
    case (sel) 0: mux_17224 = 1'h0; 1: mux_17224 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17225;
  function [0:0] mux_17225(input [0:0] sel);
    case (sel) 0: mux_17225 = 1'h0; 1: mux_17225 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17226;
  wire [0:0] v_17227;
  wire [0:0] v_17228;
  wire [0:0] v_17229;
  function [0:0] mux_17229(input [0:0] sel);
    case (sel) 0: mux_17229 = 1'h0; 1: mux_17229 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17230;
  function [0:0] mux_17230(input [0:0] sel);
    case (sel) 0: mux_17230 = 1'h0; 1: mux_17230 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17231;
  wire [0:0] v_17232;
  wire [0:0] v_17233;
  wire [0:0] v_17234;
  wire [0:0] v_17235;
  wire [0:0] v_17236;
  function [0:0] mux_17236(input [0:0] sel);
    case (sel) 0: mux_17236 = 1'h0; 1: mux_17236 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17237;
  wire [0:0] v_17238;
  wire [0:0] v_17239;
  wire [0:0] v_17240;
  wire [0:0] v_17241;
  function [0:0] mux_17241(input [0:0] sel);
    case (sel) 0: mux_17241 = 1'h0; 1: mux_17241 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17242;
  wire [0:0] v_17243;
  wire [0:0] v_17244;
  wire [0:0] v_17245;
  function [0:0] mux_17245(input [0:0] sel);
    case (sel) 0: mux_17245 = 1'h0; 1: mux_17245 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17246;
  function [0:0] mux_17246(input [0:0] sel);
    case (sel) 0: mux_17246 = 1'h0; 1: mux_17246 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_17247 = 1'h0;
  wire [0:0] v_17248;
  wire [0:0] v_17249;
  wire [0:0] act_17250;
  wire [0:0] v_17251;
  wire [0:0] v_17252;
  wire [0:0] v_17253;
  reg [0:0] v_17254 = 1'h0;
  wire [0:0] v_17255;
  wire [0:0] v_17256;
  wire [0:0] act_17257;
  wire [0:0] v_17258;
  wire [0:0] v_17259;
  wire [0:0] v_17260;
  wire [0:0] vin0_consume_en_17261;
  wire [0:0] vout_canPeek_17261;
  wire [7:0] vout_peek_17261;
  wire [0:0] v_17262;
  wire [0:0] v_17263;
  function [0:0] mux_17263(input [0:0] sel);
    case (sel) 0: mux_17263 = 1'h0; 1: mux_17263 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17264;
  wire [0:0] v_17265;
  wire [0:0] v_17266;
  wire [0:0] v_17267;
  wire [0:0] v_17268;
  function [0:0] mux_17268(input [0:0] sel);
    case (sel) 0: mux_17268 = 1'h0; 1: mux_17268 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17269;
  wire [0:0] vin0_consume_en_17270;
  wire [0:0] vout_canPeek_17270;
  wire [7:0] vout_peek_17270;
  wire [0:0] v_17271;
  wire [0:0] v_17272;
  function [0:0] mux_17272(input [0:0] sel);
    case (sel) 0: mux_17272 = 1'h0; 1: mux_17272 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17273;
  function [0:0] mux_17273(input [0:0] sel);
    case (sel) 0: mux_17273 = 1'h0; 1: mux_17273 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17274;
  wire [0:0] v_17275;
  wire [0:0] v_17276;
  wire [0:0] v_17277;
  wire [0:0] v_17278;
  wire [0:0] v_17279;
  wire [0:0] v_17280;
  function [0:0] mux_17280(input [0:0] sel);
    case (sel) 0: mux_17280 = 1'h0; 1: mux_17280 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17281;
  wire [0:0] v_17282;
  wire [0:0] v_17283;
  wire [0:0] v_17284;
  wire [0:0] v_17285;
  function [0:0] mux_17285(input [0:0] sel);
    case (sel) 0: mux_17285 = 1'h0; 1: mux_17285 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17286;
  wire [0:0] v_17287;
  wire [0:0] v_17288;
  wire [0:0] v_17289;
  function [0:0] mux_17289(input [0:0] sel);
    case (sel) 0: mux_17289 = 1'h0; 1: mux_17289 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17290;
  function [0:0] mux_17290(input [0:0] sel);
    case (sel) 0: mux_17290 = 1'h0; 1: mux_17290 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_17291 = 1'h0;
  wire [0:0] v_17292;
  wire [0:0] v_17293;
  wire [0:0] act_17294;
  wire [0:0] v_17295;
  wire [0:0] v_17296;
  wire [0:0] v_17297;
  wire [0:0] vin0_consume_en_17298;
  wire [0:0] vout_canPeek_17298;
  wire [7:0] vout_peek_17298;
  wire [0:0] v_17299;
  wire [0:0] v_17300;
  function [0:0] mux_17300(input [0:0] sel);
    case (sel) 0: mux_17300 = 1'h0; 1: mux_17300 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17301;
  wire [0:0] v_17302;
  wire [0:0] v_17303;
  wire [0:0] v_17304;
  wire [0:0] v_17305;
  function [0:0] mux_17305(input [0:0] sel);
    case (sel) 0: mux_17305 = 1'h0; 1: mux_17305 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17306;
  wire [0:0] vin0_consume_en_17307;
  wire [0:0] vout_canPeek_17307;
  wire [7:0] vout_peek_17307;
  wire [0:0] v_17308;
  wire [0:0] v_17309;
  function [0:0] mux_17309(input [0:0] sel);
    case (sel) 0: mux_17309 = 1'h0; 1: mux_17309 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17310;
  function [0:0] mux_17310(input [0:0] sel);
    case (sel) 0: mux_17310 = 1'h0; 1: mux_17310 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17311;
  wire [0:0] v_17312;
  wire [0:0] v_17313;
  wire [0:0] v_17314;
  wire [0:0] v_17315;
  wire [0:0] v_17316;
  wire [0:0] v_17317;
  function [0:0] mux_17317(input [0:0] sel);
    case (sel) 0: mux_17317 = 1'h0; 1: mux_17317 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17318;
  function [0:0] mux_17318(input [0:0] sel);
    case (sel) 0: mux_17318 = 1'h0; 1: mux_17318 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17319;
  wire [0:0] v_17320;
  wire [0:0] v_17321;
  wire [0:0] v_17322;
  function [0:0] mux_17322(input [0:0] sel);
    case (sel) 0: mux_17322 = 1'h0; 1: mux_17322 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17323;
  function [0:0] mux_17323(input [0:0] sel);
    case (sel) 0: mux_17323 = 1'h0; 1: mux_17323 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17324;
  wire [0:0] v_17325;
  wire [0:0] v_17326;
  wire [0:0] v_17327;
  wire [0:0] v_17328;
  wire [0:0] v_17329;
  function [0:0] mux_17329(input [0:0] sel);
    case (sel) 0: mux_17329 = 1'h0; 1: mux_17329 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17330;
  function [0:0] mux_17330(input [0:0] sel);
    case (sel) 0: mux_17330 = 1'h0; 1: mux_17330 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17331;
  wire [0:0] v_17332;
  wire [0:0] v_17333;
  wire [0:0] v_17334;
  function [0:0] mux_17334(input [0:0] sel);
    case (sel) 0: mux_17334 = 1'h0; 1: mux_17334 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17335;
  function [0:0] mux_17335(input [0:0] sel);
    case (sel) 0: mux_17335 = 1'h0; 1: mux_17335 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17336;
  wire [0:0] v_17337;
  wire [0:0] v_17338;
  wire [0:0] v_17339;
  wire [0:0] v_17340;
  wire [0:0] v_17341;
  function [0:0] mux_17341(input [0:0] sel);
    case (sel) 0: mux_17341 = 1'h0; 1: mux_17341 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17342;
  function [0:0] mux_17342(input [0:0] sel);
    case (sel) 0: mux_17342 = 1'h0; 1: mux_17342 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17343;
  wire [0:0] v_17344;
  wire [0:0] v_17345;
  wire [0:0] v_17346;
  function [0:0] mux_17346(input [0:0] sel);
    case (sel) 0: mux_17346 = 1'h0; 1: mux_17346 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17347;
  function [0:0] mux_17347(input [0:0] sel);
    case (sel) 0: mux_17347 = 1'h0; 1: mux_17347 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17348;
  wire [0:0] v_17349;
  wire [0:0] v_17350;
  wire [0:0] v_17351;
  wire [0:0] v_17352;
  wire [0:0] v_17353;
  function [0:0] mux_17353(input [0:0] sel);
    case (sel) 0: mux_17353 = 1'h0; 1: mux_17353 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17354;
  wire [0:0] v_17355;
  wire [0:0] v_17356;
  wire [0:0] v_17357;
  wire [0:0] v_17358;
  function [0:0] mux_17358(input [0:0] sel);
    case (sel) 0: mux_17358 = 1'h0; 1: mux_17358 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17359;
  wire [0:0] v_17360;
  wire [0:0] v_17361;
  wire [0:0] v_17362;
  function [0:0] mux_17362(input [0:0] sel);
    case (sel) 0: mux_17362 = 1'h0; 1: mux_17362 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17363;
  function [0:0] mux_17363(input [0:0] sel);
    case (sel) 0: mux_17363 = 1'h0; 1: mux_17363 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_17364 = 1'h0;
  wire [0:0] v_17365;
  wire [0:0] v_17366;
  wire [0:0] act_17367;
  wire [0:0] v_17368;
  wire [0:0] v_17369;
  wire [0:0] v_17370;
  reg [0:0] v_17371 = 1'h0;
  wire [0:0] v_17372;
  wire [0:0] v_17373;
  wire [0:0] act_17374;
  wire [0:0] v_17375;
  wire [0:0] v_17376;
  wire [0:0] v_17377;
  reg [0:0] v_17378 = 1'h0;
  wire [0:0] v_17379;
  wire [0:0] v_17380;
  wire [0:0] act_17381;
  wire [0:0] v_17382;
  wire [0:0] v_17383;
  wire [0:0] v_17384;
  reg [0:0] v_17385 = 1'h0;
  wire [0:0] v_17386;
  wire [0:0] v_17387;
  wire [0:0] act_17388;
  wire [0:0] v_17389;
  wire [0:0] v_17390;
  wire [0:0] v_17391;
  wire [0:0] vin0_consume_en_17392;
  wire [0:0] vout_canPeek_17392;
  wire [7:0] vout_peek_17392;
  wire [0:0] v_17393;
  wire [0:0] v_17394;
  function [0:0] mux_17394(input [0:0] sel);
    case (sel) 0: mux_17394 = 1'h0; 1: mux_17394 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17395;
  wire [0:0] v_17396;
  wire [0:0] v_17397;
  wire [0:0] v_17398;
  wire [0:0] v_17399;
  function [0:0] mux_17399(input [0:0] sel);
    case (sel) 0: mux_17399 = 1'h0; 1: mux_17399 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17400;
  wire [0:0] vin0_consume_en_17401;
  wire [0:0] vout_canPeek_17401;
  wire [7:0] vout_peek_17401;
  wire [0:0] v_17402;
  wire [0:0] v_17403;
  function [0:0] mux_17403(input [0:0] sel);
    case (sel) 0: mux_17403 = 1'h0; 1: mux_17403 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17404;
  function [0:0] mux_17404(input [0:0] sel);
    case (sel) 0: mux_17404 = 1'h0; 1: mux_17404 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17405;
  wire [0:0] v_17406;
  wire [0:0] v_17407;
  wire [0:0] v_17408;
  wire [0:0] v_17409;
  wire [0:0] v_17410;
  wire [0:0] v_17411;
  function [0:0] mux_17411(input [0:0] sel);
    case (sel) 0: mux_17411 = 1'h0; 1: mux_17411 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17412;
  wire [0:0] v_17413;
  wire [0:0] v_17414;
  wire [0:0] v_17415;
  wire [0:0] v_17416;
  function [0:0] mux_17416(input [0:0] sel);
    case (sel) 0: mux_17416 = 1'h0; 1: mux_17416 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17417;
  wire [0:0] v_17418;
  wire [0:0] v_17419;
  wire [0:0] v_17420;
  function [0:0] mux_17420(input [0:0] sel);
    case (sel) 0: mux_17420 = 1'h0; 1: mux_17420 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17421;
  function [0:0] mux_17421(input [0:0] sel);
    case (sel) 0: mux_17421 = 1'h0; 1: mux_17421 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_17422 = 1'h0;
  wire [0:0] v_17423;
  wire [0:0] v_17424;
  wire [0:0] act_17425;
  wire [0:0] v_17426;
  wire [0:0] v_17427;
  wire [0:0] v_17428;
  wire [0:0] vin0_consume_en_17429;
  wire [0:0] vout_canPeek_17429;
  wire [7:0] vout_peek_17429;
  wire [0:0] v_17430;
  wire [0:0] v_17431;
  function [0:0] mux_17431(input [0:0] sel);
    case (sel) 0: mux_17431 = 1'h0; 1: mux_17431 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17432;
  wire [0:0] v_17433;
  wire [0:0] v_17434;
  wire [0:0] v_17435;
  wire [0:0] v_17436;
  function [0:0] mux_17436(input [0:0] sel);
    case (sel) 0: mux_17436 = 1'h0; 1: mux_17436 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17437;
  wire [0:0] vin0_consume_en_17438;
  wire [0:0] vout_canPeek_17438;
  wire [7:0] vout_peek_17438;
  wire [0:0] v_17439;
  wire [0:0] v_17440;
  function [0:0] mux_17440(input [0:0] sel);
    case (sel) 0: mux_17440 = 1'h0; 1: mux_17440 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17441;
  function [0:0] mux_17441(input [0:0] sel);
    case (sel) 0: mux_17441 = 1'h0; 1: mux_17441 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17442;
  wire [0:0] v_17443;
  wire [0:0] v_17444;
  wire [0:0] v_17445;
  wire [0:0] v_17446;
  wire [0:0] v_17447;
  wire [0:0] v_17448;
  function [0:0] mux_17448(input [0:0] sel);
    case (sel) 0: mux_17448 = 1'h0; 1: mux_17448 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17449;
  function [0:0] mux_17449(input [0:0] sel);
    case (sel) 0: mux_17449 = 1'h0; 1: mux_17449 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17450;
  wire [0:0] v_17451;
  wire [0:0] v_17452;
  wire [0:0] v_17453;
  function [0:0] mux_17453(input [0:0] sel);
    case (sel) 0: mux_17453 = 1'h0; 1: mux_17453 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17454;
  function [0:0] mux_17454(input [0:0] sel);
    case (sel) 0: mux_17454 = 1'h0; 1: mux_17454 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17455;
  wire [0:0] v_17456;
  wire [0:0] v_17457;
  wire [0:0] v_17458;
  wire [0:0] v_17459;
  wire [0:0] v_17460;
  function [0:0] mux_17460(input [0:0] sel);
    case (sel) 0: mux_17460 = 1'h0; 1: mux_17460 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17461;
  wire [0:0] v_17462;
  wire [0:0] v_17463;
  wire [0:0] v_17464;
  wire [0:0] v_17465;
  function [0:0] mux_17465(input [0:0] sel);
    case (sel) 0: mux_17465 = 1'h0; 1: mux_17465 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17466;
  wire [0:0] v_17467;
  wire [0:0] v_17468;
  wire [0:0] v_17469;
  function [0:0] mux_17469(input [0:0] sel);
    case (sel) 0: mux_17469 = 1'h0; 1: mux_17469 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17470;
  function [0:0] mux_17470(input [0:0] sel);
    case (sel) 0: mux_17470 = 1'h0; 1: mux_17470 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_17471 = 1'h0;
  wire [0:0] v_17472;
  wire [0:0] v_17473;
  wire [0:0] act_17474;
  wire [0:0] v_17475;
  wire [0:0] v_17476;
  wire [0:0] v_17477;
  reg [0:0] v_17478 = 1'h0;
  wire [0:0] v_17479;
  wire [0:0] v_17480;
  wire [0:0] act_17481;
  wire [0:0] v_17482;
  wire [0:0] v_17483;
  wire [0:0] v_17484;
  wire [0:0] vin0_consume_en_17485;
  wire [0:0] vout_canPeek_17485;
  wire [7:0] vout_peek_17485;
  wire [0:0] v_17486;
  wire [0:0] v_17487;
  function [0:0] mux_17487(input [0:0] sel);
    case (sel) 0: mux_17487 = 1'h0; 1: mux_17487 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17488;
  wire [0:0] v_17489;
  wire [0:0] v_17490;
  wire [0:0] v_17491;
  wire [0:0] v_17492;
  function [0:0] mux_17492(input [0:0] sel);
    case (sel) 0: mux_17492 = 1'h0; 1: mux_17492 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17493;
  wire [0:0] vin0_consume_en_17494;
  wire [0:0] vout_canPeek_17494;
  wire [7:0] vout_peek_17494;
  wire [0:0] v_17495;
  wire [0:0] v_17496;
  function [0:0] mux_17496(input [0:0] sel);
    case (sel) 0: mux_17496 = 1'h0; 1: mux_17496 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17497;
  function [0:0] mux_17497(input [0:0] sel);
    case (sel) 0: mux_17497 = 1'h0; 1: mux_17497 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17498;
  wire [0:0] v_17499;
  wire [0:0] v_17500;
  wire [0:0] v_17501;
  wire [0:0] v_17502;
  wire [0:0] v_17503;
  wire [0:0] v_17504;
  function [0:0] mux_17504(input [0:0] sel);
    case (sel) 0: mux_17504 = 1'h0; 1: mux_17504 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17505;
  wire [0:0] v_17506;
  wire [0:0] v_17507;
  wire [0:0] v_17508;
  wire [0:0] v_17509;
  function [0:0] mux_17509(input [0:0] sel);
    case (sel) 0: mux_17509 = 1'h0; 1: mux_17509 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17510;
  wire [0:0] v_17511;
  wire [0:0] v_17512;
  wire [0:0] v_17513;
  function [0:0] mux_17513(input [0:0] sel);
    case (sel) 0: mux_17513 = 1'h0; 1: mux_17513 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17514;
  function [0:0] mux_17514(input [0:0] sel);
    case (sel) 0: mux_17514 = 1'h0; 1: mux_17514 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_17515 = 1'h0;
  wire [0:0] v_17516;
  wire [0:0] v_17517;
  wire [0:0] act_17518;
  wire [0:0] v_17519;
  wire [0:0] v_17520;
  wire [0:0] v_17521;
  wire [0:0] vin0_consume_en_17522;
  wire [0:0] vout_canPeek_17522;
  wire [7:0] vout_peek_17522;
  wire [0:0] v_17523;
  wire [0:0] v_17524;
  function [0:0] mux_17524(input [0:0] sel);
    case (sel) 0: mux_17524 = 1'h0; 1: mux_17524 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17525;
  wire [0:0] v_17526;
  wire [0:0] v_17527;
  wire [0:0] v_17528;
  wire [0:0] v_17529;
  function [0:0] mux_17529(input [0:0] sel);
    case (sel) 0: mux_17529 = 1'h0; 1: mux_17529 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17530;
  wire [0:0] vin0_consume_en_17531;
  wire [0:0] vout_canPeek_17531;
  wire [7:0] vout_peek_17531;
  wire [0:0] v_17532;
  wire [0:0] v_17533;
  function [0:0] mux_17533(input [0:0] sel);
    case (sel) 0: mux_17533 = 1'h0; 1: mux_17533 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17534;
  function [0:0] mux_17534(input [0:0] sel);
    case (sel) 0: mux_17534 = 1'h0; 1: mux_17534 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17535;
  wire [0:0] v_17536;
  wire [0:0] v_17537;
  wire [0:0] v_17538;
  wire [0:0] v_17539;
  wire [0:0] v_17540;
  wire [0:0] v_17541;
  function [0:0] mux_17541(input [0:0] sel);
    case (sel) 0: mux_17541 = 1'h0; 1: mux_17541 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17542;
  function [0:0] mux_17542(input [0:0] sel);
    case (sel) 0: mux_17542 = 1'h0; 1: mux_17542 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17543;
  wire [0:0] v_17544;
  wire [0:0] v_17545;
  wire [0:0] v_17546;
  function [0:0] mux_17546(input [0:0] sel);
    case (sel) 0: mux_17546 = 1'h0; 1: mux_17546 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17547;
  function [0:0] mux_17547(input [0:0] sel);
    case (sel) 0: mux_17547 = 1'h0; 1: mux_17547 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17548;
  wire [0:0] v_17549;
  wire [0:0] v_17550;
  wire [0:0] v_17551;
  wire [0:0] v_17552;
  wire [0:0] v_17553;
  function [0:0] mux_17553(input [0:0] sel);
    case (sel) 0: mux_17553 = 1'h0; 1: mux_17553 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17554;
  function [0:0] mux_17554(input [0:0] sel);
    case (sel) 0: mux_17554 = 1'h0; 1: mux_17554 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17555;
  wire [0:0] v_17556;
  wire [0:0] v_17557;
  wire [0:0] v_17558;
  function [0:0] mux_17558(input [0:0] sel);
    case (sel) 0: mux_17558 = 1'h0; 1: mux_17558 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17559;
  function [0:0] mux_17559(input [0:0] sel);
    case (sel) 0: mux_17559 = 1'h0; 1: mux_17559 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17560;
  wire [0:0] v_17561;
  wire [0:0] v_17562;
  wire [0:0] v_17563;
  wire [0:0] v_17564;
  wire [0:0] v_17565;
  function [0:0] mux_17565(input [0:0] sel);
    case (sel) 0: mux_17565 = 1'h0; 1: mux_17565 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17566;
  wire [0:0] v_17567;
  wire [0:0] v_17568;
  wire [0:0] v_17569;
  wire [0:0] v_17570;
  function [0:0] mux_17570(input [0:0] sel);
    case (sel) 0: mux_17570 = 1'h0; 1: mux_17570 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17571;
  wire [0:0] v_17572;
  wire [0:0] v_17573;
  wire [0:0] v_17574;
  function [0:0] mux_17574(input [0:0] sel);
    case (sel) 0: mux_17574 = 1'h0; 1: mux_17574 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17575;
  function [0:0] mux_17575(input [0:0] sel);
    case (sel) 0: mux_17575 = 1'h0; 1: mux_17575 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_17576 = 1'h0;
  wire [0:0] v_17577;
  wire [0:0] v_17578;
  wire [0:0] act_17579;
  wire [0:0] v_17580;
  wire [0:0] v_17581;
  wire [0:0] v_17582;
  reg [0:0] v_17583 = 1'h0;
  wire [0:0] v_17584;
  wire [0:0] v_17585;
  wire [0:0] act_17586;
  wire [0:0] v_17587;
  wire [0:0] v_17588;
  wire [0:0] v_17589;
  reg [0:0] v_17590 = 1'h0;
  wire [0:0] v_17591;
  wire [0:0] v_17592;
  wire [0:0] act_17593;
  wire [0:0] v_17594;
  wire [0:0] v_17595;
  wire [0:0] v_17596;
  wire [0:0] vin0_consume_en_17597;
  wire [0:0] vout_canPeek_17597;
  wire [7:0] vout_peek_17597;
  wire [0:0] v_17598;
  wire [0:0] v_17599;
  function [0:0] mux_17599(input [0:0] sel);
    case (sel) 0: mux_17599 = 1'h0; 1: mux_17599 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17600;
  wire [0:0] v_17601;
  wire [0:0] v_17602;
  wire [0:0] v_17603;
  wire [0:0] v_17604;
  function [0:0] mux_17604(input [0:0] sel);
    case (sel) 0: mux_17604 = 1'h0; 1: mux_17604 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17605;
  wire [0:0] vin0_consume_en_17606;
  wire [0:0] vout_canPeek_17606;
  wire [7:0] vout_peek_17606;
  wire [0:0] v_17607;
  wire [0:0] v_17608;
  function [0:0] mux_17608(input [0:0] sel);
    case (sel) 0: mux_17608 = 1'h0; 1: mux_17608 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17609;
  function [0:0] mux_17609(input [0:0] sel);
    case (sel) 0: mux_17609 = 1'h0; 1: mux_17609 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17610;
  wire [0:0] v_17611;
  wire [0:0] v_17612;
  wire [0:0] v_17613;
  wire [0:0] v_17614;
  wire [0:0] v_17615;
  wire [0:0] v_17616;
  function [0:0] mux_17616(input [0:0] sel);
    case (sel) 0: mux_17616 = 1'h0; 1: mux_17616 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17617;
  wire [0:0] v_17618;
  wire [0:0] v_17619;
  wire [0:0] v_17620;
  wire [0:0] v_17621;
  function [0:0] mux_17621(input [0:0] sel);
    case (sel) 0: mux_17621 = 1'h0; 1: mux_17621 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17622;
  wire [0:0] v_17623;
  wire [0:0] v_17624;
  wire [0:0] v_17625;
  function [0:0] mux_17625(input [0:0] sel);
    case (sel) 0: mux_17625 = 1'h0; 1: mux_17625 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17626;
  function [0:0] mux_17626(input [0:0] sel);
    case (sel) 0: mux_17626 = 1'h0; 1: mux_17626 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_17627 = 1'h0;
  wire [0:0] v_17628;
  wire [0:0] v_17629;
  wire [0:0] act_17630;
  wire [0:0] v_17631;
  wire [0:0] v_17632;
  wire [0:0] v_17633;
  wire [0:0] vin0_consume_en_17634;
  wire [0:0] vout_canPeek_17634;
  wire [7:0] vout_peek_17634;
  wire [0:0] v_17635;
  wire [0:0] v_17636;
  function [0:0] mux_17636(input [0:0] sel);
    case (sel) 0: mux_17636 = 1'h0; 1: mux_17636 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17637;
  wire [0:0] v_17638;
  wire [0:0] v_17639;
  wire [0:0] v_17640;
  wire [0:0] v_17641;
  function [0:0] mux_17641(input [0:0] sel);
    case (sel) 0: mux_17641 = 1'h0; 1: mux_17641 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17642;
  wire [0:0] vin0_consume_en_17643;
  wire [0:0] vout_canPeek_17643;
  wire [7:0] vout_peek_17643;
  wire [0:0] v_17644;
  wire [0:0] v_17645;
  function [0:0] mux_17645(input [0:0] sel);
    case (sel) 0: mux_17645 = 1'h0; 1: mux_17645 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17646;
  function [0:0] mux_17646(input [0:0] sel);
    case (sel) 0: mux_17646 = 1'h0; 1: mux_17646 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17647;
  wire [0:0] v_17648;
  wire [0:0] v_17649;
  wire [0:0] v_17650;
  wire [0:0] v_17651;
  wire [0:0] v_17652;
  wire [0:0] v_17653;
  function [0:0] mux_17653(input [0:0] sel);
    case (sel) 0: mux_17653 = 1'h0; 1: mux_17653 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17654;
  function [0:0] mux_17654(input [0:0] sel);
    case (sel) 0: mux_17654 = 1'h0; 1: mux_17654 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17655;
  wire [0:0] v_17656;
  wire [0:0] v_17657;
  wire [0:0] v_17658;
  function [0:0] mux_17658(input [0:0] sel);
    case (sel) 0: mux_17658 = 1'h0; 1: mux_17658 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17659;
  function [0:0] mux_17659(input [0:0] sel);
    case (sel) 0: mux_17659 = 1'h0; 1: mux_17659 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17660;
  wire [0:0] v_17661;
  wire [0:0] v_17662;
  wire [0:0] v_17663;
  wire [0:0] v_17664;
  wire [0:0] v_17665;
  function [0:0] mux_17665(input [0:0] sel);
    case (sel) 0: mux_17665 = 1'h0; 1: mux_17665 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17666;
  wire [0:0] v_17667;
  wire [0:0] v_17668;
  wire [0:0] v_17669;
  wire [0:0] v_17670;
  function [0:0] mux_17670(input [0:0] sel);
    case (sel) 0: mux_17670 = 1'h0; 1: mux_17670 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17671;
  wire [0:0] v_17672;
  wire [0:0] v_17673;
  wire [0:0] v_17674;
  function [0:0] mux_17674(input [0:0] sel);
    case (sel) 0: mux_17674 = 1'h0; 1: mux_17674 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17675;
  function [0:0] mux_17675(input [0:0] sel);
    case (sel) 0: mux_17675 = 1'h0; 1: mux_17675 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_17676 = 1'h0;
  wire [0:0] v_17677;
  wire [0:0] v_17678;
  wire [0:0] act_17679;
  wire [0:0] v_17680;
  wire [0:0] v_17681;
  wire [0:0] v_17682;
  reg [0:0] v_17683 = 1'h0;
  wire [0:0] v_17684;
  wire [0:0] v_17685;
  wire [0:0] act_17686;
  wire [0:0] v_17687;
  wire [0:0] v_17688;
  wire [0:0] v_17689;
  wire [0:0] vin0_consume_en_17690;
  wire [0:0] vout_canPeek_17690;
  wire [7:0] vout_peek_17690;
  wire [0:0] v_17691;
  wire [0:0] v_17692;
  function [0:0] mux_17692(input [0:0] sel);
    case (sel) 0: mux_17692 = 1'h0; 1: mux_17692 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17693;
  wire [0:0] v_17694;
  wire [0:0] v_17695;
  wire [0:0] v_17696;
  wire [0:0] v_17697;
  function [0:0] mux_17697(input [0:0] sel);
    case (sel) 0: mux_17697 = 1'h0; 1: mux_17697 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17698;
  wire [0:0] vin0_consume_en_17699;
  wire [0:0] vout_canPeek_17699;
  wire [7:0] vout_peek_17699;
  wire [0:0] v_17700;
  wire [0:0] v_17701;
  function [0:0] mux_17701(input [0:0] sel);
    case (sel) 0: mux_17701 = 1'h0; 1: mux_17701 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17702;
  function [0:0] mux_17702(input [0:0] sel);
    case (sel) 0: mux_17702 = 1'h0; 1: mux_17702 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17703;
  wire [0:0] v_17704;
  wire [0:0] v_17705;
  wire [0:0] v_17706;
  wire [0:0] v_17707;
  wire [0:0] v_17708;
  wire [0:0] v_17709;
  function [0:0] mux_17709(input [0:0] sel);
    case (sel) 0: mux_17709 = 1'h0; 1: mux_17709 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17710;
  wire [0:0] v_17711;
  wire [0:0] v_17712;
  wire [0:0] v_17713;
  wire [0:0] v_17714;
  function [0:0] mux_17714(input [0:0] sel);
    case (sel) 0: mux_17714 = 1'h0; 1: mux_17714 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17715;
  wire [0:0] v_17716;
  wire [0:0] v_17717;
  wire [0:0] v_17718;
  function [0:0] mux_17718(input [0:0] sel);
    case (sel) 0: mux_17718 = 1'h0; 1: mux_17718 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17719;
  function [0:0] mux_17719(input [0:0] sel);
    case (sel) 0: mux_17719 = 1'h0; 1: mux_17719 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_17720 = 1'h0;
  wire [0:0] v_17721;
  wire [0:0] v_17722;
  wire [0:0] act_17723;
  wire [0:0] v_17724;
  wire [0:0] v_17725;
  wire [0:0] v_17726;
  wire [0:0] vin0_consume_en_17727;
  wire [0:0] vout_canPeek_17727;
  wire [7:0] vout_peek_17727;
  wire [0:0] v_17728;
  wire [0:0] v_17729;
  function [0:0] mux_17729(input [0:0] sel);
    case (sel) 0: mux_17729 = 1'h0; 1: mux_17729 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17730;
  wire [0:0] v_17731;
  wire [0:0] v_17732;
  wire [0:0] v_17733;
  wire [0:0] v_17734;
  function [0:0] mux_17734(input [0:0] sel);
    case (sel) 0: mux_17734 = 1'h0; 1: mux_17734 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17735;
  wire [0:0] vin0_consume_en_17736;
  wire [0:0] vout_canPeek_17736;
  wire [7:0] vout_peek_17736;
  wire [0:0] v_17737;
  wire [0:0] v_17738;
  function [0:0] mux_17738(input [0:0] sel);
    case (sel) 0: mux_17738 = 1'h0; 1: mux_17738 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17739;
  function [0:0] mux_17739(input [0:0] sel);
    case (sel) 0: mux_17739 = 1'h0; 1: mux_17739 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17740;
  wire [0:0] v_17741;
  wire [0:0] v_17742;
  wire [0:0] v_17743;
  wire [0:0] v_17744;
  wire [0:0] v_17745;
  wire [0:0] v_17746;
  function [0:0] mux_17746(input [0:0] sel);
    case (sel) 0: mux_17746 = 1'h0; 1: mux_17746 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17747;
  function [0:0] mux_17747(input [0:0] sel);
    case (sel) 0: mux_17747 = 1'h0; 1: mux_17747 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17748;
  wire [0:0] v_17749;
  wire [0:0] v_17750;
  wire [0:0] v_17751;
  function [0:0] mux_17751(input [0:0] sel);
    case (sel) 0: mux_17751 = 1'h0; 1: mux_17751 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17752;
  function [0:0] mux_17752(input [0:0] sel);
    case (sel) 0: mux_17752 = 1'h0; 1: mux_17752 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17753;
  wire [0:0] v_17754;
  wire [0:0] v_17755;
  wire [0:0] v_17756;
  wire [0:0] v_17757;
  wire [0:0] v_17758;
  function [0:0] mux_17758(input [0:0] sel);
    case (sel) 0: mux_17758 = 1'h0; 1: mux_17758 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17759;
  function [0:0] mux_17759(input [0:0] sel);
    case (sel) 0: mux_17759 = 1'h0; 1: mux_17759 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17760;
  wire [0:0] v_17761;
  wire [0:0] v_17762;
  wire [0:0] v_17763;
  function [0:0] mux_17763(input [0:0] sel);
    case (sel) 0: mux_17763 = 1'h0; 1: mux_17763 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17764;
  function [0:0] mux_17764(input [0:0] sel);
    case (sel) 0: mux_17764 = 1'h0; 1: mux_17764 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17765;
  wire [0:0] v_17766;
  wire [0:0] v_17767;
  wire [0:0] v_17768;
  wire [0:0] v_17769;
  wire [0:0] v_17770;
  function [0:0] mux_17770(input [0:0] sel);
    case (sel) 0: mux_17770 = 1'h0; 1: mux_17770 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17771;
  function [0:0] mux_17771(input [0:0] sel);
    case (sel) 0: mux_17771 = 1'h0; 1: mux_17771 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17772;
  wire [0:0] v_17773;
  wire [0:0] v_17774;
  wire [0:0] v_17775;
  function [0:0] mux_17775(input [0:0] sel);
    case (sel) 0: mux_17775 = 1'h0; 1: mux_17775 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17776;
  function [0:0] mux_17776(input [0:0] sel);
    case (sel) 0: mux_17776 = 1'h0; 1: mux_17776 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17777;
  wire [0:0] v_17778;
  wire [0:0] v_17779;
  wire [0:0] v_17780;
  wire [0:0] v_17781;
  wire [0:0] v_17782;
  function [0:0] mux_17782(input [0:0] sel);
    case (sel) 0: mux_17782 = 1'h0; 1: mux_17782 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17783;
  function [0:0] mux_17783(input [0:0] sel);
    case (sel) 0: mux_17783 = 1'h0; 1: mux_17783 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17784;
  wire [0:0] v_17785;
  wire [0:0] v_17786;
  wire [0:0] v_17787;
  function [0:0] mux_17787(input [0:0] sel);
    case (sel) 0: mux_17787 = 1'h0; 1: mux_17787 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17788;
  function [0:0] mux_17788(input [0:0] sel);
    case (sel) 0: mux_17788 = 1'h0; 1: mux_17788 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17789;
  wire [0:0] v_17790;
  wire [0:0] v_17791;
  wire [0:0] v_17792;
  wire [0:0] v_17793;
  wire [0:0] v_17794;
  function [0:0] mux_17794(input [0:0] sel);
    case (sel) 0: mux_17794 = 1'h0; 1: mux_17794 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17795;
  wire [0:0] v_17796;
  wire [0:0] v_17797;
  wire [0:0] v_17798;
  wire [0:0] v_17799;
  function [0:0] mux_17799(input [0:0] sel);
    case (sel) 0: mux_17799 = 1'h0; 1: mux_17799 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17800;
  wire [0:0] v_17801;
  wire [0:0] v_17802;
  wire [0:0] v_17803;
  function [0:0] mux_17803(input [0:0] sel);
    case (sel) 0: mux_17803 = 1'h0; 1: mux_17803 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17804;
  function [0:0] mux_17804(input [0:0] sel);
    case (sel) 0: mux_17804 = 1'h0; 1: mux_17804 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_17805 = 1'h0;
  wire [0:0] v_17806;
  wire [0:0] v_17807;
  wire [0:0] act_17808;
  wire [0:0] v_17809;
  wire [0:0] v_17810;
  wire [0:0] v_17811;
  reg [0:0] v_17812 = 1'h0;
  wire [0:0] v_17813;
  wire [0:0] v_17814;
  wire [0:0] act_17815;
  wire [0:0] v_17816;
  wire [0:0] v_17817;
  wire [0:0] v_17818;
  reg [0:0] v_17819 = 1'h0;
  wire [0:0] v_17820;
  wire [0:0] v_17821;
  wire [0:0] act_17822;
  wire [0:0] v_17823;
  wire [0:0] v_17824;
  wire [0:0] v_17825;
  reg [0:0] v_17826 = 1'h0;
  wire [0:0] v_17827;
  wire [0:0] v_17828;
  wire [0:0] act_17829;
  wire [0:0] v_17830;
  wire [0:0] v_17831;
  wire [0:0] v_17832;
  reg [0:0] v_17833 = 1'h0;
  wire [0:0] v_17834;
  wire [0:0] v_17835;
  wire [0:0] act_17836;
  wire [0:0] v_17837;
  wire [0:0] v_17838;
  wire [0:0] v_17839;
  wire [0:0] vin0_consume_en_17840;
  wire [0:0] vout_canPeek_17840;
  wire [7:0] vout_peek_17840;
  wire [0:0] v_17841;
  wire [0:0] v_17842;
  function [0:0] mux_17842(input [0:0] sel);
    case (sel) 0: mux_17842 = 1'h0; 1: mux_17842 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17843;
  wire [0:0] v_17844;
  wire [0:0] v_17845;
  wire [0:0] v_17846;
  wire [0:0] v_17847;
  function [0:0] mux_17847(input [0:0] sel);
    case (sel) 0: mux_17847 = 1'h0; 1: mux_17847 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17848;
  wire [0:0] vin0_consume_en_17849;
  wire [0:0] vout_canPeek_17849;
  wire [7:0] vout_peek_17849;
  wire [0:0] v_17850;
  wire [0:0] v_17851;
  function [0:0] mux_17851(input [0:0] sel);
    case (sel) 0: mux_17851 = 1'h0; 1: mux_17851 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17852;
  function [0:0] mux_17852(input [0:0] sel);
    case (sel) 0: mux_17852 = 1'h0; 1: mux_17852 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17853;
  wire [0:0] v_17854;
  wire [0:0] v_17855;
  wire [0:0] v_17856;
  wire [0:0] v_17857;
  wire [0:0] v_17858;
  wire [0:0] v_17859;
  function [0:0] mux_17859(input [0:0] sel);
    case (sel) 0: mux_17859 = 1'h0; 1: mux_17859 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17860;
  wire [0:0] v_17861;
  wire [0:0] v_17862;
  wire [0:0] v_17863;
  wire [0:0] v_17864;
  function [0:0] mux_17864(input [0:0] sel);
    case (sel) 0: mux_17864 = 1'h0; 1: mux_17864 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17865;
  wire [0:0] v_17866;
  wire [0:0] v_17867;
  wire [0:0] v_17868;
  function [0:0] mux_17868(input [0:0] sel);
    case (sel) 0: mux_17868 = 1'h0; 1: mux_17868 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17869;
  function [0:0] mux_17869(input [0:0] sel);
    case (sel) 0: mux_17869 = 1'h0; 1: mux_17869 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_17870 = 1'h0;
  wire [0:0] v_17871;
  wire [0:0] v_17872;
  wire [0:0] act_17873;
  wire [0:0] v_17874;
  wire [0:0] v_17875;
  wire [0:0] v_17876;
  wire [0:0] vin0_consume_en_17877;
  wire [0:0] vout_canPeek_17877;
  wire [7:0] vout_peek_17877;
  wire [0:0] v_17878;
  wire [0:0] v_17879;
  function [0:0] mux_17879(input [0:0] sel);
    case (sel) 0: mux_17879 = 1'h0; 1: mux_17879 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17880;
  wire [0:0] v_17881;
  wire [0:0] v_17882;
  wire [0:0] v_17883;
  wire [0:0] v_17884;
  function [0:0] mux_17884(input [0:0] sel);
    case (sel) 0: mux_17884 = 1'h0; 1: mux_17884 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17885;
  wire [0:0] vin0_consume_en_17886;
  wire [0:0] vout_canPeek_17886;
  wire [7:0] vout_peek_17886;
  wire [0:0] v_17887;
  wire [0:0] v_17888;
  function [0:0] mux_17888(input [0:0] sel);
    case (sel) 0: mux_17888 = 1'h0; 1: mux_17888 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17889;
  function [0:0] mux_17889(input [0:0] sel);
    case (sel) 0: mux_17889 = 1'h0; 1: mux_17889 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17890;
  wire [0:0] v_17891;
  wire [0:0] v_17892;
  wire [0:0] v_17893;
  wire [0:0] v_17894;
  wire [0:0] v_17895;
  wire [0:0] v_17896;
  function [0:0] mux_17896(input [0:0] sel);
    case (sel) 0: mux_17896 = 1'h0; 1: mux_17896 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17897;
  function [0:0] mux_17897(input [0:0] sel);
    case (sel) 0: mux_17897 = 1'h0; 1: mux_17897 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17898;
  wire [0:0] v_17899;
  wire [0:0] v_17900;
  wire [0:0] v_17901;
  function [0:0] mux_17901(input [0:0] sel);
    case (sel) 0: mux_17901 = 1'h0; 1: mux_17901 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17902;
  function [0:0] mux_17902(input [0:0] sel);
    case (sel) 0: mux_17902 = 1'h0; 1: mux_17902 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17903;
  wire [0:0] v_17904;
  wire [0:0] v_17905;
  wire [0:0] v_17906;
  wire [0:0] v_17907;
  wire [0:0] v_17908;
  function [0:0] mux_17908(input [0:0] sel);
    case (sel) 0: mux_17908 = 1'h0; 1: mux_17908 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17909;
  wire [0:0] v_17910;
  wire [0:0] v_17911;
  wire [0:0] v_17912;
  wire [0:0] v_17913;
  function [0:0] mux_17913(input [0:0] sel);
    case (sel) 0: mux_17913 = 1'h0; 1: mux_17913 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17914;
  wire [0:0] v_17915;
  wire [0:0] v_17916;
  wire [0:0] v_17917;
  function [0:0] mux_17917(input [0:0] sel);
    case (sel) 0: mux_17917 = 1'h0; 1: mux_17917 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17918;
  function [0:0] mux_17918(input [0:0] sel);
    case (sel) 0: mux_17918 = 1'h0; 1: mux_17918 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_17919 = 1'h0;
  wire [0:0] v_17920;
  wire [0:0] v_17921;
  wire [0:0] act_17922;
  wire [0:0] v_17923;
  wire [0:0] v_17924;
  wire [0:0] v_17925;
  reg [0:0] v_17926 = 1'h0;
  wire [0:0] v_17927;
  wire [0:0] v_17928;
  wire [0:0] act_17929;
  wire [0:0] v_17930;
  wire [0:0] v_17931;
  wire [0:0] v_17932;
  wire [0:0] vin0_consume_en_17933;
  wire [0:0] vout_canPeek_17933;
  wire [7:0] vout_peek_17933;
  wire [0:0] v_17934;
  wire [0:0] v_17935;
  function [0:0] mux_17935(input [0:0] sel);
    case (sel) 0: mux_17935 = 1'h0; 1: mux_17935 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17936;
  wire [0:0] v_17937;
  wire [0:0] v_17938;
  wire [0:0] v_17939;
  wire [0:0] v_17940;
  function [0:0] mux_17940(input [0:0] sel);
    case (sel) 0: mux_17940 = 1'h0; 1: mux_17940 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17941;
  wire [0:0] vin0_consume_en_17942;
  wire [0:0] vout_canPeek_17942;
  wire [7:0] vout_peek_17942;
  wire [0:0] v_17943;
  wire [0:0] v_17944;
  function [0:0] mux_17944(input [0:0] sel);
    case (sel) 0: mux_17944 = 1'h0; 1: mux_17944 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17945;
  function [0:0] mux_17945(input [0:0] sel);
    case (sel) 0: mux_17945 = 1'h0; 1: mux_17945 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17946;
  wire [0:0] v_17947;
  wire [0:0] v_17948;
  wire [0:0] v_17949;
  wire [0:0] v_17950;
  wire [0:0] v_17951;
  wire [0:0] v_17952;
  function [0:0] mux_17952(input [0:0] sel);
    case (sel) 0: mux_17952 = 1'h0; 1: mux_17952 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17953;
  wire [0:0] v_17954;
  wire [0:0] v_17955;
  wire [0:0] v_17956;
  wire [0:0] v_17957;
  function [0:0] mux_17957(input [0:0] sel);
    case (sel) 0: mux_17957 = 1'h0; 1: mux_17957 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17958;
  wire [0:0] v_17959;
  wire [0:0] v_17960;
  wire [0:0] v_17961;
  function [0:0] mux_17961(input [0:0] sel);
    case (sel) 0: mux_17961 = 1'h0; 1: mux_17961 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17962;
  function [0:0] mux_17962(input [0:0] sel);
    case (sel) 0: mux_17962 = 1'h0; 1: mux_17962 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_17963 = 1'h0;
  wire [0:0] v_17964;
  wire [0:0] v_17965;
  wire [0:0] act_17966;
  wire [0:0] v_17967;
  wire [0:0] v_17968;
  wire [0:0] v_17969;
  wire [0:0] vin0_consume_en_17970;
  wire [0:0] vout_canPeek_17970;
  wire [7:0] vout_peek_17970;
  wire [0:0] v_17971;
  wire [0:0] v_17972;
  function [0:0] mux_17972(input [0:0] sel);
    case (sel) 0: mux_17972 = 1'h0; 1: mux_17972 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17973;
  wire [0:0] v_17974;
  wire [0:0] v_17975;
  wire [0:0] v_17976;
  wire [0:0] v_17977;
  function [0:0] mux_17977(input [0:0] sel);
    case (sel) 0: mux_17977 = 1'h0; 1: mux_17977 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17978;
  wire [0:0] vin0_consume_en_17979;
  wire [0:0] vout_canPeek_17979;
  wire [7:0] vout_peek_17979;
  wire [0:0] v_17980;
  wire [0:0] v_17981;
  function [0:0] mux_17981(input [0:0] sel);
    case (sel) 0: mux_17981 = 1'h0; 1: mux_17981 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17982;
  function [0:0] mux_17982(input [0:0] sel);
    case (sel) 0: mux_17982 = 1'h0; 1: mux_17982 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17983;
  wire [0:0] v_17984;
  wire [0:0] v_17985;
  wire [0:0] v_17986;
  wire [0:0] v_17987;
  wire [0:0] v_17988;
  wire [0:0] v_17989;
  function [0:0] mux_17989(input [0:0] sel);
    case (sel) 0: mux_17989 = 1'h0; 1: mux_17989 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17990;
  function [0:0] mux_17990(input [0:0] sel);
    case (sel) 0: mux_17990 = 1'h0; 1: mux_17990 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17991;
  wire [0:0] v_17992;
  wire [0:0] v_17993;
  wire [0:0] v_17994;
  function [0:0] mux_17994(input [0:0] sel);
    case (sel) 0: mux_17994 = 1'h0; 1: mux_17994 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_17995;
  function [0:0] mux_17995(input [0:0] sel);
    case (sel) 0: mux_17995 = 1'h0; 1: mux_17995 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_17996;
  wire [0:0] v_17997;
  wire [0:0] v_17998;
  wire [0:0] v_17999;
  wire [0:0] v_18000;
  wire [0:0] v_18001;
  function [0:0] mux_18001(input [0:0] sel);
    case (sel) 0: mux_18001 = 1'h0; 1: mux_18001 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18002;
  function [0:0] mux_18002(input [0:0] sel);
    case (sel) 0: mux_18002 = 1'h0; 1: mux_18002 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18003;
  wire [0:0] v_18004;
  wire [0:0] v_18005;
  wire [0:0] v_18006;
  function [0:0] mux_18006(input [0:0] sel);
    case (sel) 0: mux_18006 = 1'h0; 1: mux_18006 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18007;
  function [0:0] mux_18007(input [0:0] sel);
    case (sel) 0: mux_18007 = 1'h0; 1: mux_18007 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18008;
  wire [0:0] v_18009;
  wire [0:0] v_18010;
  wire [0:0] v_18011;
  wire [0:0] v_18012;
  wire [0:0] v_18013;
  function [0:0] mux_18013(input [0:0] sel);
    case (sel) 0: mux_18013 = 1'h0; 1: mux_18013 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18014;
  wire [0:0] v_18015;
  wire [0:0] v_18016;
  wire [0:0] v_18017;
  wire [0:0] v_18018;
  function [0:0] mux_18018(input [0:0] sel);
    case (sel) 0: mux_18018 = 1'h0; 1: mux_18018 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18019;
  wire [0:0] v_18020;
  wire [0:0] v_18021;
  wire [0:0] v_18022;
  function [0:0] mux_18022(input [0:0] sel);
    case (sel) 0: mux_18022 = 1'h0; 1: mux_18022 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18023;
  function [0:0] mux_18023(input [0:0] sel);
    case (sel) 0: mux_18023 = 1'h0; 1: mux_18023 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_18024 = 1'h0;
  wire [0:0] v_18025;
  wire [0:0] v_18026;
  wire [0:0] act_18027;
  wire [0:0] v_18028;
  wire [0:0] v_18029;
  wire [0:0] v_18030;
  reg [0:0] v_18031 = 1'h0;
  wire [0:0] v_18032;
  wire [0:0] v_18033;
  wire [0:0] act_18034;
  wire [0:0] v_18035;
  wire [0:0] v_18036;
  wire [0:0] v_18037;
  reg [0:0] v_18038 = 1'h0;
  wire [0:0] v_18039;
  wire [0:0] v_18040;
  wire [0:0] act_18041;
  wire [0:0] v_18042;
  wire [0:0] v_18043;
  wire [0:0] v_18044;
  wire [0:0] vin0_consume_en_18045;
  wire [0:0] vout_canPeek_18045;
  wire [7:0] vout_peek_18045;
  wire [0:0] v_18046;
  wire [0:0] v_18047;
  function [0:0] mux_18047(input [0:0] sel);
    case (sel) 0: mux_18047 = 1'h0; 1: mux_18047 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18048;
  wire [0:0] v_18049;
  wire [0:0] v_18050;
  wire [0:0] v_18051;
  wire [0:0] v_18052;
  function [0:0] mux_18052(input [0:0] sel);
    case (sel) 0: mux_18052 = 1'h0; 1: mux_18052 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18053;
  wire [0:0] vin0_consume_en_18054;
  wire [0:0] vout_canPeek_18054;
  wire [7:0] vout_peek_18054;
  wire [0:0] v_18055;
  wire [0:0] v_18056;
  function [0:0] mux_18056(input [0:0] sel);
    case (sel) 0: mux_18056 = 1'h0; 1: mux_18056 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18057;
  function [0:0] mux_18057(input [0:0] sel);
    case (sel) 0: mux_18057 = 1'h0; 1: mux_18057 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18058;
  wire [0:0] v_18059;
  wire [0:0] v_18060;
  wire [0:0] v_18061;
  wire [0:0] v_18062;
  wire [0:0] v_18063;
  wire [0:0] v_18064;
  function [0:0] mux_18064(input [0:0] sel);
    case (sel) 0: mux_18064 = 1'h0; 1: mux_18064 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18065;
  wire [0:0] v_18066;
  wire [0:0] v_18067;
  wire [0:0] v_18068;
  wire [0:0] v_18069;
  function [0:0] mux_18069(input [0:0] sel);
    case (sel) 0: mux_18069 = 1'h0; 1: mux_18069 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18070;
  wire [0:0] v_18071;
  wire [0:0] v_18072;
  wire [0:0] v_18073;
  function [0:0] mux_18073(input [0:0] sel);
    case (sel) 0: mux_18073 = 1'h0; 1: mux_18073 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18074;
  function [0:0] mux_18074(input [0:0] sel);
    case (sel) 0: mux_18074 = 1'h0; 1: mux_18074 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_18075 = 1'h0;
  wire [0:0] v_18076;
  wire [0:0] v_18077;
  wire [0:0] act_18078;
  wire [0:0] v_18079;
  wire [0:0] v_18080;
  wire [0:0] v_18081;
  wire [0:0] vin0_consume_en_18082;
  wire [0:0] vout_canPeek_18082;
  wire [7:0] vout_peek_18082;
  wire [0:0] v_18083;
  wire [0:0] v_18084;
  function [0:0] mux_18084(input [0:0] sel);
    case (sel) 0: mux_18084 = 1'h0; 1: mux_18084 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18085;
  wire [0:0] v_18086;
  wire [0:0] v_18087;
  wire [0:0] v_18088;
  wire [0:0] v_18089;
  function [0:0] mux_18089(input [0:0] sel);
    case (sel) 0: mux_18089 = 1'h0; 1: mux_18089 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18090;
  wire [0:0] vin0_consume_en_18091;
  wire [0:0] vout_canPeek_18091;
  wire [7:0] vout_peek_18091;
  wire [0:0] v_18092;
  wire [0:0] v_18093;
  function [0:0] mux_18093(input [0:0] sel);
    case (sel) 0: mux_18093 = 1'h0; 1: mux_18093 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18094;
  function [0:0] mux_18094(input [0:0] sel);
    case (sel) 0: mux_18094 = 1'h0; 1: mux_18094 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18095;
  wire [0:0] v_18096;
  wire [0:0] v_18097;
  wire [0:0] v_18098;
  wire [0:0] v_18099;
  wire [0:0] v_18100;
  wire [0:0] v_18101;
  function [0:0] mux_18101(input [0:0] sel);
    case (sel) 0: mux_18101 = 1'h0; 1: mux_18101 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18102;
  function [0:0] mux_18102(input [0:0] sel);
    case (sel) 0: mux_18102 = 1'h0; 1: mux_18102 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18103;
  wire [0:0] v_18104;
  wire [0:0] v_18105;
  wire [0:0] v_18106;
  function [0:0] mux_18106(input [0:0] sel);
    case (sel) 0: mux_18106 = 1'h0; 1: mux_18106 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18107;
  function [0:0] mux_18107(input [0:0] sel);
    case (sel) 0: mux_18107 = 1'h0; 1: mux_18107 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18108;
  wire [0:0] v_18109;
  wire [0:0] v_18110;
  wire [0:0] v_18111;
  wire [0:0] v_18112;
  wire [0:0] v_18113;
  function [0:0] mux_18113(input [0:0] sel);
    case (sel) 0: mux_18113 = 1'h0; 1: mux_18113 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18114;
  wire [0:0] v_18115;
  wire [0:0] v_18116;
  wire [0:0] v_18117;
  wire [0:0] v_18118;
  function [0:0] mux_18118(input [0:0] sel);
    case (sel) 0: mux_18118 = 1'h0; 1: mux_18118 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18119;
  wire [0:0] v_18120;
  wire [0:0] v_18121;
  wire [0:0] v_18122;
  function [0:0] mux_18122(input [0:0] sel);
    case (sel) 0: mux_18122 = 1'h0; 1: mux_18122 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18123;
  function [0:0] mux_18123(input [0:0] sel);
    case (sel) 0: mux_18123 = 1'h0; 1: mux_18123 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_18124 = 1'h0;
  wire [0:0] v_18125;
  wire [0:0] v_18126;
  wire [0:0] act_18127;
  wire [0:0] v_18128;
  wire [0:0] v_18129;
  wire [0:0] v_18130;
  reg [0:0] v_18131 = 1'h0;
  wire [0:0] v_18132;
  wire [0:0] v_18133;
  wire [0:0] act_18134;
  wire [0:0] v_18135;
  wire [0:0] v_18136;
  wire [0:0] v_18137;
  wire [0:0] vin0_consume_en_18138;
  wire [0:0] vout_canPeek_18138;
  wire [7:0] vout_peek_18138;
  wire [0:0] v_18139;
  wire [0:0] v_18140;
  function [0:0] mux_18140(input [0:0] sel);
    case (sel) 0: mux_18140 = 1'h0; 1: mux_18140 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18141;
  wire [0:0] v_18142;
  wire [0:0] v_18143;
  wire [0:0] v_18144;
  wire [0:0] v_18145;
  function [0:0] mux_18145(input [0:0] sel);
    case (sel) 0: mux_18145 = 1'h0; 1: mux_18145 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18146;
  wire [0:0] vin0_consume_en_18147;
  wire [0:0] vout_canPeek_18147;
  wire [7:0] vout_peek_18147;
  wire [0:0] v_18148;
  wire [0:0] v_18149;
  function [0:0] mux_18149(input [0:0] sel);
    case (sel) 0: mux_18149 = 1'h0; 1: mux_18149 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18150;
  function [0:0] mux_18150(input [0:0] sel);
    case (sel) 0: mux_18150 = 1'h0; 1: mux_18150 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18151;
  wire [0:0] v_18152;
  wire [0:0] v_18153;
  wire [0:0] v_18154;
  wire [0:0] v_18155;
  wire [0:0] v_18156;
  wire [0:0] v_18157;
  function [0:0] mux_18157(input [0:0] sel);
    case (sel) 0: mux_18157 = 1'h0; 1: mux_18157 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18158;
  wire [0:0] v_18159;
  wire [0:0] v_18160;
  wire [0:0] v_18161;
  wire [0:0] v_18162;
  function [0:0] mux_18162(input [0:0] sel);
    case (sel) 0: mux_18162 = 1'h0; 1: mux_18162 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18163;
  wire [0:0] v_18164;
  wire [0:0] v_18165;
  wire [0:0] v_18166;
  function [0:0] mux_18166(input [0:0] sel);
    case (sel) 0: mux_18166 = 1'h0; 1: mux_18166 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18167;
  function [0:0] mux_18167(input [0:0] sel);
    case (sel) 0: mux_18167 = 1'h0; 1: mux_18167 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_18168 = 1'h0;
  wire [0:0] v_18169;
  wire [0:0] v_18170;
  wire [0:0] act_18171;
  wire [0:0] v_18172;
  wire [0:0] v_18173;
  wire [0:0] v_18174;
  wire [0:0] vin0_consume_en_18175;
  wire [0:0] vout_canPeek_18175;
  wire [7:0] vout_peek_18175;
  wire [0:0] v_18176;
  wire [0:0] v_18177;
  function [0:0] mux_18177(input [0:0] sel);
    case (sel) 0: mux_18177 = 1'h0; 1: mux_18177 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18178;
  wire [0:0] v_18179;
  wire [0:0] v_18180;
  wire [0:0] v_18181;
  wire [0:0] v_18182;
  function [0:0] mux_18182(input [0:0] sel);
    case (sel) 0: mux_18182 = 1'h0; 1: mux_18182 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18183;
  wire [0:0] vin0_consume_en_18184;
  wire [0:0] vout_canPeek_18184;
  wire [7:0] vout_peek_18184;
  wire [0:0] v_18185;
  wire [0:0] v_18186;
  function [0:0] mux_18186(input [0:0] sel);
    case (sel) 0: mux_18186 = 1'h0; 1: mux_18186 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18187;
  function [0:0] mux_18187(input [0:0] sel);
    case (sel) 0: mux_18187 = 1'h0; 1: mux_18187 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18188;
  wire [0:0] v_18189;
  wire [0:0] v_18190;
  wire [0:0] v_18191;
  wire [0:0] v_18192;
  wire [0:0] v_18193;
  wire [0:0] v_18194;
  function [0:0] mux_18194(input [0:0] sel);
    case (sel) 0: mux_18194 = 1'h0; 1: mux_18194 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18195;
  function [0:0] mux_18195(input [0:0] sel);
    case (sel) 0: mux_18195 = 1'h0; 1: mux_18195 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18196;
  wire [0:0] v_18197;
  wire [0:0] v_18198;
  wire [0:0] v_18199;
  function [0:0] mux_18199(input [0:0] sel);
    case (sel) 0: mux_18199 = 1'h0; 1: mux_18199 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18200;
  function [0:0] mux_18200(input [0:0] sel);
    case (sel) 0: mux_18200 = 1'h0; 1: mux_18200 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18201;
  wire [0:0] v_18202;
  wire [0:0] v_18203;
  wire [0:0] v_18204;
  wire [0:0] v_18205;
  wire [0:0] v_18206;
  function [0:0] mux_18206(input [0:0] sel);
    case (sel) 0: mux_18206 = 1'h0; 1: mux_18206 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18207;
  function [0:0] mux_18207(input [0:0] sel);
    case (sel) 0: mux_18207 = 1'h0; 1: mux_18207 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18208;
  wire [0:0] v_18209;
  wire [0:0] v_18210;
  wire [0:0] v_18211;
  function [0:0] mux_18211(input [0:0] sel);
    case (sel) 0: mux_18211 = 1'h0; 1: mux_18211 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18212;
  function [0:0] mux_18212(input [0:0] sel);
    case (sel) 0: mux_18212 = 1'h0; 1: mux_18212 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18213;
  wire [0:0] v_18214;
  wire [0:0] v_18215;
  wire [0:0] v_18216;
  wire [0:0] v_18217;
  wire [0:0] v_18218;
  function [0:0] mux_18218(input [0:0] sel);
    case (sel) 0: mux_18218 = 1'h0; 1: mux_18218 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18219;
  function [0:0] mux_18219(input [0:0] sel);
    case (sel) 0: mux_18219 = 1'h0; 1: mux_18219 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18220;
  wire [0:0] v_18221;
  wire [0:0] v_18222;
  wire [0:0] v_18223;
  function [0:0] mux_18223(input [0:0] sel);
    case (sel) 0: mux_18223 = 1'h0; 1: mux_18223 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18224;
  function [0:0] mux_18224(input [0:0] sel);
    case (sel) 0: mux_18224 = 1'h0; 1: mux_18224 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18225;
  wire [0:0] v_18226;
  wire [0:0] v_18227;
  wire [0:0] v_18228;
  wire [0:0] v_18229;
  wire [0:0] v_18230;
  function [0:0] mux_18230(input [0:0] sel);
    case (sel) 0: mux_18230 = 1'h0; 1: mux_18230 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18231;
  wire [0:0] v_18232;
  wire [0:0] v_18233;
  wire [0:0] v_18234;
  wire [0:0] v_18235;
  function [0:0] mux_18235(input [0:0] sel);
    case (sel) 0: mux_18235 = 1'h0; 1: mux_18235 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18236;
  wire [0:0] v_18237;
  wire [0:0] v_18238;
  wire [0:0] v_18239;
  function [0:0] mux_18239(input [0:0] sel);
    case (sel) 0: mux_18239 = 1'h0; 1: mux_18239 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18240;
  function [0:0] mux_18240(input [0:0] sel);
    case (sel) 0: mux_18240 = 1'h0; 1: mux_18240 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_18241 = 1'h0;
  wire [0:0] v_18242;
  wire [0:0] v_18243;
  wire [0:0] act_18244;
  wire [0:0] v_18245;
  wire [0:0] v_18246;
  wire [0:0] v_18247;
  reg [0:0] v_18248 = 1'h0;
  wire [0:0] v_18249;
  wire [0:0] v_18250;
  wire [0:0] act_18251;
  wire [0:0] v_18252;
  wire [0:0] v_18253;
  wire [0:0] v_18254;
  reg [0:0] v_18255 = 1'h0;
  wire [0:0] v_18256;
  wire [0:0] v_18257;
  wire [0:0] act_18258;
  wire [0:0] v_18259;
  wire [0:0] v_18260;
  wire [0:0] v_18261;
  reg [0:0] v_18262 = 1'h0;
  wire [0:0] v_18263;
  wire [0:0] v_18264;
  wire [0:0] act_18265;
  wire [0:0] v_18266;
  wire [0:0] v_18267;
  wire [0:0] v_18268;
  wire [0:0] vin0_consume_en_18269;
  wire [0:0] vout_canPeek_18269;
  wire [7:0] vout_peek_18269;
  wire [0:0] v_18270;
  wire [0:0] v_18271;
  function [0:0] mux_18271(input [0:0] sel);
    case (sel) 0: mux_18271 = 1'h0; 1: mux_18271 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18272;
  wire [0:0] v_18273;
  wire [0:0] v_18274;
  wire [0:0] v_18275;
  wire [0:0] v_18276;
  function [0:0] mux_18276(input [0:0] sel);
    case (sel) 0: mux_18276 = 1'h0; 1: mux_18276 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18277;
  wire [0:0] vin0_consume_en_18278;
  wire [0:0] vout_canPeek_18278;
  wire [7:0] vout_peek_18278;
  wire [0:0] v_18279;
  wire [0:0] v_18280;
  function [0:0] mux_18280(input [0:0] sel);
    case (sel) 0: mux_18280 = 1'h0; 1: mux_18280 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18281;
  function [0:0] mux_18281(input [0:0] sel);
    case (sel) 0: mux_18281 = 1'h0; 1: mux_18281 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18282;
  wire [0:0] v_18283;
  wire [0:0] v_18284;
  wire [0:0] v_18285;
  wire [0:0] v_18286;
  wire [0:0] v_18287;
  wire [0:0] v_18288;
  function [0:0] mux_18288(input [0:0] sel);
    case (sel) 0: mux_18288 = 1'h0; 1: mux_18288 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18289;
  wire [0:0] v_18290;
  wire [0:0] v_18291;
  wire [0:0] v_18292;
  wire [0:0] v_18293;
  function [0:0] mux_18293(input [0:0] sel);
    case (sel) 0: mux_18293 = 1'h0; 1: mux_18293 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18294;
  wire [0:0] v_18295;
  wire [0:0] v_18296;
  wire [0:0] v_18297;
  function [0:0] mux_18297(input [0:0] sel);
    case (sel) 0: mux_18297 = 1'h0; 1: mux_18297 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18298;
  function [0:0] mux_18298(input [0:0] sel);
    case (sel) 0: mux_18298 = 1'h0; 1: mux_18298 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_18299 = 1'h0;
  wire [0:0] v_18300;
  wire [0:0] v_18301;
  wire [0:0] act_18302;
  wire [0:0] v_18303;
  wire [0:0] v_18304;
  wire [0:0] v_18305;
  wire [0:0] vin0_consume_en_18306;
  wire [0:0] vout_canPeek_18306;
  wire [7:0] vout_peek_18306;
  wire [0:0] v_18307;
  wire [0:0] v_18308;
  function [0:0] mux_18308(input [0:0] sel);
    case (sel) 0: mux_18308 = 1'h0; 1: mux_18308 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18309;
  wire [0:0] v_18310;
  wire [0:0] v_18311;
  wire [0:0] v_18312;
  wire [0:0] v_18313;
  function [0:0] mux_18313(input [0:0] sel);
    case (sel) 0: mux_18313 = 1'h0; 1: mux_18313 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18314;
  wire [0:0] vin0_consume_en_18315;
  wire [0:0] vout_canPeek_18315;
  wire [7:0] vout_peek_18315;
  wire [0:0] v_18316;
  wire [0:0] v_18317;
  function [0:0] mux_18317(input [0:0] sel);
    case (sel) 0: mux_18317 = 1'h0; 1: mux_18317 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18318;
  function [0:0] mux_18318(input [0:0] sel);
    case (sel) 0: mux_18318 = 1'h0; 1: mux_18318 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18319;
  wire [0:0] v_18320;
  wire [0:0] v_18321;
  wire [0:0] v_18322;
  wire [0:0] v_18323;
  wire [0:0] v_18324;
  wire [0:0] v_18325;
  function [0:0] mux_18325(input [0:0] sel);
    case (sel) 0: mux_18325 = 1'h0; 1: mux_18325 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18326;
  function [0:0] mux_18326(input [0:0] sel);
    case (sel) 0: mux_18326 = 1'h0; 1: mux_18326 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18327;
  wire [0:0] v_18328;
  wire [0:0] v_18329;
  wire [0:0] v_18330;
  function [0:0] mux_18330(input [0:0] sel);
    case (sel) 0: mux_18330 = 1'h0; 1: mux_18330 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18331;
  function [0:0] mux_18331(input [0:0] sel);
    case (sel) 0: mux_18331 = 1'h0; 1: mux_18331 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18332;
  wire [0:0] v_18333;
  wire [0:0] v_18334;
  wire [0:0] v_18335;
  wire [0:0] v_18336;
  wire [0:0] v_18337;
  function [0:0] mux_18337(input [0:0] sel);
    case (sel) 0: mux_18337 = 1'h0; 1: mux_18337 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18338;
  wire [0:0] v_18339;
  wire [0:0] v_18340;
  wire [0:0] v_18341;
  wire [0:0] v_18342;
  function [0:0] mux_18342(input [0:0] sel);
    case (sel) 0: mux_18342 = 1'h0; 1: mux_18342 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18343;
  wire [0:0] v_18344;
  wire [0:0] v_18345;
  wire [0:0] v_18346;
  function [0:0] mux_18346(input [0:0] sel);
    case (sel) 0: mux_18346 = 1'h0; 1: mux_18346 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18347;
  function [0:0] mux_18347(input [0:0] sel);
    case (sel) 0: mux_18347 = 1'h0; 1: mux_18347 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_18348 = 1'h0;
  wire [0:0] v_18349;
  wire [0:0] v_18350;
  wire [0:0] act_18351;
  wire [0:0] v_18352;
  wire [0:0] v_18353;
  wire [0:0] v_18354;
  reg [0:0] v_18355 = 1'h0;
  wire [0:0] v_18356;
  wire [0:0] v_18357;
  wire [0:0] act_18358;
  wire [0:0] v_18359;
  wire [0:0] v_18360;
  wire [0:0] v_18361;
  wire [0:0] vin0_consume_en_18362;
  wire [0:0] vout_canPeek_18362;
  wire [7:0] vout_peek_18362;
  wire [0:0] v_18363;
  wire [0:0] v_18364;
  function [0:0] mux_18364(input [0:0] sel);
    case (sel) 0: mux_18364 = 1'h0; 1: mux_18364 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18365;
  wire [0:0] v_18366;
  wire [0:0] v_18367;
  wire [0:0] v_18368;
  wire [0:0] v_18369;
  function [0:0] mux_18369(input [0:0] sel);
    case (sel) 0: mux_18369 = 1'h0; 1: mux_18369 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18370;
  wire [0:0] vin0_consume_en_18371;
  wire [0:0] vout_canPeek_18371;
  wire [7:0] vout_peek_18371;
  wire [0:0] v_18372;
  wire [0:0] v_18373;
  function [0:0] mux_18373(input [0:0] sel);
    case (sel) 0: mux_18373 = 1'h0; 1: mux_18373 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18374;
  function [0:0] mux_18374(input [0:0] sel);
    case (sel) 0: mux_18374 = 1'h0; 1: mux_18374 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18375;
  wire [0:0] v_18376;
  wire [0:0] v_18377;
  wire [0:0] v_18378;
  wire [0:0] v_18379;
  wire [0:0] v_18380;
  wire [0:0] v_18381;
  function [0:0] mux_18381(input [0:0] sel);
    case (sel) 0: mux_18381 = 1'h0; 1: mux_18381 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18382;
  wire [0:0] v_18383;
  wire [0:0] v_18384;
  wire [0:0] v_18385;
  wire [0:0] v_18386;
  function [0:0] mux_18386(input [0:0] sel);
    case (sel) 0: mux_18386 = 1'h0; 1: mux_18386 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18387;
  wire [0:0] v_18388;
  wire [0:0] v_18389;
  wire [0:0] v_18390;
  function [0:0] mux_18390(input [0:0] sel);
    case (sel) 0: mux_18390 = 1'h0; 1: mux_18390 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18391;
  function [0:0] mux_18391(input [0:0] sel);
    case (sel) 0: mux_18391 = 1'h0; 1: mux_18391 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_18392 = 1'h0;
  wire [0:0] v_18393;
  wire [0:0] v_18394;
  wire [0:0] act_18395;
  wire [0:0] v_18396;
  wire [0:0] v_18397;
  wire [0:0] v_18398;
  wire [0:0] vin0_consume_en_18399;
  wire [0:0] vout_canPeek_18399;
  wire [7:0] vout_peek_18399;
  wire [0:0] v_18400;
  wire [0:0] v_18401;
  function [0:0] mux_18401(input [0:0] sel);
    case (sel) 0: mux_18401 = 1'h0; 1: mux_18401 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18402;
  wire [0:0] v_18403;
  wire [0:0] v_18404;
  wire [0:0] v_18405;
  wire [0:0] v_18406;
  function [0:0] mux_18406(input [0:0] sel);
    case (sel) 0: mux_18406 = 1'h0; 1: mux_18406 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18407;
  wire [0:0] vin0_consume_en_18408;
  wire [0:0] vout_canPeek_18408;
  wire [7:0] vout_peek_18408;
  wire [0:0] v_18409;
  wire [0:0] v_18410;
  function [0:0] mux_18410(input [0:0] sel);
    case (sel) 0: mux_18410 = 1'h0; 1: mux_18410 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18411;
  function [0:0] mux_18411(input [0:0] sel);
    case (sel) 0: mux_18411 = 1'h0; 1: mux_18411 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18412;
  wire [0:0] v_18413;
  wire [0:0] v_18414;
  wire [0:0] v_18415;
  wire [0:0] v_18416;
  wire [0:0] v_18417;
  wire [0:0] v_18418;
  function [0:0] mux_18418(input [0:0] sel);
    case (sel) 0: mux_18418 = 1'h0; 1: mux_18418 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18419;
  function [0:0] mux_18419(input [0:0] sel);
    case (sel) 0: mux_18419 = 1'h0; 1: mux_18419 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18420;
  wire [0:0] v_18421;
  wire [0:0] v_18422;
  wire [0:0] v_18423;
  function [0:0] mux_18423(input [0:0] sel);
    case (sel) 0: mux_18423 = 1'h0; 1: mux_18423 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18424;
  function [0:0] mux_18424(input [0:0] sel);
    case (sel) 0: mux_18424 = 1'h0; 1: mux_18424 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18425;
  wire [0:0] v_18426;
  wire [0:0] v_18427;
  wire [0:0] v_18428;
  wire [0:0] v_18429;
  wire [0:0] v_18430;
  function [0:0] mux_18430(input [0:0] sel);
    case (sel) 0: mux_18430 = 1'h0; 1: mux_18430 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18431;
  function [0:0] mux_18431(input [0:0] sel);
    case (sel) 0: mux_18431 = 1'h0; 1: mux_18431 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18432;
  wire [0:0] v_18433;
  wire [0:0] v_18434;
  wire [0:0] v_18435;
  function [0:0] mux_18435(input [0:0] sel);
    case (sel) 0: mux_18435 = 1'h0; 1: mux_18435 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18436;
  function [0:0] mux_18436(input [0:0] sel);
    case (sel) 0: mux_18436 = 1'h0; 1: mux_18436 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18437;
  wire [0:0] v_18438;
  wire [0:0] v_18439;
  wire [0:0] v_18440;
  wire [0:0] v_18441;
  wire [0:0] v_18442;
  function [0:0] mux_18442(input [0:0] sel);
    case (sel) 0: mux_18442 = 1'h0; 1: mux_18442 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18443;
  wire [0:0] v_18444;
  wire [0:0] v_18445;
  wire [0:0] v_18446;
  wire [0:0] v_18447;
  function [0:0] mux_18447(input [0:0] sel);
    case (sel) 0: mux_18447 = 1'h0; 1: mux_18447 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18448;
  wire [0:0] v_18449;
  wire [0:0] v_18450;
  wire [0:0] v_18451;
  function [0:0] mux_18451(input [0:0] sel);
    case (sel) 0: mux_18451 = 1'h0; 1: mux_18451 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18452;
  function [0:0] mux_18452(input [0:0] sel);
    case (sel) 0: mux_18452 = 1'h0; 1: mux_18452 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_18453 = 1'h0;
  wire [0:0] v_18454;
  wire [0:0] v_18455;
  wire [0:0] act_18456;
  wire [0:0] v_18457;
  wire [0:0] v_18458;
  wire [0:0] v_18459;
  reg [0:0] v_18460 = 1'h0;
  wire [0:0] v_18461;
  wire [0:0] v_18462;
  wire [0:0] act_18463;
  wire [0:0] v_18464;
  wire [0:0] v_18465;
  wire [0:0] v_18466;
  reg [0:0] v_18467 = 1'h0;
  wire [0:0] v_18468;
  wire [0:0] v_18469;
  wire [0:0] act_18470;
  wire [0:0] v_18471;
  wire [0:0] v_18472;
  wire [0:0] v_18473;
  wire [0:0] vin0_consume_en_18474;
  wire [0:0] vout_canPeek_18474;
  wire [7:0] vout_peek_18474;
  wire [0:0] v_18475;
  wire [0:0] v_18476;
  function [0:0] mux_18476(input [0:0] sel);
    case (sel) 0: mux_18476 = 1'h0; 1: mux_18476 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18477;
  wire [0:0] v_18478;
  wire [0:0] v_18479;
  wire [0:0] v_18480;
  wire [0:0] v_18481;
  function [0:0] mux_18481(input [0:0] sel);
    case (sel) 0: mux_18481 = 1'h0; 1: mux_18481 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18482;
  wire [0:0] vin0_consume_en_18483;
  wire [0:0] vout_canPeek_18483;
  wire [7:0] vout_peek_18483;
  wire [0:0] v_18484;
  wire [0:0] v_18485;
  function [0:0] mux_18485(input [0:0] sel);
    case (sel) 0: mux_18485 = 1'h0; 1: mux_18485 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18486;
  function [0:0] mux_18486(input [0:0] sel);
    case (sel) 0: mux_18486 = 1'h0; 1: mux_18486 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18487;
  wire [0:0] v_18488;
  wire [0:0] v_18489;
  wire [0:0] v_18490;
  wire [0:0] v_18491;
  wire [0:0] v_18492;
  wire [0:0] v_18493;
  function [0:0] mux_18493(input [0:0] sel);
    case (sel) 0: mux_18493 = 1'h0; 1: mux_18493 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18494;
  wire [0:0] v_18495;
  wire [0:0] v_18496;
  wire [0:0] v_18497;
  wire [0:0] v_18498;
  function [0:0] mux_18498(input [0:0] sel);
    case (sel) 0: mux_18498 = 1'h0; 1: mux_18498 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18499;
  wire [0:0] v_18500;
  wire [0:0] v_18501;
  wire [0:0] v_18502;
  function [0:0] mux_18502(input [0:0] sel);
    case (sel) 0: mux_18502 = 1'h0; 1: mux_18502 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18503;
  function [0:0] mux_18503(input [0:0] sel);
    case (sel) 0: mux_18503 = 1'h0; 1: mux_18503 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_18504 = 1'h0;
  wire [0:0] v_18505;
  wire [0:0] v_18506;
  wire [0:0] act_18507;
  wire [0:0] v_18508;
  wire [0:0] v_18509;
  wire [0:0] v_18510;
  wire [0:0] vin0_consume_en_18511;
  wire [0:0] vout_canPeek_18511;
  wire [7:0] vout_peek_18511;
  wire [0:0] v_18512;
  wire [0:0] v_18513;
  function [0:0] mux_18513(input [0:0] sel);
    case (sel) 0: mux_18513 = 1'h0; 1: mux_18513 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18514;
  wire [0:0] v_18515;
  wire [0:0] v_18516;
  wire [0:0] v_18517;
  wire [0:0] v_18518;
  function [0:0] mux_18518(input [0:0] sel);
    case (sel) 0: mux_18518 = 1'h0; 1: mux_18518 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18519;
  wire [0:0] vin0_consume_en_18520;
  wire [0:0] vout_canPeek_18520;
  wire [7:0] vout_peek_18520;
  wire [0:0] v_18521;
  wire [0:0] v_18522;
  function [0:0] mux_18522(input [0:0] sel);
    case (sel) 0: mux_18522 = 1'h0; 1: mux_18522 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18523;
  function [0:0] mux_18523(input [0:0] sel);
    case (sel) 0: mux_18523 = 1'h0; 1: mux_18523 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18524;
  wire [0:0] v_18525;
  wire [0:0] v_18526;
  wire [0:0] v_18527;
  wire [0:0] v_18528;
  wire [0:0] v_18529;
  wire [0:0] v_18530;
  function [0:0] mux_18530(input [0:0] sel);
    case (sel) 0: mux_18530 = 1'h0; 1: mux_18530 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18531;
  function [0:0] mux_18531(input [0:0] sel);
    case (sel) 0: mux_18531 = 1'h0; 1: mux_18531 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18532;
  wire [0:0] v_18533;
  wire [0:0] v_18534;
  wire [0:0] v_18535;
  function [0:0] mux_18535(input [0:0] sel);
    case (sel) 0: mux_18535 = 1'h0; 1: mux_18535 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18536;
  function [0:0] mux_18536(input [0:0] sel);
    case (sel) 0: mux_18536 = 1'h0; 1: mux_18536 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18537;
  wire [0:0] v_18538;
  wire [0:0] v_18539;
  wire [0:0] v_18540;
  wire [0:0] v_18541;
  wire [0:0] v_18542;
  function [0:0] mux_18542(input [0:0] sel);
    case (sel) 0: mux_18542 = 1'h0; 1: mux_18542 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18543;
  wire [0:0] v_18544;
  wire [0:0] v_18545;
  wire [0:0] v_18546;
  wire [0:0] v_18547;
  function [0:0] mux_18547(input [0:0] sel);
    case (sel) 0: mux_18547 = 1'h0; 1: mux_18547 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18548;
  wire [0:0] v_18549;
  wire [0:0] v_18550;
  wire [0:0] v_18551;
  function [0:0] mux_18551(input [0:0] sel);
    case (sel) 0: mux_18551 = 1'h0; 1: mux_18551 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18552;
  function [0:0] mux_18552(input [0:0] sel);
    case (sel) 0: mux_18552 = 1'h0; 1: mux_18552 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_18553 = 1'h0;
  wire [0:0] v_18554;
  wire [0:0] v_18555;
  wire [0:0] act_18556;
  wire [0:0] v_18557;
  wire [0:0] v_18558;
  wire [0:0] v_18559;
  reg [0:0] v_18560 = 1'h0;
  wire [0:0] v_18561;
  wire [0:0] v_18562;
  wire [0:0] act_18563;
  wire [0:0] v_18564;
  wire [0:0] v_18565;
  wire [0:0] v_18566;
  wire [0:0] vin0_consume_en_18567;
  wire [0:0] vout_canPeek_18567;
  wire [7:0] vout_peek_18567;
  wire [0:0] v_18568;
  wire [0:0] v_18569;
  function [0:0] mux_18569(input [0:0] sel);
    case (sel) 0: mux_18569 = 1'h0; 1: mux_18569 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18570;
  wire [0:0] v_18571;
  wire [0:0] v_18572;
  wire [0:0] v_18573;
  wire [0:0] v_18574;
  function [0:0] mux_18574(input [0:0] sel);
    case (sel) 0: mux_18574 = 1'h0; 1: mux_18574 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18575;
  wire [0:0] vin0_consume_en_18576;
  wire [0:0] vout_canPeek_18576;
  wire [7:0] vout_peek_18576;
  wire [0:0] v_18577;
  wire [0:0] v_18578;
  function [0:0] mux_18578(input [0:0] sel);
    case (sel) 0: mux_18578 = 1'h0; 1: mux_18578 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18579;
  function [0:0] mux_18579(input [0:0] sel);
    case (sel) 0: mux_18579 = 1'h0; 1: mux_18579 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18580;
  wire [0:0] v_18581;
  wire [0:0] v_18582;
  wire [0:0] v_18583;
  wire [0:0] v_18584;
  wire [0:0] v_18585;
  wire [0:0] v_18586;
  function [0:0] mux_18586(input [0:0] sel);
    case (sel) 0: mux_18586 = 1'h0; 1: mux_18586 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18587;
  wire [0:0] v_18588;
  wire [0:0] v_18589;
  wire [0:0] v_18590;
  wire [0:0] v_18591;
  function [0:0] mux_18591(input [0:0] sel);
    case (sel) 0: mux_18591 = 1'h0; 1: mux_18591 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18592;
  wire [0:0] v_18593;
  wire [0:0] v_18594;
  wire [0:0] v_18595;
  function [0:0] mux_18595(input [0:0] sel);
    case (sel) 0: mux_18595 = 1'h0; 1: mux_18595 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18596;
  function [0:0] mux_18596(input [0:0] sel);
    case (sel) 0: mux_18596 = 1'h0; 1: mux_18596 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_18597 = 1'h0;
  wire [0:0] v_18598;
  wire [0:0] v_18599;
  wire [0:0] act_18600;
  wire [0:0] v_18601;
  wire [0:0] v_18602;
  wire [0:0] v_18603;
  wire [0:0] vin0_consume_en_18604;
  wire [0:0] vout_canPeek_18604;
  wire [7:0] vout_peek_18604;
  wire [0:0] v_18605;
  wire [0:0] v_18606;
  function [0:0] mux_18606(input [0:0] sel);
    case (sel) 0: mux_18606 = 1'h0; 1: mux_18606 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18607;
  wire [0:0] v_18608;
  wire [0:0] v_18609;
  wire [0:0] v_18610;
  wire [0:0] v_18611;
  function [0:0] mux_18611(input [0:0] sel);
    case (sel) 0: mux_18611 = 1'h0; 1: mux_18611 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18612;
  wire [0:0] vin0_consume_en_18613;
  wire [0:0] vout_canPeek_18613;
  wire [7:0] vout_peek_18613;
  wire [0:0] v_18614;
  wire [0:0] v_18615;
  function [0:0] mux_18615(input [0:0] sel);
    case (sel) 0: mux_18615 = 1'h0; 1: mux_18615 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18616;
  function [0:0] mux_18616(input [0:0] sel);
    case (sel) 0: mux_18616 = 1'h0; 1: mux_18616 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18617;
  wire [0:0] v_18618;
  wire [0:0] v_18619;
  wire [0:0] v_18620;
  wire [0:0] v_18621;
  wire [0:0] v_18622;
  wire [0:0] v_18623;
  function [0:0] mux_18623(input [0:0] sel);
    case (sel) 0: mux_18623 = 1'h0; 1: mux_18623 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18624;
  function [0:0] mux_18624(input [0:0] sel);
    case (sel) 0: mux_18624 = 1'h0; 1: mux_18624 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18625;
  wire [0:0] v_18626;
  wire [0:0] v_18627;
  wire [0:0] v_18628;
  function [0:0] mux_18628(input [0:0] sel);
    case (sel) 0: mux_18628 = 1'h0; 1: mux_18628 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18629;
  function [0:0] mux_18629(input [0:0] sel);
    case (sel) 0: mux_18629 = 1'h0; 1: mux_18629 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18630;
  wire [0:0] v_18631;
  wire [0:0] v_18632;
  wire [0:0] v_18633;
  wire [0:0] v_18634;
  wire [0:0] v_18635;
  function [0:0] mux_18635(input [0:0] sel);
    case (sel) 0: mux_18635 = 1'h0; 1: mux_18635 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18636;
  function [0:0] mux_18636(input [0:0] sel);
    case (sel) 0: mux_18636 = 1'h0; 1: mux_18636 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18637;
  wire [0:0] v_18638;
  wire [0:0] v_18639;
  wire [0:0] v_18640;
  function [0:0] mux_18640(input [0:0] sel);
    case (sel) 0: mux_18640 = 1'h0; 1: mux_18640 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18641;
  function [0:0] mux_18641(input [0:0] sel);
    case (sel) 0: mux_18641 = 1'h0; 1: mux_18641 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18642;
  wire [0:0] v_18643;
  wire [0:0] v_18644;
  wire [0:0] v_18645;
  wire [0:0] v_18646;
  wire [0:0] v_18647;
  function [0:0] mux_18647(input [0:0] sel);
    case (sel) 0: mux_18647 = 1'h0; 1: mux_18647 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18648;
  function [0:0] mux_18648(input [0:0] sel);
    case (sel) 0: mux_18648 = 1'h0; 1: mux_18648 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18649;
  wire [0:0] v_18650;
  wire [0:0] v_18651;
  wire [0:0] v_18652;
  function [0:0] mux_18652(input [0:0] sel);
    case (sel) 0: mux_18652 = 1'h0; 1: mux_18652 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18653;
  function [0:0] mux_18653(input [0:0] sel);
    case (sel) 0: mux_18653 = 1'h0; 1: mux_18653 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18654;
  wire [0:0] v_18655;
  wire [0:0] v_18656;
  wire [0:0] v_18657;
  wire [0:0] v_18658;
  wire [0:0] v_18659;
  function [0:0] mux_18659(input [0:0] sel);
    case (sel) 0: mux_18659 = 1'h0; 1: mux_18659 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18660;
  function [0:0] mux_18660(input [0:0] sel);
    case (sel) 0: mux_18660 = 1'h0; 1: mux_18660 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18661;
  wire [0:0] v_18662;
  wire [0:0] v_18663;
  wire [0:0] v_18664;
  function [0:0] mux_18664(input [0:0] sel);
    case (sel) 0: mux_18664 = 1'h0; 1: mux_18664 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18665;
  function [0:0] mux_18665(input [0:0] sel);
    case (sel) 0: mux_18665 = 1'h0; 1: mux_18665 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18666;
  wire [0:0] v_18667;
  wire [0:0] v_18668;
  wire [0:0] v_18669;
  wire [0:0] v_18670;
  wire [0:0] v_18671;
  function [0:0] mux_18671(input [0:0] sel);
    case (sel) 0: mux_18671 = 1'h0; 1: mux_18671 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18672;
  function [0:0] mux_18672(input [0:0] sel);
    case (sel) 0: mux_18672 = 1'h0; 1: mux_18672 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18673;
  wire [0:0] v_18674;
  wire [0:0] v_18675;
  wire [0:0] v_18676;
  function [0:0] mux_18676(input [0:0] sel);
    case (sel) 0: mux_18676 = 1'h0; 1: mux_18676 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18677;
  function [0:0] mux_18677(input [0:0] sel);
    case (sel) 0: mux_18677 = 1'h0; 1: mux_18677 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18678;
  wire [0:0] v_18679;
  wire [0:0] v_18680;
  wire [0:0] v_18681;
  wire [0:0] v_18682;
  wire [0:0] v_18683;
  function [0:0] mux_18683(input [0:0] sel);
    case (sel) 0: mux_18683 = 1'h0; 1: mux_18683 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18684;
  function [0:0] mux_18684(input [0:0] sel);
    case (sel) 0: mux_18684 = 1'h0; 1: mux_18684 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18685;
  wire [0:0] v_18686;
  wire [0:0] v_18687;
  wire [0:0] v_18688;
  function [0:0] mux_18688(input [0:0] sel);
    case (sel) 0: mux_18688 = 1'h0; 1: mux_18688 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18689;
  function [0:0] mux_18689(input [0:0] sel);
    case (sel) 0: mux_18689 = 1'h0; 1: mux_18689 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18690;
  wire [0:0] v_18691;
  wire [0:0] v_18692;
  wire [0:0] v_18693;
  wire [0:0] v_18694;
  wire [0:0] v_18695;
  function [0:0] mux_18695(input [0:0] sel);
    case (sel) 0: mux_18695 = 1'h0; 1: mux_18695 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18696;
  wire [0:0] v_18697;
  wire [0:0] v_18698;
  wire [0:0] v_18699;
  wire [0:0] v_18700;
  function [0:0] mux_18700(input [0:0] sel);
    case (sel) 0: mux_18700 = 1'h0; 1: mux_18700 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18701;
  wire [0:0] v_18702;
  wire [0:0] v_18703;
  wire [0:0] v_18704;
  function [0:0] mux_18704(input [0:0] sel);
    case (sel) 0: mux_18704 = 1'h0; 1: mux_18704 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18705;
  function [0:0] mux_18705(input [0:0] sel);
    case (sel) 0: mux_18705 = 1'h0; 1: mux_18705 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_18706 = 1'h0;
  wire [0:0] v_18707;
  wire [0:0] v_18708;
  wire [0:0] act_18709;
  wire [0:0] v_18710;
  wire [0:0] v_18711;
  wire [0:0] v_18712;
  reg [0:0] v_18713 = 1'h0;
  wire [0:0] v_18714;
  wire [0:0] v_18715;
  wire [0:0] act_18716;
  wire [0:0] v_18717;
  wire [0:0] v_18718;
  wire [0:0] v_18719;
  reg [0:0] v_18720 = 1'h0;
  wire [0:0] v_18721;
  wire [0:0] v_18722;
  wire [0:0] act_18723;
  wire [0:0] v_18724;
  wire [0:0] v_18725;
  wire [0:0] v_18726;
  reg [0:0] v_18727 = 1'h0;
  wire [0:0] v_18728;
  wire [0:0] v_18729;
  wire [0:0] act_18730;
  wire [0:0] v_18731;
  wire [0:0] v_18732;
  wire [0:0] v_18733;
  reg [0:0] v_18734 = 1'h0;
  wire [0:0] v_18735;
  wire [0:0] v_18736;
  wire [0:0] act_18737;
  wire [0:0] v_18738;
  wire [0:0] v_18739;
  wire [0:0] v_18740;
  reg [0:0] v_18741 = 1'h0;
  wire [0:0] v_18742;
  wire [0:0] v_18743;
  wire [0:0] act_18744;
  wire [0:0] v_18745;
  wire [0:0] v_18746;
  wire [0:0] v_18747;
  reg [0:0] v_18748 = 1'h0;
  wire [0:0] v_18749;
  wire [0:0] v_18750;
  wire [0:0] act_18751;
  wire [0:0] v_18752;
  wire [0:0] v_18753;
  wire [0:0] v_18754;
  wire [0:0] vin0_consume_en_18755;
  wire [0:0] vout_canPeek_18755;
  wire [7:0] vout_peek_18755;
  wire [0:0] v_18756;
  wire [0:0] v_18757;
  function [0:0] mux_18757(input [0:0] sel);
    case (sel) 0: mux_18757 = 1'h0; 1: mux_18757 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18758;
  wire [0:0] v_18759;
  wire [0:0] v_18760;
  wire [0:0] v_18761;
  wire [0:0] v_18762;
  function [0:0] mux_18762(input [0:0] sel);
    case (sel) 0: mux_18762 = 1'h0; 1: mux_18762 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18763;
  wire [0:0] vin0_consume_en_18764;
  wire [0:0] vout_canPeek_18764;
  wire [7:0] vout_peek_18764;
  wire [0:0] v_18765;
  wire [0:0] v_18766;
  function [0:0] mux_18766(input [0:0] sel);
    case (sel) 0: mux_18766 = 1'h0; 1: mux_18766 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18767;
  function [0:0] mux_18767(input [0:0] sel);
    case (sel) 0: mux_18767 = 1'h0; 1: mux_18767 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18768;
  wire [0:0] v_18769;
  wire [0:0] v_18770;
  wire [0:0] v_18771;
  wire [0:0] v_18772;
  wire [0:0] v_18773;
  wire [0:0] v_18774;
  function [0:0] mux_18774(input [0:0] sel);
    case (sel) 0: mux_18774 = 1'h0; 1: mux_18774 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18775;
  wire [0:0] v_18776;
  wire [0:0] v_18777;
  wire [0:0] v_18778;
  wire [0:0] v_18779;
  function [0:0] mux_18779(input [0:0] sel);
    case (sel) 0: mux_18779 = 1'h0; 1: mux_18779 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18780;
  wire [0:0] v_18781;
  wire [0:0] v_18782;
  wire [0:0] v_18783;
  function [0:0] mux_18783(input [0:0] sel);
    case (sel) 0: mux_18783 = 1'h0; 1: mux_18783 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18784;
  function [0:0] mux_18784(input [0:0] sel);
    case (sel) 0: mux_18784 = 1'h0; 1: mux_18784 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_18785 = 1'h0;
  wire [0:0] v_18786;
  wire [0:0] v_18787;
  wire [0:0] act_18788;
  wire [0:0] v_18789;
  wire [0:0] v_18790;
  wire [0:0] v_18791;
  wire [0:0] vin0_consume_en_18792;
  wire [0:0] vout_canPeek_18792;
  wire [7:0] vout_peek_18792;
  wire [0:0] v_18793;
  wire [0:0] v_18794;
  function [0:0] mux_18794(input [0:0] sel);
    case (sel) 0: mux_18794 = 1'h0; 1: mux_18794 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18795;
  wire [0:0] v_18796;
  wire [0:0] v_18797;
  wire [0:0] v_18798;
  wire [0:0] v_18799;
  function [0:0] mux_18799(input [0:0] sel);
    case (sel) 0: mux_18799 = 1'h0; 1: mux_18799 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18800;
  wire [0:0] vin0_consume_en_18801;
  wire [0:0] vout_canPeek_18801;
  wire [7:0] vout_peek_18801;
  wire [0:0] v_18802;
  wire [0:0] v_18803;
  function [0:0] mux_18803(input [0:0] sel);
    case (sel) 0: mux_18803 = 1'h0; 1: mux_18803 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18804;
  function [0:0] mux_18804(input [0:0] sel);
    case (sel) 0: mux_18804 = 1'h0; 1: mux_18804 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18805;
  wire [0:0] v_18806;
  wire [0:0] v_18807;
  wire [0:0] v_18808;
  wire [0:0] v_18809;
  wire [0:0] v_18810;
  wire [0:0] v_18811;
  function [0:0] mux_18811(input [0:0] sel);
    case (sel) 0: mux_18811 = 1'h0; 1: mux_18811 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18812;
  function [0:0] mux_18812(input [0:0] sel);
    case (sel) 0: mux_18812 = 1'h0; 1: mux_18812 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18813;
  wire [0:0] v_18814;
  wire [0:0] v_18815;
  wire [0:0] v_18816;
  function [0:0] mux_18816(input [0:0] sel);
    case (sel) 0: mux_18816 = 1'h0; 1: mux_18816 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18817;
  function [0:0] mux_18817(input [0:0] sel);
    case (sel) 0: mux_18817 = 1'h0; 1: mux_18817 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18818;
  wire [0:0] v_18819;
  wire [0:0] v_18820;
  wire [0:0] v_18821;
  wire [0:0] v_18822;
  wire [0:0] v_18823;
  function [0:0] mux_18823(input [0:0] sel);
    case (sel) 0: mux_18823 = 1'h0; 1: mux_18823 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18824;
  wire [0:0] v_18825;
  wire [0:0] v_18826;
  wire [0:0] v_18827;
  wire [0:0] v_18828;
  function [0:0] mux_18828(input [0:0] sel);
    case (sel) 0: mux_18828 = 1'h0; 1: mux_18828 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18829;
  wire [0:0] v_18830;
  wire [0:0] v_18831;
  wire [0:0] v_18832;
  function [0:0] mux_18832(input [0:0] sel);
    case (sel) 0: mux_18832 = 1'h0; 1: mux_18832 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18833;
  function [0:0] mux_18833(input [0:0] sel);
    case (sel) 0: mux_18833 = 1'h0; 1: mux_18833 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_18834 = 1'h0;
  wire [0:0] v_18835;
  wire [0:0] v_18836;
  wire [0:0] act_18837;
  wire [0:0] v_18838;
  wire [0:0] v_18839;
  wire [0:0] v_18840;
  reg [0:0] v_18841 = 1'h0;
  wire [0:0] v_18842;
  wire [0:0] v_18843;
  wire [0:0] act_18844;
  wire [0:0] v_18845;
  wire [0:0] v_18846;
  wire [0:0] v_18847;
  wire [0:0] vin0_consume_en_18848;
  wire [0:0] vout_canPeek_18848;
  wire [7:0] vout_peek_18848;
  wire [0:0] v_18849;
  wire [0:0] v_18850;
  function [0:0] mux_18850(input [0:0] sel);
    case (sel) 0: mux_18850 = 1'h0; 1: mux_18850 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18851;
  wire [0:0] v_18852;
  wire [0:0] v_18853;
  wire [0:0] v_18854;
  wire [0:0] v_18855;
  function [0:0] mux_18855(input [0:0] sel);
    case (sel) 0: mux_18855 = 1'h0; 1: mux_18855 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18856;
  wire [0:0] vin0_consume_en_18857;
  wire [0:0] vout_canPeek_18857;
  wire [7:0] vout_peek_18857;
  wire [0:0] v_18858;
  wire [0:0] v_18859;
  function [0:0] mux_18859(input [0:0] sel);
    case (sel) 0: mux_18859 = 1'h0; 1: mux_18859 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18860;
  function [0:0] mux_18860(input [0:0] sel);
    case (sel) 0: mux_18860 = 1'h0; 1: mux_18860 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18861;
  wire [0:0] v_18862;
  wire [0:0] v_18863;
  wire [0:0] v_18864;
  wire [0:0] v_18865;
  wire [0:0] v_18866;
  wire [0:0] v_18867;
  function [0:0] mux_18867(input [0:0] sel);
    case (sel) 0: mux_18867 = 1'h0; 1: mux_18867 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18868;
  wire [0:0] v_18869;
  wire [0:0] v_18870;
  wire [0:0] v_18871;
  wire [0:0] v_18872;
  function [0:0] mux_18872(input [0:0] sel);
    case (sel) 0: mux_18872 = 1'h0; 1: mux_18872 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18873;
  wire [0:0] v_18874;
  wire [0:0] v_18875;
  wire [0:0] v_18876;
  function [0:0] mux_18876(input [0:0] sel);
    case (sel) 0: mux_18876 = 1'h0; 1: mux_18876 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18877;
  function [0:0] mux_18877(input [0:0] sel);
    case (sel) 0: mux_18877 = 1'h0; 1: mux_18877 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_18878 = 1'h0;
  wire [0:0] v_18879;
  wire [0:0] v_18880;
  wire [0:0] act_18881;
  wire [0:0] v_18882;
  wire [0:0] v_18883;
  wire [0:0] v_18884;
  wire [0:0] vin0_consume_en_18885;
  wire [0:0] vout_canPeek_18885;
  wire [7:0] vout_peek_18885;
  wire [0:0] v_18886;
  wire [0:0] v_18887;
  function [0:0] mux_18887(input [0:0] sel);
    case (sel) 0: mux_18887 = 1'h0; 1: mux_18887 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18888;
  wire [0:0] v_18889;
  wire [0:0] v_18890;
  wire [0:0] v_18891;
  wire [0:0] v_18892;
  function [0:0] mux_18892(input [0:0] sel);
    case (sel) 0: mux_18892 = 1'h0; 1: mux_18892 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18893;
  wire [0:0] vin0_consume_en_18894;
  wire [0:0] vout_canPeek_18894;
  wire [7:0] vout_peek_18894;
  wire [0:0] v_18895;
  wire [0:0] v_18896;
  function [0:0] mux_18896(input [0:0] sel);
    case (sel) 0: mux_18896 = 1'h0; 1: mux_18896 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18897;
  function [0:0] mux_18897(input [0:0] sel);
    case (sel) 0: mux_18897 = 1'h0; 1: mux_18897 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18898;
  wire [0:0] v_18899;
  wire [0:0] v_18900;
  wire [0:0] v_18901;
  wire [0:0] v_18902;
  wire [0:0] v_18903;
  wire [0:0] v_18904;
  function [0:0] mux_18904(input [0:0] sel);
    case (sel) 0: mux_18904 = 1'h0; 1: mux_18904 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18905;
  function [0:0] mux_18905(input [0:0] sel);
    case (sel) 0: mux_18905 = 1'h0; 1: mux_18905 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18906;
  wire [0:0] v_18907;
  wire [0:0] v_18908;
  wire [0:0] v_18909;
  function [0:0] mux_18909(input [0:0] sel);
    case (sel) 0: mux_18909 = 1'h0; 1: mux_18909 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18910;
  function [0:0] mux_18910(input [0:0] sel);
    case (sel) 0: mux_18910 = 1'h0; 1: mux_18910 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18911;
  wire [0:0] v_18912;
  wire [0:0] v_18913;
  wire [0:0] v_18914;
  wire [0:0] v_18915;
  wire [0:0] v_18916;
  function [0:0] mux_18916(input [0:0] sel);
    case (sel) 0: mux_18916 = 1'h0; 1: mux_18916 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18917;
  function [0:0] mux_18917(input [0:0] sel);
    case (sel) 0: mux_18917 = 1'h0; 1: mux_18917 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18918;
  wire [0:0] v_18919;
  wire [0:0] v_18920;
  wire [0:0] v_18921;
  function [0:0] mux_18921(input [0:0] sel);
    case (sel) 0: mux_18921 = 1'h0; 1: mux_18921 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18922;
  function [0:0] mux_18922(input [0:0] sel);
    case (sel) 0: mux_18922 = 1'h0; 1: mux_18922 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18923;
  wire [0:0] v_18924;
  wire [0:0] v_18925;
  wire [0:0] v_18926;
  wire [0:0] v_18927;
  wire [0:0] v_18928;
  function [0:0] mux_18928(input [0:0] sel);
    case (sel) 0: mux_18928 = 1'h0; 1: mux_18928 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18929;
  wire [0:0] v_18930;
  wire [0:0] v_18931;
  wire [0:0] v_18932;
  wire [0:0] v_18933;
  function [0:0] mux_18933(input [0:0] sel);
    case (sel) 0: mux_18933 = 1'h0; 1: mux_18933 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18934;
  wire [0:0] v_18935;
  wire [0:0] v_18936;
  wire [0:0] v_18937;
  function [0:0] mux_18937(input [0:0] sel);
    case (sel) 0: mux_18937 = 1'h0; 1: mux_18937 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18938;
  function [0:0] mux_18938(input [0:0] sel);
    case (sel) 0: mux_18938 = 1'h0; 1: mux_18938 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_18939 = 1'h0;
  wire [0:0] v_18940;
  wire [0:0] v_18941;
  wire [0:0] act_18942;
  wire [0:0] v_18943;
  wire [0:0] v_18944;
  wire [0:0] v_18945;
  reg [0:0] v_18946 = 1'h0;
  wire [0:0] v_18947;
  wire [0:0] v_18948;
  wire [0:0] act_18949;
  wire [0:0] v_18950;
  wire [0:0] v_18951;
  wire [0:0] v_18952;
  reg [0:0] v_18953 = 1'h0;
  wire [0:0] v_18954;
  wire [0:0] v_18955;
  wire [0:0] act_18956;
  wire [0:0] v_18957;
  wire [0:0] v_18958;
  wire [0:0] v_18959;
  wire [0:0] vin0_consume_en_18960;
  wire [0:0] vout_canPeek_18960;
  wire [7:0] vout_peek_18960;
  wire [0:0] v_18961;
  wire [0:0] v_18962;
  function [0:0] mux_18962(input [0:0] sel);
    case (sel) 0: mux_18962 = 1'h0; 1: mux_18962 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18963;
  wire [0:0] v_18964;
  wire [0:0] v_18965;
  wire [0:0] v_18966;
  wire [0:0] v_18967;
  function [0:0] mux_18967(input [0:0] sel);
    case (sel) 0: mux_18967 = 1'h0; 1: mux_18967 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18968;
  wire [0:0] vin0_consume_en_18969;
  wire [0:0] vout_canPeek_18969;
  wire [7:0] vout_peek_18969;
  wire [0:0] v_18970;
  wire [0:0] v_18971;
  function [0:0] mux_18971(input [0:0] sel);
    case (sel) 0: mux_18971 = 1'h0; 1: mux_18971 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18972;
  function [0:0] mux_18972(input [0:0] sel);
    case (sel) 0: mux_18972 = 1'h0; 1: mux_18972 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18973;
  wire [0:0] v_18974;
  wire [0:0] v_18975;
  wire [0:0] v_18976;
  wire [0:0] v_18977;
  wire [0:0] v_18978;
  wire [0:0] v_18979;
  function [0:0] mux_18979(input [0:0] sel);
    case (sel) 0: mux_18979 = 1'h0; 1: mux_18979 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18980;
  wire [0:0] v_18981;
  wire [0:0] v_18982;
  wire [0:0] v_18983;
  wire [0:0] v_18984;
  function [0:0] mux_18984(input [0:0] sel);
    case (sel) 0: mux_18984 = 1'h0; 1: mux_18984 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_18985;
  wire [0:0] v_18986;
  wire [0:0] v_18987;
  wire [0:0] v_18988;
  function [0:0] mux_18988(input [0:0] sel);
    case (sel) 0: mux_18988 = 1'h0; 1: mux_18988 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_18989;
  function [0:0] mux_18989(input [0:0] sel);
    case (sel) 0: mux_18989 = 1'h0; 1: mux_18989 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_18990 = 1'h0;
  wire [0:0] v_18991;
  wire [0:0] v_18992;
  wire [0:0] act_18993;
  wire [0:0] v_18994;
  wire [0:0] v_18995;
  wire [0:0] v_18996;
  wire [0:0] vin0_consume_en_18997;
  wire [0:0] vout_canPeek_18997;
  wire [7:0] vout_peek_18997;
  wire [0:0] v_18998;
  wire [0:0] v_18999;
  function [0:0] mux_18999(input [0:0] sel);
    case (sel) 0: mux_18999 = 1'h0; 1: mux_18999 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19000;
  wire [0:0] v_19001;
  wire [0:0] v_19002;
  wire [0:0] v_19003;
  wire [0:0] v_19004;
  function [0:0] mux_19004(input [0:0] sel);
    case (sel) 0: mux_19004 = 1'h0; 1: mux_19004 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19005;
  wire [0:0] vin0_consume_en_19006;
  wire [0:0] vout_canPeek_19006;
  wire [7:0] vout_peek_19006;
  wire [0:0] v_19007;
  wire [0:0] v_19008;
  function [0:0] mux_19008(input [0:0] sel);
    case (sel) 0: mux_19008 = 1'h0; 1: mux_19008 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19009;
  function [0:0] mux_19009(input [0:0] sel);
    case (sel) 0: mux_19009 = 1'h0; 1: mux_19009 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19010;
  wire [0:0] v_19011;
  wire [0:0] v_19012;
  wire [0:0] v_19013;
  wire [0:0] v_19014;
  wire [0:0] v_19015;
  wire [0:0] v_19016;
  function [0:0] mux_19016(input [0:0] sel);
    case (sel) 0: mux_19016 = 1'h0; 1: mux_19016 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19017;
  function [0:0] mux_19017(input [0:0] sel);
    case (sel) 0: mux_19017 = 1'h0; 1: mux_19017 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19018;
  wire [0:0] v_19019;
  wire [0:0] v_19020;
  wire [0:0] v_19021;
  function [0:0] mux_19021(input [0:0] sel);
    case (sel) 0: mux_19021 = 1'h0; 1: mux_19021 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19022;
  function [0:0] mux_19022(input [0:0] sel);
    case (sel) 0: mux_19022 = 1'h0; 1: mux_19022 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19023;
  wire [0:0] v_19024;
  wire [0:0] v_19025;
  wire [0:0] v_19026;
  wire [0:0] v_19027;
  wire [0:0] v_19028;
  function [0:0] mux_19028(input [0:0] sel);
    case (sel) 0: mux_19028 = 1'h0; 1: mux_19028 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19029;
  wire [0:0] v_19030;
  wire [0:0] v_19031;
  wire [0:0] v_19032;
  wire [0:0] v_19033;
  function [0:0] mux_19033(input [0:0] sel);
    case (sel) 0: mux_19033 = 1'h0; 1: mux_19033 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19034;
  wire [0:0] v_19035;
  wire [0:0] v_19036;
  wire [0:0] v_19037;
  function [0:0] mux_19037(input [0:0] sel);
    case (sel) 0: mux_19037 = 1'h0; 1: mux_19037 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19038;
  function [0:0] mux_19038(input [0:0] sel);
    case (sel) 0: mux_19038 = 1'h0; 1: mux_19038 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_19039 = 1'h0;
  wire [0:0] v_19040;
  wire [0:0] v_19041;
  wire [0:0] act_19042;
  wire [0:0] v_19043;
  wire [0:0] v_19044;
  wire [0:0] v_19045;
  reg [0:0] v_19046 = 1'h0;
  wire [0:0] v_19047;
  wire [0:0] v_19048;
  wire [0:0] act_19049;
  wire [0:0] v_19050;
  wire [0:0] v_19051;
  wire [0:0] v_19052;
  wire [0:0] vin0_consume_en_19053;
  wire [0:0] vout_canPeek_19053;
  wire [7:0] vout_peek_19053;
  wire [0:0] v_19054;
  wire [0:0] v_19055;
  function [0:0] mux_19055(input [0:0] sel);
    case (sel) 0: mux_19055 = 1'h0; 1: mux_19055 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19056;
  wire [0:0] v_19057;
  wire [0:0] v_19058;
  wire [0:0] v_19059;
  wire [0:0] v_19060;
  function [0:0] mux_19060(input [0:0] sel);
    case (sel) 0: mux_19060 = 1'h0; 1: mux_19060 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19061;
  wire [0:0] vin0_consume_en_19062;
  wire [0:0] vout_canPeek_19062;
  wire [7:0] vout_peek_19062;
  wire [0:0] v_19063;
  wire [0:0] v_19064;
  function [0:0] mux_19064(input [0:0] sel);
    case (sel) 0: mux_19064 = 1'h0; 1: mux_19064 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19065;
  function [0:0] mux_19065(input [0:0] sel);
    case (sel) 0: mux_19065 = 1'h0; 1: mux_19065 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19066;
  wire [0:0] v_19067;
  wire [0:0] v_19068;
  wire [0:0] v_19069;
  wire [0:0] v_19070;
  wire [0:0] v_19071;
  wire [0:0] v_19072;
  function [0:0] mux_19072(input [0:0] sel);
    case (sel) 0: mux_19072 = 1'h0; 1: mux_19072 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19073;
  wire [0:0] v_19074;
  wire [0:0] v_19075;
  wire [0:0] v_19076;
  wire [0:0] v_19077;
  function [0:0] mux_19077(input [0:0] sel);
    case (sel) 0: mux_19077 = 1'h0; 1: mux_19077 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19078;
  wire [0:0] v_19079;
  wire [0:0] v_19080;
  wire [0:0] v_19081;
  function [0:0] mux_19081(input [0:0] sel);
    case (sel) 0: mux_19081 = 1'h0; 1: mux_19081 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19082;
  function [0:0] mux_19082(input [0:0] sel);
    case (sel) 0: mux_19082 = 1'h0; 1: mux_19082 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_19083 = 1'h0;
  wire [0:0] v_19084;
  wire [0:0] v_19085;
  wire [0:0] act_19086;
  wire [0:0] v_19087;
  wire [0:0] v_19088;
  wire [0:0] v_19089;
  wire [0:0] vin0_consume_en_19090;
  wire [0:0] vout_canPeek_19090;
  wire [7:0] vout_peek_19090;
  wire [0:0] v_19091;
  wire [0:0] v_19092;
  function [0:0] mux_19092(input [0:0] sel);
    case (sel) 0: mux_19092 = 1'h0; 1: mux_19092 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19093;
  wire [0:0] v_19094;
  wire [0:0] v_19095;
  wire [0:0] v_19096;
  wire [0:0] v_19097;
  function [0:0] mux_19097(input [0:0] sel);
    case (sel) 0: mux_19097 = 1'h0; 1: mux_19097 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19098;
  wire [0:0] vin0_consume_en_19099;
  wire [0:0] vout_canPeek_19099;
  wire [7:0] vout_peek_19099;
  wire [0:0] v_19100;
  wire [0:0] v_19101;
  function [0:0] mux_19101(input [0:0] sel);
    case (sel) 0: mux_19101 = 1'h0; 1: mux_19101 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19102;
  function [0:0] mux_19102(input [0:0] sel);
    case (sel) 0: mux_19102 = 1'h0; 1: mux_19102 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19103;
  wire [0:0] v_19104;
  wire [0:0] v_19105;
  wire [0:0] v_19106;
  wire [0:0] v_19107;
  wire [0:0] v_19108;
  wire [0:0] v_19109;
  function [0:0] mux_19109(input [0:0] sel);
    case (sel) 0: mux_19109 = 1'h0; 1: mux_19109 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19110;
  function [0:0] mux_19110(input [0:0] sel);
    case (sel) 0: mux_19110 = 1'h0; 1: mux_19110 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19111;
  wire [0:0] v_19112;
  wire [0:0] v_19113;
  wire [0:0] v_19114;
  function [0:0] mux_19114(input [0:0] sel);
    case (sel) 0: mux_19114 = 1'h0; 1: mux_19114 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19115;
  function [0:0] mux_19115(input [0:0] sel);
    case (sel) 0: mux_19115 = 1'h0; 1: mux_19115 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19116;
  wire [0:0] v_19117;
  wire [0:0] v_19118;
  wire [0:0] v_19119;
  wire [0:0] v_19120;
  wire [0:0] v_19121;
  function [0:0] mux_19121(input [0:0] sel);
    case (sel) 0: mux_19121 = 1'h0; 1: mux_19121 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19122;
  function [0:0] mux_19122(input [0:0] sel);
    case (sel) 0: mux_19122 = 1'h0; 1: mux_19122 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19123;
  wire [0:0] v_19124;
  wire [0:0] v_19125;
  wire [0:0] v_19126;
  function [0:0] mux_19126(input [0:0] sel);
    case (sel) 0: mux_19126 = 1'h0; 1: mux_19126 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19127;
  function [0:0] mux_19127(input [0:0] sel);
    case (sel) 0: mux_19127 = 1'h0; 1: mux_19127 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19128;
  wire [0:0] v_19129;
  wire [0:0] v_19130;
  wire [0:0] v_19131;
  wire [0:0] v_19132;
  wire [0:0] v_19133;
  function [0:0] mux_19133(input [0:0] sel);
    case (sel) 0: mux_19133 = 1'h0; 1: mux_19133 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19134;
  function [0:0] mux_19134(input [0:0] sel);
    case (sel) 0: mux_19134 = 1'h0; 1: mux_19134 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19135;
  wire [0:0] v_19136;
  wire [0:0] v_19137;
  wire [0:0] v_19138;
  function [0:0] mux_19138(input [0:0] sel);
    case (sel) 0: mux_19138 = 1'h0; 1: mux_19138 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19139;
  function [0:0] mux_19139(input [0:0] sel);
    case (sel) 0: mux_19139 = 1'h0; 1: mux_19139 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19140;
  wire [0:0] v_19141;
  wire [0:0] v_19142;
  wire [0:0] v_19143;
  wire [0:0] v_19144;
  wire [0:0] v_19145;
  function [0:0] mux_19145(input [0:0] sel);
    case (sel) 0: mux_19145 = 1'h0; 1: mux_19145 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19146;
  wire [0:0] v_19147;
  wire [0:0] v_19148;
  wire [0:0] v_19149;
  wire [0:0] v_19150;
  function [0:0] mux_19150(input [0:0] sel);
    case (sel) 0: mux_19150 = 1'h0; 1: mux_19150 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19151;
  wire [0:0] v_19152;
  wire [0:0] v_19153;
  wire [0:0] v_19154;
  function [0:0] mux_19154(input [0:0] sel);
    case (sel) 0: mux_19154 = 1'h0; 1: mux_19154 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19155;
  function [0:0] mux_19155(input [0:0] sel);
    case (sel) 0: mux_19155 = 1'h0; 1: mux_19155 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_19156 = 1'h0;
  wire [0:0] v_19157;
  wire [0:0] v_19158;
  wire [0:0] act_19159;
  wire [0:0] v_19160;
  wire [0:0] v_19161;
  wire [0:0] v_19162;
  reg [0:0] v_19163 = 1'h0;
  wire [0:0] v_19164;
  wire [0:0] v_19165;
  wire [0:0] act_19166;
  wire [0:0] v_19167;
  wire [0:0] v_19168;
  wire [0:0] v_19169;
  reg [0:0] v_19170 = 1'h0;
  wire [0:0] v_19171;
  wire [0:0] v_19172;
  wire [0:0] act_19173;
  wire [0:0] v_19174;
  wire [0:0] v_19175;
  wire [0:0] v_19176;
  reg [0:0] v_19177 = 1'h0;
  wire [0:0] v_19178;
  wire [0:0] v_19179;
  wire [0:0] act_19180;
  wire [0:0] v_19181;
  wire [0:0] v_19182;
  wire [0:0] v_19183;
  wire [0:0] vin0_consume_en_19184;
  wire [0:0] vout_canPeek_19184;
  wire [7:0] vout_peek_19184;
  wire [0:0] v_19185;
  wire [0:0] v_19186;
  function [0:0] mux_19186(input [0:0] sel);
    case (sel) 0: mux_19186 = 1'h0; 1: mux_19186 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19187;
  wire [0:0] v_19188;
  wire [0:0] v_19189;
  wire [0:0] v_19190;
  wire [0:0] v_19191;
  function [0:0] mux_19191(input [0:0] sel);
    case (sel) 0: mux_19191 = 1'h0; 1: mux_19191 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19192;
  wire [0:0] vin0_consume_en_19193;
  wire [0:0] vout_canPeek_19193;
  wire [7:0] vout_peek_19193;
  wire [0:0] v_19194;
  wire [0:0] v_19195;
  function [0:0] mux_19195(input [0:0] sel);
    case (sel) 0: mux_19195 = 1'h0; 1: mux_19195 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19196;
  function [0:0] mux_19196(input [0:0] sel);
    case (sel) 0: mux_19196 = 1'h0; 1: mux_19196 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19197;
  wire [0:0] v_19198;
  wire [0:0] v_19199;
  wire [0:0] v_19200;
  wire [0:0] v_19201;
  wire [0:0] v_19202;
  wire [0:0] v_19203;
  function [0:0] mux_19203(input [0:0] sel);
    case (sel) 0: mux_19203 = 1'h0; 1: mux_19203 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19204;
  wire [0:0] v_19205;
  wire [0:0] v_19206;
  wire [0:0] v_19207;
  wire [0:0] v_19208;
  function [0:0] mux_19208(input [0:0] sel);
    case (sel) 0: mux_19208 = 1'h0; 1: mux_19208 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19209;
  wire [0:0] v_19210;
  wire [0:0] v_19211;
  wire [0:0] v_19212;
  function [0:0] mux_19212(input [0:0] sel);
    case (sel) 0: mux_19212 = 1'h0; 1: mux_19212 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19213;
  function [0:0] mux_19213(input [0:0] sel);
    case (sel) 0: mux_19213 = 1'h0; 1: mux_19213 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_19214 = 1'h0;
  wire [0:0] v_19215;
  wire [0:0] v_19216;
  wire [0:0] act_19217;
  wire [0:0] v_19218;
  wire [0:0] v_19219;
  wire [0:0] v_19220;
  wire [0:0] vin0_consume_en_19221;
  wire [0:0] vout_canPeek_19221;
  wire [7:0] vout_peek_19221;
  wire [0:0] v_19222;
  wire [0:0] v_19223;
  function [0:0] mux_19223(input [0:0] sel);
    case (sel) 0: mux_19223 = 1'h0; 1: mux_19223 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19224;
  wire [0:0] v_19225;
  wire [0:0] v_19226;
  wire [0:0] v_19227;
  wire [0:0] v_19228;
  function [0:0] mux_19228(input [0:0] sel);
    case (sel) 0: mux_19228 = 1'h0; 1: mux_19228 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19229;
  wire [0:0] vin0_consume_en_19230;
  wire [0:0] vout_canPeek_19230;
  wire [7:0] vout_peek_19230;
  wire [0:0] v_19231;
  wire [0:0] v_19232;
  function [0:0] mux_19232(input [0:0] sel);
    case (sel) 0: mux_19232 = 1'h0; 1: mux_19232 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19233;
  function [0:0] mux_19233(input [0:0] sel);
    case (sel) 0: mux_19233 = 1'h0; 1: mux_19233 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19234;
  wire [0:0] v_19235;
  wire [0:0] v_19236;
  wire [0:0] v_19237;
  wire [0:0] v_19238;
  wire [0:0] v_19239;
  wire [0:0] v_19240;
  function [0:0] mux_19240(input [0:0] sel);
    case (sel) 0: mux_19240 = 1'h0; 1: mux_19240 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19241;
  function [0:0] mux_19241(input [0:0] sel);
    case (sel) 0: mux_19241 = 1'h0; 1: mux_19241 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19242;
  wire [0:0] v_19243;
  wire [0:0] v_19244;
  wire [0:0] v_19245;
  function [0:0] mux_19245(input [0:0] sel);
    case (sel) 0: mux_19245 = 1'h0; 1: mux_19245 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19246;
  function [0:0] mux_19246(input [0:0] sel);
    case (sel) 0: mux_19246 = 1'h0; 1: mux_19246 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19247;
  wire [0:0] v_19248;
  wire [0:0] v_19249;
  wire [0:0] v_19250;
  wire [0:0] v_19251;
  wire [0:0] v_19252;
  function [0:0] mux_19252(input [0:0] sel);
    case (sel) 0: mux_19252 = 1'h0; 1: mux_19252 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19253;
  wire [0:0] v_19254;
  wire [0:0] v_19255;
  wire [0:0] v_19256;
  wire [0:0] v_19257;
  function [0:0] mux_19257(input [0:0] sel);
    case (sel) 0: mux_19257 = 1'h0; 1: mux_19257 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19258;
  wire [0:0] v_19259;
  wire [0:0] v_19260;
  wire [0:0] v_19261;
  function [0:0] mux_19261(input [0:0] sel);
    case (sel) 0: mux_19261 = 1'h0; 1: mux_19261 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19262;
  function [0:0] mux_19262(input [0:0] sel);
    case (sel) 0: mux_19262 = 1'h0; 1: mux_19262 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_19263 = 1'h0;
  wire [0:0] v_19264;
  wire [0:0] v_19265;
  wire [0:0] act_19266;
  wire [0:0] v_19267;
  wire [0:0] v_19268;
  wire [0:0] v_19269;
  reg [0:0] v_19270 = 1'h0;
  wire [0:0] v_19271;
  wire [0:0] v_19272;
  wire [0:0] act_19273;
  wire [0:0] v_19274;
  wire [0:0] v_19275;
  wire [0:0] v_19276;
  wire [0:0] vin0_consume_en_19277;
  wire [0:0] vout_canPeek_19277;
  wire [7:0] vout_peek_19277;
  wire [0:0] v_19278;
  wire [0:0] v_19279;
  function [0:0] mux_19279(input [0:0] sel);
    case (sel) 0: mux_19279 = 1'h0; 1: mux_19279 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19280;
  wire [0:0] v_19281;
  wire [0:0] v_19282;
  wire [0:0] v_19283;
  wire [0:0] v_19284;
  function [0:0] mux_19284(input [0:0] sel);
    case (sel) 0: mux_19284 = 1'h0; 1: mux_19284 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19285;
  wire [0:0] vin0_consume_en_19286;
  wire [0:0] vout_canPeek_19286;
  wire [7:0] vout_peek_19286;
  wire [0:0] v_19287;
  wire [0:0] v_19288;
  function [0:0] mux_19288(input [0:0] sel);
    case (sel) 0: mux_19288 = 1'h0; 1: mux_19288 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19289;
  function [0:0] mux_19289(input [0:0] sel);
    case (sel) 0: mux_19289 = 1'h0; 1: mux_19289 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19290;
  wire [0:0] v_19291;
  wire [0:0] v_19292;
  wire [0:0] v_19293;
  wire [0:0] v_19294;
  wire [0:0] v_19295;
  wire [0:0] v_19296;
  function [0:0] mux_19296(input [0:0] sel);
    case (sel) 0: mux_19296 = 1'h0; 1: mux_19296 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19297;
  wire [0:0] v_19298;
  wire [0:0] v_19299;
  wire [0:0] v_19300;
  wire [0:0] v_19301;
  function [0:0] mux_19301(input [0:0] sel);
    case (sel) 0: mux_19301 = 1'h0; 1: mux_19301 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19302;
  wire [0:0] v_19303;
  wire [0:0] v_19304;
  wire [0:0] v_19305;
  function [0:0] mux_19305(input [0:0] sel);
    case (sel) 0: mux_19305 = 1'h0; 1: mux_19305 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19306;
  function [0:0] mux_19306(input [0:0] sel);
    case (sel) 0: mux_19306 = 1'h0; 1: mux_19306 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_19307 = 1'h0;
  wire [0:0] v_19308;
  wire [0:0] v_19309;
  wire [0:0] act_19310;
  wire [0:0] v_19311;
  wire [0:0] v_19312;
  wire [0:0] v_19313;
  wire [0:0] vin0_consume_en_19314;
  wire [0:0] vout_canPeek_19314;
  wire [7:0] vout_peek_19314;
  wire [0:0] v_19315;
  wire [0:0] v_19316;
  function [0:0] mux_19316(input [0:0] sel);
    case (sel) 0: mux_19316 = 1'h0; 1: mux_19316 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19317;
  wire [0:0] v_19318;
  wire [0:0] v_19319;
  wire [0:0] v_19320;
  wire [0:0] v_19321;
  function [0:0] mux_19321(input [0:0] sel);
    case (sel) 0: mux_19321 = 1'h0; 1: mux_19321 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19322;
  wire [0:0] vin0_consume_en_19323;
  wire [0:0] vout_canPeek_19323;
  wire [7:0] vout_peek_19323;
  wire [0:0] v_19324;
  wire [0:0] v_19325;
  function [0:0] mux_19325(input [0:0] sel);
    case (sel) 0: mux_19325 = 1'h0; 1: mux_19325 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19326;
  function [0:0] mux_19326(input [0:0] sel);
    case (sel) 0: mux_19326 = 1'h0; 1: mux_19326 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19327;
  wire [0:0] v_19328;
  wire [0:0] v_19329;
  wire [0:0] v_19330;
  wire [0:0] v_19331;
  wire [0:0] v_19332;
  wire [0:0] v_19333;
  function [0:0] mux_19333(input [0:0] sel);
    case (sel) 0: mux_19333 = 1'h0; 1: mux_19333 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19334;
  function [0:0] mux_19334(input [0:0] sel);
    case (sel) 0: mux_19334 = 1'h0; 1: mux_19334 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19335;
  wire [0:0] v_19336;
  wire [0:0] v_19337;
  wire [0:0] v_19338;
  function [0:0] mux_19338(input [0:0] sel);
    case (sel) 0: mux_19338 = 1'h0; 1: mux_19338 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19339;
  function [0:0] mux_19339(input [0:0] sel);
    case (sel) 0: mux_19339 = 1'h0; 1: mux_19339 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19340;
  wire [0:0] v_19341;
  wire [0:0] v_19342;
  wire [0:0] v_19343;
  wire [0:0] v_19344;
  wire [0:0] v_19345;
  function [0:0] mux_19345(input [0:0] sel);
    case (sel) 0: mux_19345 = 1'h0; 1: mux_19345 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19346;
  function [0:0] mux_19346(input [0:0] sel);
    case (sel) 0: mux_19346 = 1'h0; 1: mux_19346 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19347;
  wire [0:0] v_19348;
  wire [0:0] v_19349;
  wire [0:0] v_19350;
  function [0:0] mux_19350(input [0:0] sel);
    case (sel) 0: mux_19350 = 1'h0; 1: mux_19350 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19351;
  function [0:0] mux_19351(input [0:0] sel);
    case (sel) 0: mux_19351 = 1'h0; 1: mux_19351 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19352;
  wire [0:0] v_19353;
  wire [0:0] v_19354;
  wire [0:0] v_19355;
  wire [0:0] v_19356;
  wire [0:0] v_19357;
  function [0:0] mux_19357(input [0:0] sel);
    case (sel) 0: mux_19357 = 1'h0; 1: mux_19357 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19358;
  wire [0:0] v_19359;
  wire [0:0] v_19360;
  wire [0:0] v_19361;
  wire [0:0] v_19362;
  function [0:0] mux_19362(input [0:0] sel);
    case (sel) 0: mux_19362 = 1'h0; 1: mux_19362 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19363;
  wire [0:0] v_19364;
  wire [0:0] v_19365;
  wire [0:0] v_19366;
  function [0:0] mux_19366(input [0:0] sel);
    case (sel) 0: mux_19366 = 1'h0; 1: mux_19366 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19367;
  function [0:0] mux_19367(input [0:0] sel);
    case (sel) 0: mux_19367 = 1'h0; 1: mux_19367 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_19368 = 1'h0;
  wire [0:0] v_19369;
  wire [0:0] v_19370;
  wire [0:0] act_19371;
  wire [0:0] v_19372;
  wire [0:0] v_19373;
  wire [0:0] v_19374;
  reg [0:0] v_19375 = 1'h0;
  wire [0:0] v_19376;
  wire [0:0] v_19377;
  wire [0:0] act_19378;
  wire [0:0] v_19379;
  wire [0:0] v_19380;
  wire [0:0] v_19381;
  reg [0:0] v_19382 = 1'h0;
  wire [0:0] v_19383;
  wire [0:0] v_19384;
  wire [0:0] act_19385;
  wire [0:0] v_19386;
  wire [0:0] v_19387;
  wire [0:0] v_19388;
  wire [0:0] vin0_consume_en_19389;
  wire [0:0] vout_canPeek_19389;
  wire [7:0] vout_peek_19389;
  wire [0:0] v_19390;
  wire [0:0] v_19391;
  function [0:0] mux_19391(input [0:0] sel);
    case (sel) 0: mux_19391 = 1'h0; 1: mux_19391 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19392;
  wire [0:0] v_19393;
  wire [0:0] v_19394;
  wire [0:0] v_19395;
  wire [0:0] v_19396;
  function [0:0] mux_19396(input [0:0] sel);
    case (sel) 0: mux_19396 = 1'h0; 1: mux_19396 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19397;
  wire [0:0] vin0_consume_en_19398;
  wire [0:0] vout_canPeek_19398;
  wire [7:0] vout_peek_19398;
  wire [0:0] v_19399;
  wire [0:0] v_19400;
  function [0:0] mux_19400(input [0:0] sel);
    case (sel) 0: mux_19400 = 1'h0; 1: mux_19400 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19401;
  function [0:0] mux_19401(input [0:0] sel);
    case (sel) 0: mux_19401 = 1'h0; 1: mux_19401 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19402;
  wire [0:0] v_19403;
  wire [0:0] v_19404;
  wire [0:0] v_19405;
  wire [0:0] v_19406;
  wire [0:0] v_19407;
  wire [0:0] v_19408;
  function [0:0] mux_19408(input [0:0] sel);
    case (sel) 0: mux_19408 = 1'h0; 1: mux_19408 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19409;
  wire [0:0] v_19410;
  wire [0:0] v_19411;
  wire [0:0] v_19412;
  wire [0:0] v_19413;
  function [0:0] mux_19413(input [0:0] sel);
    case (sel) 0: mux_19413 = 1'h0; 1: mux_19413 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19414;
  wire [0:0] v_19415;
  wire [0:0] v_19416;
  wire [0:0] v_19417;
  function [0:0] mux_19417(input [0:0] sel);
    case (sel) 0: mux_19417 = 1'h0; 1: mux_19417 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19418;
  function [0:0] mux_19418(input [0:0] sel);
    case (sel) 0: mux_19418 = 1'h0; 1: mux_19418 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_19419 = 1'h0;
  wire [0:0] v_19420;
  wire [0:0] v_19421;
  wire [0:0] act_19422;
  wire [0:0] v_19423;
  wire [0:0] v_19424;
  wire [0:0] v_19425;
  wire [0:0] vin0_consume_en_19426;
  wire [0:0] vout_canPeek_19426;
  wire [7:0] vout_peek_19426;
  wire [0:0] v_19427;
  wire [0:0] v_19428;
  function [0:0] mux_19428(input [0:0] sel);
    case (sel) 0: mux_19428 = 1'h0; 1: mux_19428 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19429;
  wire [0:0] v_19430;
  wire [0:0] v_19431;
  wire [0:0] v_19432;
  wire [0:0] v_19433;
  function [0:0] mux_19433(input [0:0] sel);
    case (sel) 0: mux_19433 = 1'h0; 1: mux_19433 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19434;
  wire [0:0] vin0_consume_en_19435;
  wire [0:0] vout_canPeek_19435;
  wire [7:0] vout_peek_19435;
  wire [0:0] v_19436;
  wire [0:0] v_19437;
  function [0:0] mux_19437(input [0:0] sel);
    case (sel) 0: mux_19437 = 1'h0; 1: mux_19437 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19438;
  function [0:0] mux_19438(input [0:0] sel);
    case (sel) 0: mux_19438 = 1'h0; 1: mux_19438 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19439;
  wire [0:0] v_19440;
  wire [0:0] v_19441;
  wire [0:0] v_19442;
  wire [0:0] v_19443;
  wire [0:0] v_19444;
  wire [0:0] v_19445;
  function [0:0] mux_19445(input [0:0] sel);
    case (sel) 0: mux_19445 = 1'h0; 1: mux_19445 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19446;
  function [0:0] mux_19446(input [0:0] sel);
    case (sel) 0: mux_19446 = 1'h0; 1: mux_19446 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19447;
  wire [0:0] v_19448;
  wire [0:0] v_19449;
  wire [0:0] v_19450;
  function [0:0] mux_19450(input [0:0] sel);
    case (sel) 0: mux_19450 = 1'h0; 1: mux_19450 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19451;
  function [0:0] mux_19451(input [0:0] sel);
    case (sel) 0: mux_19451 = 1'h0; 1: mux_19451 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19452;
  wire [0:0] v_19453;
  wire [0:0] v_19454;
  wire [0:0] v_19455;
  wire [0:0] v_19456;
  wire [0:0] v_19457;
  function [0:0] mux_19457(input [0:0] sel);
    case (sel) 0: mux_19457 = 1'h0; 1: mux_19457 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19458;
  wire [0:0] v_19459;
  wire [0:0] v_19460;
  wire [0:0] v_19461;
  wire [0:0] v_19462;
  function [0:0] mux_19462(input [0:0] sel);
    case (sel) 0: mux_19462 = 1'h0; 1: mux_19462 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19463;
  wire [0:0] v_19464;
  wire [0:0] v_19465;
  wire [0:0] v_19466;
  function [0:0] mux_19466(input [0:0] sel);
    case (sel) 0: mux_19466 = 1'h0; 1: mux_19466 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19467;
  function [0:0] mux_19467(input [0:0] sel);
    case (sel) 0: mux_19467 = 1'h0; 1: mux_19467 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_19468 = 1'h0;
  wire [0:0] v_19469;
  wire [0:0] v_19470;
  wire [0:0] act_19471;
  wire [0:0] v_19472;
  wire [0:0] v_19473;
  wire [0:0] v_19474;
  reg [0:0] v_19475 = 1'h0;
  wire [0:0] v_19476;
  wire [0:0] v_19477;
  wire [0:0] act_19478;
  wire [0:0] v_19479;
  wire [0:0] v_19480;
  wire [0:0] v_19481;
  wire [0:0] vin0_consume_en_19482;
  wire [0:0] vout_canPeek_19482;
  wire [7:0] vout_peek_19482;
  wire [0:0] v_19483;
  wire [0:0] v_19484;
  function [0:0] mux_19484(input [0:0] sel);
    case (sel) 0: mux_19484 = 1'h0; 1: mux_19484 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19485;
  wire [0:0] v_19486;
  wire [0:0] v_19487;
  wire [0:0] v_19488;
  wire [0:0] v_19489;
  function [0:0] mux_19489(input [0:0] sel);
    case (sel) 0: mux_19489 = 1'h0; 1: mux_19489 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19490;
  wire [0:0] vin0_consume_en_19491;
  wire [0:0] vout_canPeek_19491;
  wire [7:0] vout_peek_19491;
  wire [0:0] v_19492;
  wire [0:0] v_19493;
  function [0:0] mux_19493(input [0:0] sel);
    case (sel) 0: mux_19493 = 1'h0; 1: mux_19493 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19494;
  function [0:0] mux_19494(input [0:0] sel);
    case (sel) 0: mux_19494 = 1'h0; 1: mux_19494 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19495;
  wire [0:0] v_19496;
  wire [0:0] v_19497;
  wire [0:0] v_19498;
  wire [0:0] v_19499;
  wire [0:0] v_19500;
  wire [0:0] v_19501;
  function [0:0] mux_19501(input [0:0] sel);
    case (sel) 0: mux_19501 = 1'h0; 1: mux_19501 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19502;
  wire [0:0] v_19503;
  wire [0:0] v_19504;
  wire [0:0] v_19505;
  wire [0:0] v_19506;
  function [0:0] mux_19506(input [0:0] sel);
    case (sel) 0: mux_19506 = 1'h0; 1: mux_19506 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19507;
  wire [0:0] v_19508;
  wire [0:0] v_19509;
  wire [0:0] v_19510;
  function [0:0] mux_19510(input [0:0] sel);
    case (sel) 0: mux_19510 = 1'h0; 1: mux_19510 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19511;
  function [0:0] mux_19511(input [0:0] sel);
    case (sel) 0: mux_19511 = 1'h0; 1: mux_19511 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_19512 = 1'h0;
  wire [0:0] v_19513;
  wire [0:0] v_19514;
  wire [0:0] act_19515;
  wire [0:0] v_19516;
  wire [0:0] v_19517;
  wire [0:0] v_19518;
  wire [0:0] vin0_consume_en_19519;
  wire [0:0] vout_canPeek_19519;
  wire [7:0] vout_peek_19519;
  wire [0:0] v_19520;
  wire [0:0] v_19521;
  function [0:0] mux_19521(input [0:0] sel);
    case (sel) 0: mux_19521 = 1'h0; 1: mux_19521 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19522;
  wire [0:0] v_19523;
  wire [0:0] v_19524;
  wire [0:0] v_19525;
  wire [0:0] v_19526;
  function [0:0] mux_19526(input [0:0] sel);
    case (sel) 0: mux_19526 = 1'h0; 1: mux_19526 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19527;
  wire [0:0] vin0_consume_en_19528;
  wire [0:0] vout_canPeek_19528;
  wire [7:0] vout_peek_19528;
  wire [0:0] v_19529;
  wire [0:0] v_19530;
  function [0:0] mux_19530(input [0:0] sel);
    case (sel) 0: mux_19530 = 1'h0; 1: mux_19530 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19531;
  function [0:0] mux_19531(input [0:0] sel);
    case (sel) 0: mux_19531 = 1'h0; 1: mux_19531 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19532;
  wire [0:0] v_19533;
  wire [0:0] v_19534;
  wire [0:0] v_19535;
  wire [0:0] v_19536;
  wire [0:0] v_19537;
  wire [0:0] v_19538;
  function [0:0] mux_19538(input [0:0] sel);
    case (sel) 0: mux_19538 = 1'h0; 1: mux_19538 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19539;
  function [0:0] mux_19539(input [0:0] sel);
    case (sel) 0: mux_19539 = 1'h0; 1: mux_19539 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19540;
  wire [0:0] v_19541;
  wire [0:0] v_19542;
  wire [0:0] v_19543;
  function [0:0] mux_19543(input [0:0] sel);
    case (sel) 0: mux_19543 = 1'h0; 1: mux_19543 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19544;
  function [0:0] mux_19544(input [0:0] sel);
    case (sel) 0: mux_19544 = 1'h0; 1: mux_19544 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19545;
  wire [0:0] v_19546;
  wire [0:0] v_19547;
  wire [0:0] v_19548;
  wire [0:0] v_19549;
  wire [0:0] v_19550;
  function [0:0] mux_19550(input [0:0] sel);
    case (sel) 0: mux_19550 = 1'h0; 1: mux_19550 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19551;
  function [0:0] mux_19551(input [0:0] sel);
    case (sel) 0: mux_19551 = 1'h0; 1: mux_19551 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19552;
  wire [0:0] v_19553;
  wire [0:0] v_19554;
  wire [0:0] v_19555;
  function [0:0] mux_19555(input [0:0] sel);
    case (sel) 0: mux_19555 = 1'h0; 1: mux_19555 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19556;
  function [0:0] mux_19556(input [0:0] sel);
    case (sel) 0: mux_19556 = 1'h0; 1: mux_19556 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19557;
  wire [0:0] v_19558;
  wire [0:0] v_19559;
  wire [0:0] v_19560;
  wire [0:0] v_19561;
  wire [0:0] v_19562;
  function [0:0] mux_19562(input [0:0] sel);
    case (sel) 0: mux_19562 = 1'h0; 1: mux_19562 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19563;
  function [0:0] mux_19563(input [0:0] sel);
    case (sel) 0: mux_19563 = 1'h0; 1: mux_19563 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19564;
  wire [0:0] v_19565;
  wire [0:0] v_19566;
  wire [0:0] v_19567;
  function [0:0] mux_19567(input [0:0] sel);
    case (sel) 0: mux_19567 = 1'h0; 1: mux_19567 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19568;
  function [0:0] mux_19568(input [0:0] sel);
    case (sel) 0: mux_19568 = 1'h0; 1: mux_19568 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19569;
  wire [0:0] v_19570;
  wire [0:0] v_19571;
  wire [0:0] v_19572;
  wire [0:0] v_19573;
  wire [0:0] v_19574;
  function [0:0] mux_19574(input [0:0] sel);
    case (sel) 0: mux_19574 = 1'h0; 1: mux_19574 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19575;
  function [0:0] mux_19575(input [0:0] sel);
    case (sel) 0: mux_19575 = 1'h0; 1: mux_19575 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19576;
  wire [0:0] v_19577;
  wire [0:0] v_19578;
  wire [0:0] v_19579;
  function [0:0] mux_19579(input [0:0] sel);
    case (sel) 0: mux_19579 = 1'h0; 1: mux_19579 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19580;
  function [0:0] mux_19580(input [0:0] sel);
    case (sel) 0: mux_19580 = 1'h0; 1: mux_19580 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19581;
  wire [0:0] v_19582;
  wire [0:0] v_19583;
  wire [0:0] v_19584;
  wire [0:0] v_19585;
  wire [0:0] v_19586;
  function [0:0] mux_19586(input [0:0] sel);
    case (sel) 0: mux_19586 = 1'h0; 1: mux_19586 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19587;
  wire [0:0] v_19588;
  wire [0:0] v_19589;
  wire [0:0] v_19590;
  wire [0:0] v_19591;
  function [0:0] mux_19591(input [0:0] sel);
    case (sel) 0: mux_19591 = 1'h0; 1: mux_19591 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19592;
  wire [0:0] v_19593;
  wire [0:0] v_19594;
  wire [0:0] v_19595;
  function [0:0] mux_19595(input [0:0] sel);
    case (sel) 0: mux_19595 = 1'h0; 1: mux_19595 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19596;
  function [0:0] mux_19596(input [0:0] sel);
    case (sel) 0: mux_19596 = 1'h0; 1: mux_19596 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_19597 = 1'h0;
  wire [0:0] v_19598;
  wire [0:0] v_19599;
  wire [0:0] act_19600;
  wire [0:0] v_19601;
  wire [0:0] v_19602;
  wire [0:0] v_19603;
  reg [0:0] v_19604 = 1'h0;
  wire [0:0] v_19605;
  wire [0:0] v_19606;
  wire [0:0] act_19607;
  wire [0:0] v_19608;
  wire [0:0] v_19609;
  wire [0:0] v_19610;
  reg [0:0] v_19611 = 1'h0;
  wire [0:0] v_19612;
  wire [0:0] v_19613;
  wire [0:0] act_19614;
  wire [0:0] v_19615;
  wire [0:0] v_19616;
  wire [0:0] v_19617;
  reg [0:0] v_19618 = 1'h0;
  wire [0:0] v_19619;
  wire [0:0] v_19620;
  wire [0:0] act_19621;
  wire [0:0] v_19622;
  wire [0:0] v_19623;
  wire [0:0] v_19624;
  reg [0:0] v_19625 = 1'h0;
  wire [0:0] v_19626;
  wire [0:0] v_19627;
  wire [0:0] act_19628;
  wire [0:0] v_19629;
  wire [0:0] v_19630;
  wire [0:0] v_19631;
  wire [0:0] vin0_consume_en_19632;
  wire [0:0] vout_canPeek_19632;
  wire [7:0] vout_peek_19632;
  wire [0:0] v_19633;
  wire [0:0] v_19634;
  function [0:0] mux_19634(input [0:0] sel);
    case (sel) 0: mux_19634 = 1'h0; 1: mux_19634 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19635;
  wire [0:0] v_19636;
  wire [0:0] v_19637;
  wire [0:0] v_19638;
  wire [0:0] v_19639;
  function [0:0] mux_19639(input [0:0] sel);
    case (sel) 0: mux_19639 = 1'h0; 1: mux_19639 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19640;
  wire [0:0] vin0_consume_en_19641;
  wire [0:0] vout_canPeek_19641;
  wire [7:0] vout_peek_19641;
  wire [0:0] v_19642;
  wire [0:0] v_19643;
  function [0:0] mux_19643(input [0:0] sel);
    case (sel) 0: mux_19643 = 1'h0; 1: mux_19643 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19644;
  function [0:0] mux_19644(input [0:0] sel);
    case (sel) 0: mux_19644 = 1'h0; 1: mux_19644 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19645;
  wire [0:0] v_19646;
  wire [0:0] v_19647;
  wire [0:0] v_19648;
  wire [0:0] v_19649;
  wire [0:0] v_19650;
  wire [0:0] v_19651;
  function [0:0] mux_19651(input [0:0] sel);
    case (sel) 0: mux_19651 = 1'h0; 1: mux_19651 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19652;
  wire [0:0] v_19653;
  wire [0:0] v_19654;
  wire [0:0] v_19655;
  wire [0:0] v_19656;
  function [0:0] mux_19656(input [0:0] sel);
    case (sel) 0: mux_19656 = 1'h0; 1: mux_19656 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19657;
  wire [0:0] v_19658;
  wire [0:0] v_19659;
  wire [0:0] v_19660;
  function [0:0] mux_19660(input [0:0] sel);
    case (sel) 0: mux_19660 = 1'h0; 1: mux_19660 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19661;
  function [0:0] mux_19661(input [0:0] sel);
    case (sel) 0: mux_19661 = 1'h0; 1: mux_19661 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_19662 = 1'h0;
  wire [0:0] v_19663;
  wire [0:0] v_19664;
  wire [0:0] act_19665;
  wire [0:0] v_19666;
  wire [0:0] v_19667;
  wire [0:0] v_19668;
  wire [0:0] vin0_consume_en_19669;
  wire [0:0] vout_canPeek_19669;
  wire [7:0] vout_peek_19669;
  wire [0:0] v_19670;
  wire [0:0] v_19671;
  function [0:0] mux_19671(input [0:0] sel);
    case (sel) 0: mux_19671 = 1'h0; 1: mux_19671 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19672;
  wire [0:0] v_19673;
  wire [0:0] v_19674;
  wire [0:0] v_19675;
  wire [0:0] v_19676;
  function [0:0] mux_19676(input [0:0] sel);
    case (sel) 0: mux_19676 = 1'h0; 1: mux_19676 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19677;
  wire [0:0] vin0_consume_en_19678;
  wire [0:0] vout_canPeek_19678;
  wire [7:0] vout_peek_19678;
  wire [0:0] v_19679;
  wire [0:0] v_19680;
  function [0:0] mux_19680(input [0:0] sel);
    case (sel) 0: mux_19680 = 1'h0; 1: mux_19680 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19681;
  function [0:0] mux_19681(input [0:0] sel);
    case (sel) 0: mux_19681 = 1'h0; 1: mux_19681 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19682;
  wire [0:0] v_19683;
  wire [0:0] v_19684;
  wire [0:0] v_19685;
  wire [0:0] v_19686;
  wire [0:0] v_19687;
  wire [0:0] v_19688;
  function [0:0] mux_19688(input [0:0] sel);
    case (sel) 0: mux_19688 = 1'h0; 1: mux_19688 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19689;
  function [0:0] mux_19689(input [0:0] sel);
    case (sel) 0: mux_19689 = 1'h0; 1: mux_19689 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19690;
  wire [0:0] v_19691;
  wire [0:0] v_19692;
  wire [0:0] v_19693;
  function [0:0] mux_19693(input [0:0] sel);
    case (sel) 0: mux_19693 = 1'h0; 1: mux_19693 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19694;
  function [0:0] mux_19694(input [0:0] sel);
    case (sel) 0: mux_19694 = 1'h0; 1: mux_19694 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19695;
  wire [0:0] v_19696;
  wire [0:0] v_19697;
  wire [0:0] v_19698;
  wire [0:0] v_19699;
  wire [0:0] v_19700;
  function [0:0] mux_19700(input [0:0] sel);
    case (sel) 0: mux_19700 = 1'h0; 1: mux_19700 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19701;
  wire [0:0] v_19702;
  wire [0:0] v_19703;
  wire [0:0] v_19704;
  wire [0:0] v_19705;
  function [0:0] mux_19705(input [0:0] sel);
    case (sel) 0: mux_19705 = 1'h0; 1: mux_19705 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19706;
  wire [0:0] v_19707;
  wire [0:0] v_19708;
  wire [0:0] v_19709;
  function [0:0] mux_19709(input [0:0] sel);
    case (sel) 0: mux_19709 = 1'h0; 1: mux_19709 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19710;
  function [0:0] mux_19710(input [0:0] sel);
    case (sel) 0: mux_19710 = 1'h0; 1: mux_19710 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_19711 = 1'h0;
  wire [0:0] v_19712;
  wire [0:0] v_19713;
  wire [0:0] act_19714;
  wire [0:0] v_19715;
  wire [0:0] v_19716;
  wire [0:0] v_19717;
  reg [0:0] v_19718 = 1'h0;
  wire [0:0] v_19719;
  wire [0:0] v_19720;
  wire [0:0] act_19721;
  wire [0:0] v_19722;
  wire [0:0] v_19723;
  wire [0:0] v_19724;
  wire [0:0] vin0_consume_en_19725;
  wire [0:0] vout_canPeek_19725;
  wire [7:0] vout_peek_19725;
  wire [0:0] v_19726;
  wire [0:0] v_19727;
  function [0:0] mux_19727(input [0:0] sel);
    case (sel) 0: mux_19727 = 1'h0; 1: mux_19727 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19728;
  wire [0:0] v_19729;
  wire [0:0] v_19730;
  wire [0:0] v_19731;
  wire [0:0] v_19732;
  function [0:0] mux_19732(input [0:0] sel);
    case (sel) 0: mux_19732 = 1'h0; 1: mux_19732 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19733;
  wire [0:0] vin0_consume_en_19734;
  wire [0:0] vout_canPeek_19734;
  wire [7:0] vout_peek_19734;
  wire [0:0] v_19735;
  wire [0:0] v_19736;
  function [0:0] mux_19736(input [0:0] sel);
    case (sel) 0: mux_19736 = 1'h0; 1: mux_19736 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19737;
  function [0:0] mux_19737(input [0:0] sel);
    case (sel) 0: mux_19737 = 1'h0; 1: mux_19737 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19738;
  wire [0:0] v_19739;
  wire [0:0] v_19740;
  wire [0:0] v_19741;
  wire [0:0] v_19742;
  wire [0:0] v_19743;
  wire [0:0] v_19744;
  function [0:0] mux_19744(input [0:0] sel);
    case (sel) 0: mux_19744 = 1'h0; 1: mux_19744 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19745;
  wire [0:0] v_19746;
  wire [0:0] v_19747;
  wire [0:0] v_19748;
  wire [0:0] v_19749;
  function [0:0] mux_19749(input [0:0] sel);
    case (sel) 0: mux_19749 = 1'h0; 1: mux_19749 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19750;
  wire [0:0] v_19751;
  wire [0:0] v_19752;
  wire [0:0] v_19753;
  function [0:0] mux_19753(input [0:0] sel);
    case (sel) 0: mux_19753 = 1'h0; 1: mux_19753 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19754;
  function [0:0] mux_19754(input [0:0] sel);
    case (sel) 0: mux_19754 = 1'h0; 1: mux_19754 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_19755 = 1'h0;
  wire [0:0] v_19756;
  wire [0:0] v_19757;
  wire [0:0] act_19758;
  wire [0:0] v_19759;
  wire [0:0] v_19760;
  wire [0:0] v_19761;
  wire [0:0] vin0_consume_en_19762;
  wire [0:0] vout_canPeek_19762;
  wire [7:0] vout_peek_19762;
  wire [0:0] v_19763;
  wire [0:0] v_19764;
  function [0:0] mux_19764(input [0:0] sel);
    case (sel) 0: mux_19764 = 1'h0; 1: mux_19764 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19765;
  wire [0:0] v_19766;
  wire [0:0] v_19767;
  wire [0:0] v_19768;
  wire [0:0] v_19769;
  function [0:0] mux_19769(input [0:0] sel);
    case (sel) 0: mux_19769 = 1'h0; 1: mux_19769 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19770;
  wire [0:0] vin0_consume_en_19771;
  wire [0:0] vout_canPeek_19771;
  wire [7:0] vout_peek_19771;
  wire [0:0] v_19772;
  wire [0:0] v_19773;
  function [0:0] mux_19773(input [0:0] sel);
    case (sel) 0: mux_19773 = 1'h0; 1: mux_19773 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19774;
  function [0:0] mux_19774(input [0:0] sel);
    case (sel) 0: mux_19774 = 1'h0; 1: mux_19774 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19775;
  wire [0:0] v_19776;
  wire [0:0] v_19777;
  wire [0:0] v_19778;
  wire [0:0] v_19779;
  wire [0:0] v_19780;
  wire [0:0] v_19781;
  function [0:0] mux_19781(input [0:0] sel);
    case (sel) 0: mux_19781 = 1'h0; 1: mux_19781 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19782;
  function [0:0] mux_19782(input [0:0] sel);
    case (sel) 0: mux_19782 = 1'h0; 1: mux_19782 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19783;
  wire [0:0] v_19784;
  wire [0:0] v_19785;
  wire [0:0] v_19786;
  function [0:0] mux_19786(input [0:0] sel);
    case (sel) 0: mux_19786 = 1'h0; 1: mux_19786 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19787;
  function [0:0] mux_19787(input [0:0] sel);
    case (sel) 0: mux_19787 = 1'h0; 1: mux_19787 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19788;
  wire [0:0] v_19789;
  wire [0:0] v_19790;
  wire [0:0] v_19791;
  wire [0:0] v_19792;
  wire [0:0] v_19793;
  function [0:0] mux_19793(input [0:0] sel);
    case (sel) 0: mux_19793 = 1'h0; 1: mux_19793 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19794;
  function [0:0] mux_19794(input [0:0] sel);
    case (sel) 0: mux_19794 = 1'h0; 1: mux_19794 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19795;
  wire [0:0] v_19796;
  wire [0:0] v_19797;
  wire [0:0] v_19798;
  function [0:0] mux_19798(input [0:0] sel);
    case (sel) 0: mux_19798 = 1'h0; 1: mux_19798 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19799;
  function [0:0] mux_19799(input [0:0] sel);
    case (sel) 0: mux_19799 = 1'h0; 1: mux_19799 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19800;
  wire [0:0] v_19801;
  wire [0:0] v_19802;
  wire [0:0] v_19803;
  wire [0:0] v_19804;
  wire [0:0] v_19805;
  function [0:0] mux_19805(input [0:0] sel);
    case (sel) 0: mux_19805 = 1'h0; 1: mux_19805 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19806;
  wire [0:0] v_19807;
  wire [0:0] v_19808;
  wire [0:0] v_19809;
  wire [0:0] v_19810;
  function [0:0] mux_19810(input [0:0] sel);
    case (sel) 0: mux_19810 = 1'h0; 1: mux_19810 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19811;
  wire [0:0] v_19812;
  wire [0:0] v_19813;
  wire [0:0] v_19814;
  function [0:0] mux_19814(input [0:0] sel);
    case (sel) 0: mux_19814 = 1'h0; 1: mux_19814 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19815;
  function [0:0] mux_19815(input [0:0] sel);
    case (sel) 0: mux_19815 = 1'h0; 1: mux_19815 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_19816 = 1'h0;
  wire [0:0] v_19817;
  wire [0:0] v_19818;
  wire [0:0] act_19819;
  wire [0:0] v_19820;
  wire [0:0] v_19821;
  wire [0:0] v_19822;
  reg [0:0] v_19823 = 1'h0;
  wire [0:0] v_19824;
  wire [0:0] v_19825;
  wire [0:0] act_19826;
  wire [0:0] v_19827;
  wire [0:0] v_19828;
  wire [0:0] v_19829;
  reg [0:0] v_19830 = 1'h0;
  wire [0:0] v_19831;
  wire [0:0] v_19832;
  wire [0:0] act_19833;
  wire [0:0] v_19834;
  wire [0:0] v_19835;
  wire [0:0] v_19836;
  wire [0:0] vin0_consume_en_19837;
  wire [0:0] vout_canPeek_19837;
  wire [7:0] vout_peek_19837;
  wire [0:0] v_19838;
  wire [0:0] v_19839;
  function [0:0] mux_19839(input [0:0] sel);
    case (sel) 0: mux_19839 = 1'h0; 1: mux_19839 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19840;
  wire [0:0] v_19841;
  wire [0:0] v_19842;
  wire [0:0] v_19843;
  wire [0:0] v_19844;
  function [0:0] mux_19844(input [0:0] sel);
    case (sel) 0: mux_19844 = 1'h0; 1: mux_19844 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19845;
  wire [0:0] vin0_consume_en_19846;
  wire [0:0] vout_canPeek_19846;
  wire [7:0] vout_peek_19846;
  wire [0:0] v_19847;
  wire [0:0] v_19848;
  function [0:0] mux_19848(input [0:0] sel);
    case (sel) 0: mux_19848 = 1'h0; 1: mux_19848 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19849;
  function [0:0] mux_19849(input [0:0] sel);
    case (sel) 0: mux_19849 = 1'h0; 1: mux_19849 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19850;
  wire [0:0] v_19851;
  wire [0:0] v_19852;
  wire [0:0] v_19853;
  wire [0:0] v_19854;
  wire [0:0] v_19855;
  wire [0:0] v_19856;
  function [0:0] mux_19856(input [0:0] sel);
    case (sel) 0: mux_19856 = 1'h0; 1: mux_19856 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19857;
  wire [0:0] v_19858;
  wire [0:0] v_19859;
  wire [0:0] v_19860;
  wire [0:0] v_19861;
  function [0:0] mux_19861(input [0:0] sel);
    case (sel) 0: mux_19861 = 1'h0; 1: mux_19861 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19862;
  wire [0:0] v_19863;
  wire [0:0] v_19864;
  wire [0:0] v_19865;
  function [0:0] mux_19865(input [0:0] sel);
    case (sel) 0: mux_19865 = 1'h0; 1: mux_19865 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19866;
  function [0:0] mux_19866(input [0:0] sel);
    case (sel) 0: mux_19866 = 1'h0; 1: mux_19866 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_19867 = 1'h0;
  wire [0:0] v_19868;
  wire [0:0] v_19869;
  wire [0:0] act_19870;
  wire [0:0] v_19871;
  wire [0:0] v_19872;
  wire [0:0] v_19873;
  wire [0:0] vin0_consume_en_19874;
  wire [0:0] vout_canPeek_19874;
  wire [7:0] vout_peek_19874;
  wire [0:0] v_19875;
  wire [0:0] v_19876;
  function [0:0] mux_19876(input [0:0] sel);
    case (sel) 0: mux_19876 = 1'h0; 1: mux_19876 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19877;
  wire [0:0] v_19878;
  wire [0:0] v_19879;
  wire [0:0] v_19880;
  wire [0:0] v_19881;
  function [0:0] mux_19881(input [0:0] sel);
    case (sel) 0: mux_19881 = 1'h0; 1: mux_19881 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19882;
  wire [0:0] vin0_consume_en_19883;
  wire [0:0] vout_canPeek_19883;
  wire [7:0] vout_peek_19883;
  wire [0:0] v_19884;
  wire [0:0] v_19885;
  function [0:0] mux_19885(input [0:0] sel);
    case (sel) 0: mux_19885 = 1'h0; 1: mux_19885 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19886;
  function [0:0] mux_19886(input [0:0] sel);
    case (sel) 0: mux_19886 = 1'h0; 1: mux_19886 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19887;
  wire [0:0] v_19888;
  wire [0:0] v_19889;
  wire [0:0] v_19890;
  wire [0:0] v_19891;
  wire [0:0] v_19892;
  wire [0:0] v_19893;
  function [0:0] mux_19893(input [0:0] sel);
    case (sel) 0: mux_19893 = 1'h0; 1: mux_19893 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19894;
  function [0:0] mux_19894(input [0:0] sel);
    case (sel) 0: mux_19894 = 1'h0; 1: mux_19894 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19895;
  wire [0:0] v_19896;
  wire [0:0] v_19897;
  wire [0:0] v_19898;
  function [0:0] mux_19898(input [0:0] sel);
    case (sel) 0: mux_19898 = 1'h0; 1: mux_19898 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19899;
  function [0:0] mux_19899(input [0:0] sel);
    case (sel) 0: mux_19899 = 1'h0; 1: mux_19899 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19900;
  wire [0:0] v_19901;
  wire [0:0] v_19902;
  wire [0:0] v_19903;
  wire [0:0] v_19904;
  wire [0:0] v_19905;
  function [0:0] mux_19905(input [0:0] sel);
    case (sel) 0: mux_19905 = 1'h0; 1: mux_19905 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19906;
  wire [0:0] v_19907;
  wire [0:0] v_19908;
  wire [0:0] v_19909;
  wire [0:0] v_19910;
  function [0:0] mux_19910(input [0:0] sel);
    case (sel) 0: mux_19910 = 1'h0; 1: mux_19910 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19911;
  wire [0:0] v_19912;
  wire [0:0] v_19913;
  wire [0:0] v_19914;
  function [0:0] mux_19914(input [0:0] sel);
    case (sel) 0: mux_19914 = 1'h0; 1: mux_19914 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19915;
  function [0:0] mux_19915(input [0:0] sel);
    case (sel) 0: mux_19915 = 1'h0; 1: mux_19915 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_19916 = 1'h0;
  wire [0:0] v_19917;
  wire [0:0] v_19918;
  wire [0:0] act_19919;
  wire [0:0] v_19920;
  wire [0:0] v_19921;
  wire [0:0] v_19922;
  reg [0:0] v_19923 = 1'h0;
  wire [0:0] v_19924;
  wire [0:0] v_19925;
  wire [0:0] act_19926;
  wire [0:0] v_19927;
  wire [0:0] v_19928;
  wire [0:0] v_19929;
  wire [0:0] vin0_consume_en_19930;
  wire [0:0] vout_canPeek_19930;
  wire [7:0] vout_peek_19930;
  wire [0:0] v_19931;
  wire [0:0] v_19932;
  function [0:0] mux_19932(input [0:0] sel);
    case (sel) 0: mux_19932 = 1'h0; 1: mux_19932 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19933;
  wire [0:0] v_19934;
  wire [0:0] v_19935;
  wire [0:0] v_19936;
  wire [0:0] v_19937;
  function [0:0] mux_19937(input [0:0] sel);
    case (sel) 0: mux_19937 = 1'h0; 1: mux_19937 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19938;
  wire [0:0] vin0_consume_en_19939;
  wire [0:0] vout_canPeek_19939;
  wire [7:0] vout_peek_19939;
  wire [0:0] v_19940;
  wire [0:0] v_19941;
  function [0:0] mux_19941(input [0:0] sel);
    case (sel) 0: mux_19941 = 1'h0; 1: mux_19941 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19942;
  function [0:0] mux_19942(input [0:0] sel);
    case (sel) 0: mux_19942 = 1'h0; 1: mux_19942 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19943;
  wire [0:0] v_19944;
  wire [0:0] v_19945;
  wire [0:0] v_19946;
  wire [0:0] v_19947;
  wire [0:0] v_19948;
  wire [0:0] v_19949;
  function [0:0] mux_19949(input [0:0] sel);
    case (sel) 0: mux_19949 = 1'h0; 1: mux_19949 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19950;
  wire [0:0] v_19951;
  wire [0:0] v_19952;
  wire [0:0] v_19953;
  wire [0:0] v_19954;
  function [0:0] mux_19954(input [0:0] sel);
    case (sel) 0: mux_19954 = 1'h0; 1: mux_19954 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19955;
  wire [0:0] v_19956;
  wire [0:0] v_19957;
  wire [0:0] v_19958;
  function [0:0] mux_19958(input [0:0] sel);
    case (sel) 0: mux_19958 = 1'h0; 1: mux_19958 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19959;
  function [0:0] mux_19959(input [0:0] sel);
    case (sel) 0: mux_19959 = 1'h0; 1: mux_19959 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_19960 = 1'h0;
  wire [0:0] v_19961;
  wire [0:0] v_19962;
  wire [0:0] act_19963;
  wire [0:0] v_19964;
  wire [0:0] v_19965;
  wire [0:0] v_19966;
  wire [0:0] vin0_consume_en_19967;
  wire [0:0] vout_canPeek_19967;
  wire [7:0] vout_peek_19967;
  wire [0:0] v_19968;
  wire [0:0] v_19969;
  function [0:0] mux_19969(input [0:0] sel);
    case (sel) 0: mux_19969 = 1'h0; 1: mux_19969 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19970;
  wire [0:0] v_19971;
  wire [0:0] v_19972;
  wire [0:0] v_19973;
  wire [0:0] v_19974;
  function [0:0] mux_19974(input [0:0] sel);
    case (sel) 0: mux_19974 = 1'h0; 1: mux_19974 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19975;
  wire [0:0] vin0_consume_en_19976;
  wire [0:0] vout_canPeek_19976;
  wire [7:0] vout_peek_19976;
  wire [0:0] v_19977;
  wire [0:0] v_19978;
  function [0:0] mux_19978(input [0:0] sel);
    case (sel) 0: mux_19978 = 1'h0; 1: mux_19978 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19979;
  function [0:0] mux_19979(input [0:0] sel);
    case (sel) 0: mux_19979 = 1'h0; 1: mux_19979 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19980;
  wire [0:0] v_19981;
  wire [0:0] v_19982;
  wire [0:0] v_19983;
  wire [0:0] v_19984;
  wire [0:0] v_19985;
  wire [0:0] v_19986;
  function [0:0] mux_19986(input [0:0] sel);
    case (sel) 0: mux_19986 = 1'h0; 1: mux_19986 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19987;
  function [0:0] mux_19987(input [0:0] sel);
    case (sel) 0: mux_19987 = 1'h0; 1: mux_19987 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19988;
  wire [0:0] v_19989;
  wire [0:0] v_19990;
  wire [0:0] v_19991;
  function [0:0] mux_19991(input [0:0] sel);
    case (sel) 0: mux_19991 = 1'h0; 1: mux_19991 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19992;
  function [0:0] mux_19992(input [0:0] sel);
    case (sel) 0: mux_19992 = 1'h0; 1: mux_19992 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19993;
  wire [0:0] v_19994;
  wire [0:0] v_19995;
  wire [0:0] v_19996;
  wire [0:0] v_19997;
  wire [0:0] v_19998;
  function [0:0] mux_19998(input [0:0] sel);
    case (sel) 0: mux_19998 = 1'h0; 1: mux_19998 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_19999;
  function [0:0] mux_19999(input [0:0] sel);
    case (sel) 0: mux_19999 = 1'h0; 1: mux_19999 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20000;
  wire [0:0] v_20001;
  wire [0:0] v_20002;
  wire [0:0] v_20003;
  function [0:0] mux_20003(input [0:0] sel);
    case (sel) 0: mux_20003 = 1'h0; 1: mux_20003 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20004;
  function [0:0] mux_20004(input [0:0] sel);
    case (sel) 0: mux_20004 = 1'h0; 1: mux_20004 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20005;
  wire [0:0] v_20006;
  wire [0:0] v_20007;
  wire [0:0] v_20008;
  wire [0:0] v_20009;
  wire [0:0] v_20010;
  function [0:0] mux_20010(input [0:0] sel);
    case (sel) 0: mux_20010 = 1'h0; 1: mux_20010 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20011;
  function [0:0] mux_20011(input [0:0] sel);
    case (sel) 0: mux_20011 = 1'h0; 1: mux_20011 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20012;
  wire [0:0] v_20013;
  wire [0:0] v_20014;
  wire [0:0] v_20015;
  function [0:0] mux_20015(input [0:0] sel);
    case (sel) 0: mux_20015 = 1'h0; 1: mux_20015 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20016;
  function [0:0] mux_20016(input [0:0] sel);
    case (sel) 0: mux_20016 = 1'h0; 1: mux_20016 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20017;
  wire [0:0] v_20018;
  wire [0:0] v_20019;
  wire [0:0] v_20020;
  wire [0:0] v_20021;
  wire [0:0] v_20022;
  function [0:0] mux_20022(input [0:0] sel);
    case (sel) 0: mux_20022 = 1'h0; 1: mux_20022 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20023;
  wire [0:0] v_20024;
  wire [0:0] v_20025;
  wire [0:0] v_20026;
  wire [0:0] v_20027;
  function [0:0] mux_20027(input [0:0] sel);
    case (sel) 0: mux_20027 = 1'h0; 1: mux_20027 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20028;
  wire [0:0] v_20029;
  wire [0:0] v_20030;
  wire [0:0] v_20031;
  function [0:0] mux_20031(input [0:0] sel);
    case (sel) 0: mux_20031 = 1'h0; 1: mux_20031 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20032;
  function [0:0] mux_20032(input [0:0] sel);
    case (sel) 0: mux_20032 = 1'h0; 1: mux_20032 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_20033 = 1'h0;
  wire [0:0] v_20034;
  wire [0:0] v_20035;
  wire [0:0] act_20036;
  wire [0:0] v_20037;
  wire [0:0] v_20038;
  wire [0:0] v_20039;
  reg [0:0] v_20040 = 1'h0;
  wire [0:0] v_20041;
  wire [0:0] v_20042;
  wire [0:0] act_20043;
  wire [0:0] v_20044;
  wire [0:0] v_20045;
  wire [0:0] v_20046;
  reg [0:0] v_20047 = 1'h0;
  wire [0:0] v_20048;
  wire [0:0] v_20049;
  wire [0:0] act_20050;
  wire [0:0] v_20051;
  wire [0:0] v_20052;
  wire [0:0] v_20053;
  reg [0:0] v_20054 = 1'h0;
  wire [0:0] v_20055;
  wire [0:0] v_20056;
  wire [0:0] act_20057;
  wire [0:0] v_20058;
  wire [0:0] v_20059;
  wire [0:0] v_20060;
  wire [0:0] vin0_consume_en_20061;
  wire [0:0] vout_canPeek_20061;
  wire [7:0] vout_peek_20061;
  wire [0:0] v_20062;
  wire [0:0] v_20063;
  function [0:0] mux_20063(input [0:0] sel);
    case (sel) 0: mux_20063 = 1'h0; 1: mux_20063 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20064;
  wire [0:0] v_20065;
  wire [0:0] v_20066;
  wire [0:0] v_20067;
  wire [0:0] v_20068;
  function [0:0] mux_20068(input [0:0] sel);
    case (sel) 0: mux_20068 = 1'h0; 1: mux_20068 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20069;
  wire [0:0] vin0_consume_en_20070;
  wire [0:0] vout_canPeek_20070;
  wire [7:0] vout_peek_20070;
  wire [0:0] v_20071;
  wire [0:0] v_20072;
  function [0:0] mux_20072(input [0:0] sel);
    case (sel) 0: mux_20072 = 1'h0; 1: mux_20072 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20073;
  function [0:0] mux_20073(input [0:0] sel);
    case (sel) 0: mux_20073 = 1'h0; 1: mux_20073 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20074;
  wire [0:0] v_20075;
  wire [0:0] v_20076;
  wire [0:0] v_20077;
  wire [0:0] v_20078;
  wire [0:0] v_20079;
  wire [0:0] v_20080;
  function [0:0] mux_20080(input [0:0] sel);
    case (sel) 0: mux_20080 = 1'h0; 1: mux_20080 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20081;
  wire [0:0] v_20082;
  wire [0:0] v_20083;
  wire [0:0] v_20084;
  wire [0:0] v_20085;
  function [0:0] mux_20085(input [0:0] sel);
    case (sel) 0: mux_20085 = 1'h0; 1: mux_20085 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20086;
  wire [0:0] v_20087;
  wire [0:0] v_20088;
  wire [0:0] v_20089;
  function [0:0] mux_20089(input [0:0] sel);
    case (sel) 0: mux_20089 = 1'h0; 1: mux_20089 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20090;
  function [0:0] mux_20090(input [0:0] sel);
    case (sel) 0: mux_20090 = 1'h0; 1: mux_20090 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_20091 = 1'h0;
  wire [0:0] v_20092;
  wire [0:0] v_20093;
  wire [0:0] act_20094;
  wire [0:0] v_20095;
  wire [0:0] v_20096;
  wire [0:0] v_20097;
  wire [0:0] vin0_consume_en_20098;
  wire [0:0] vout_canPeek_20098;
  wire [7:0] vout_peek_20098;
  wire [0:0] v_20099;
  wire [0:0] v_20100;
  function [0:0] mux_20100(input [0:0] sel);
    case (sel) 0: mux_20100 = 1'h0; 1: mux_20100 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20101;
  wire [0:0] v_20102;
  wire [0:0] v_20103;
  wire [0:0] v_20104;
  wire [0:0] v_20105;
  function [0:0] mux_20105(input [0:0] sel);
    case (sel) 0: mux_20105 = 1'h0; 1: mux_20105 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20106;
  wire [0:0] vin0_consume_en_20107;
  wire [0:0] vout_canPeek_20107;
  wire [7:0] vout_peek_20107;
  wire [0:0] v_20108;
  wire [0:0] v_20109;
  function [0:0] mux_20109(input [0:0] sel);
    case (sel) 0: mux_20109 = 1'h0; 1: mux_20109 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20110;
  function [0:0] mux_20110(input [0:0] sel);
    case (sel) 0: mux_20110 = 1'h0; 1: mux_20110 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20111;
  wire [0:0] v_20112;
  wire [0:0] v_20113;
  wire [0:0] v_20114;
  wire [0:0] v_20115;
  wire [0:0] v_20116;
  wire [0:0] v_20117;
  function [0:0] mux_20117(input [0:0] sel);
    case (sel) 0: mux_20117 = 1'h0; 1: mux_20117 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20118;
  function [0:0] mux_20118(input [0:0] sel);
    case (sel) 0: mux_20118 = 1'h0; 1: mux_20118 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20119;
  wire [0:0] v_20120;
  wire [0:0] v_20121;
  wire [0:0] v_20122;
  function [0:0] mux_20122(input [0:0] sel);
    case (sel) 0: mux_20122 = 1'h0; 1: mux_20122 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20123;
  function [0:0] mux_20123(input [0:0] sel);
    case (sel) 0: mux_20123 = 1'h0; 1: mux_20123 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20124;
  wire [0:0] v_20125;
  wire [0:0] v_20126;
  wire [0:0] v_20127;
  wire [0:0] v_20128;
  wire [0:0] v_20129;
  function [0:0] mux_20129(input [0:0] sel);
    case (sel) 0: mux_20129 = 1'h0; 1: mux_20129 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20130;
  wire [0:0] v_20131;
  wire [0:0] v_20132;
  wire [0:0] v_20133;
  wire [0:0] v_20134;
  function [0:0] mux_20134(input [0:0] sel);
    case (sel) 0: mux_20134 = 1'h0; 1: mux_20134 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20135;
  wire [0:0] v_20136;
  wire [0:0] v_20137;
  wire [0:0] v_20138;
  function [0:0] mux_20138(input [0:0] sel);
    case (sel) 0: mux_20138 = 1'h0; 1: mux_20138 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20139;
  function [0:0] mux_20139(input [0:0] sel);
    case (sel) 0: mux_20139 = 1'h0; 1: mux_20139 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_20140 = 1'h0;
  wire [0:0] v_20141;
  wire [0:0] v_20142;
  wire [0:0] act_20143;
  wire [0:0] v_20144;
  wire [0:0] v_20145;
  wire [0:0] v_20146;
  reg [0:0] v_20147 = 1'h0;
  wire [0:0] v_20148;
  wire [0:0] v_20149;
  wire [0:0] act_20150;
  wire [0:0] v_20151;
  wire [0:0] v_20152;
  wire [0:0] v_20153;
  wire [0:0] vin0_consume_en_20154;
  wire [0:0] vout_canPeek_20154;
  wire [7:0] vout_peek_20154;
  wire [0:0] v_20155;
  wire [0:0] v_20156;
  function [0:0] mux_20156(input [0:0] sel);
    case (sel) 0: mux_20156 = 1'h0; 1: mux_20156 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20157;
  wire [0:0] v_20158;
  wire [0:0] v_20159;
  wire [0:0] v_20160;
  wire [0:0] v_20161;
  function [0:0] mux_20161(input [0:0] sel);
    case (sel) 0: mux_20161 = 1'h0; 1: mux_20161 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20162;
  wire [0:0] vin0_consume_en_20163;
  wire [0:0] vout_canPeek_20163;
  wire [7:0] vout_peek_20163;
  wire [0:0] v_20164;
  wire [0:0] v_20165;
  function [0:0] mux_20165(input [0:0] sel);
    case (sel) 0: mux_20165 = 1'h0; 1: mux_20165 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20166;
  function [0:0] mux_20166(input [0:0] sel);
    case (sel) 0: mux_20166 = 1'h0; 1: mux_20166 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20167;
  wire [0:0] v_20168;
  wire [0:0] v_20169;
  wire [0:0] v_20170;
  wire [0:0] v_20171;
  wire [0:0] v_20172;
  wire [0:0] v_20173;
  function [0:0] mux_20173(input [0:0] sel);
    case (sel) 0: mux_20173 = 1'h0; 1: mux_20173 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20174;
  wire [0:0] v_20175;
  wire [0:0] v_20176;
  wire [0:0] v_20177;
  wire [0:0] v_20178;
  function [0:0] mux_20178(input [0:0] sel);
    case (sel) 0: mux_20178 = 1'h0; 1: mux_20178 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20179;
  wire [0:0] v_20180;
  wire [0:0] v_20181;
  wire [0:0] v_20182;
  function [0:0] mux_20182(input [0:0] sel);
    case (sel) 0: mux_20182 = 1'h0; 1: mux_20182 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20183;
  function [0:0] mux_20183(input [0:0] sel);
    case (sel) 0: mux_20183 = 1'h0; 1: mux_20183 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_20184 = 1'h0;
  wire [0:0] v_20185;
  wire [0:0] v_20186;
  wire [0:0] act_20187;
  wire [0:0] v_20188;
  wire [0:0] v_20189;
  wire [0:0] v_20190;
  wire [0:0] vin0_consume_en_20191;
  wire [0:0] vout_canPeek_20191;
  wire [7:0] vout_peek_20191;
  wire [0:0] v_20192;
  wire [0:0] v_20193;
  function [0:0] mux_20193(input [0:0] sel);
    case (sel) 0: mux_20193 = 1'h0; 1: mux_20193 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20194;
  wire [0:0] v_20195;
  wire [0:0] v_20196;
  wire [0:0] v_20197;
  wire [0:0] v_20198;
  function [0:0] mux_20198(input [0:0] sel);
    case (sel) 0: mux_20198 = 1'h0; 1: mux_20198 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20199;
  wire [0:0] vin0_consume_en_20200;
  wire [0:0] vout_canPeek_20200;
  wire [7:0] vout_peek_20200;
  wire [0:0] v_20201;
  wire [0:0] v_20202;
  function [0:0] mux_20202(input [0:0] sel);
    case (sel) 0: mux_20202 = 1'h0; 1: mux_20202 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20203;
  function [0:0] mux_20203(input [0:0] sel);
    case (sel) 0: mux_20203 = 1'h0; 1: mux_20203 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20204;
  wire [0:0] v_20205;
  wire [0:0] v_20206;
  wire [0:0] v_20207;
  wire [0:0] v_20208;
  wire [0:0] v_20209;
  wire [0:0] v_20210;
  function [0:0] mux_20210(input [0:0] sel);
    case (sel) 0: mux_20210 = 1'h0; 1: mux_20210 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20211;
  function [0:0] mux_20211(input [0:0] sel);
    case (sel) 0: mux_20211 = 1'h0; 1: mux_20211 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20212;
  wire [0:0] v_20213;
  wire [0:0] v_20214;
  wire [0:0] v_20215;
  function [0:0] mux_20215(input [0:0] sel);
    case (sel) 0: mux_20215 = 1'h0; 1: mux_20215 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20216;
  function [0:0] mux_20216(input [0:0] sel);
    case (sel) 0: mux_20216 = 1'h0; 1: mux_20216 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20217;
  wire [0:0] v_20218;
  wire [0:0] v_20219;
  wire [0:0] v_20220;
  wire [0:0] v_20221;
  wire [0:0] v_20222;
  function [0:0] mux_20222(input [0:0] sel);
    case (sel) 0: mux_20222 = 1'h0; 1: mux_20222 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20223;
  function [0:0] mux_20223(input [0:0] sel);
    case (sel) 0: mux_20223 = 1'h0; 1: mux_20223 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20224;
  wire [0:0] v_20225;
  wire [0:0] v_20226;
  wire [0:0] v_20227;
  function [0:0] mux_20227(input [0:0] sel);
    case (sel) 0: mux_20227 = 1'h0; 1: mux_20227 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20228;
  function [0:0] mux_20228(input [0:0] sel);
    case (sel) 0: mux_20228 = 1'h0; 1: mux_20228 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20229;
  wire [0:0] v_20230;
  wire [0:0] v_20231;
  wire [0:0] v_20232;
  wire [0:0] v_20233;
  wire [0:0] v_20234;
  function [0:0] mux_20234(input [0:0] sel);
    case (sel) 0: mux_20234 = 1'h0; 1: mux_20234 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20235;
  wire [0:0] v_20236;
  wire [0:0] v_20237;
  wire [0:0] v_20238;
  wire [0:0] v_20239;
  function [0:0] mux_20239(input [0:0] sel);
    case (sel) 0: mux_20239 = 1'h0; 1: mux_20239 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20240;
  wire [0:0] v_20241;
  wire [0:0] v_20242;
  wire [0:0] v_20243;
  function [0:0] mux_20243(input [0:0] sel);
    case (sel) 0: mux_20243 = 1'h0; 1: mux_20243 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20244;
  function [0:0] mux_20244(input [0:0] sel);
    case (sel) 0: mux_20244 = 1'h0; 1: mux_20244 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_20245 = 1'h0;
  wire [0:0] v_20246;
  wire [0:0] v_20247;
  wire [0:0] act_20248;
  wire [0:0] v_20249;
  wire [0:0] v_20250;
  wire [0:0] v_20251;
  reg [0:0] v_20252 = 1'h0;
  wire [0:0] v_20253;
  wire [0:0] v_20254;
  wire [0:0] act_20255;
  wire [0:0] v_20256;
  wire [0:0] v_20257;
  wire [0:0] v_20258;
  reg [0:0] v_20259 = 1'h0;
  wire [0:0] v_20260;
  wire [0:0] v_20261;
  wire [0:0] act_20262;
  wire [0:0] v_20263;
  wire [0:0] v_20264;
  wire [0:0] v_20265;
  wire [0:0] vin0_consume_en_20266;
  wire [0:0] vout_canPeek_20266;
  wire [7:0] vout_peek_20266;
  wire [0:0] v_20267;
  wire [0:0] v_20268;
  function [0:0] mux_20268(input [0:0] sel);
    case (sel) 0: mux_20268 = 1'h0; 1: mux_20268 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20269;
  wire [0:0] v_20270;
  wire [0:0] v_20271;
  wire [0:0] v_20272;
  wire [0:0] v_20273;
  function [0:0] mux_20273(input [0:0] sel);
    case (sel) 0: mux_20273 = 1'h0; 1: mux_20273 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20274;
  wire [0:0] vin0_consume_en_20275;
  wire [0:0] vout_canPeek_20275;
  wire [7:0] vout_peek_20275;
  wire [0:0] v_20276;
  wire [0:0] v_20277;
  function [0:0] mux_20277(input [0:0] sel);
    case (sel) 0: mux_20277 = 1'h0; 1: mux_20277 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20278;
  function [0:0] mux_20278(input [0:0] sel);
    case (sel) 0: mux_20278 = 1'h0; 1: mux_20278 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20279;
  wire [0:0] v_20280;
  wire [0:0] v_20281;
  wire [0:0] v_20282;
  wire [0:0] v_20283;
  wire [0:0] v_20284;
  wire [0:0] v_20285;
  function [0:0] mux_20285(input [0:0] sel);
    case (sel) 0: mux_20285 = 1'h0; 1: mux_20285 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20286;
  wire [0:0] v_20287;
  wire [0:0] v_20288;
  wire [0:0] v_20289;
  wire [0:0] v_20290;
  function [0:0] mux_20290(input [0:0] sel);
    case (sel) 0: mux_20290 = 1'h0; 1: mux_20290 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20291;
  wire [0:0] v_20292;
  wire [0:0] v_20293;
  wire [0:0] v_20294;
  function [0:0] mux_20294(input [0:0] sel);
    case (sel) 0: mux_20294 = 1'h0; 1: mux_20294 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20295;
  function [0:0] mux_20295(input [0:0] sel);
    case (sel) 0: mux_20295 = 1'h0; 1: mux_20295 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_20296 = 1'h0;
  wire [0:0] v_20297;
  wire [0:0] v_20298;
  wire [0:0] act_20299;
  wire [0:0] v_20300;
  wire [0:0] v_20301;
  wire [0:0] v_20302;
  wire [0:0] vin0_consume_en_20303;
  wire [0:0] vout_canPeek_20303;
  wire [7:0] vout_peek_20303;
  wire [0:0] v_20304;
  wire [0:0] v_20305;
  function [0:0] mux_20305(input [0:0] sel);
    case (sel) 0: mux_20305 = 1'h0; 1: mux_20305 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20306;
  wire [0:0] v_20307;
  wire [0:0] v_20308;
  wire [0:0] v_20309;
  wire [0:0] v_20310;
  function [0:0] mux_20310(input [0:0] sel);
    case (sel) 0: mux_20310 = 1'h0; 1: mux_20310 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20311;
  wire [0:0] vin0_consume_en_20312;
  wire [0:0] vout_canPeek_20312;
  wire [7:0] vout_peek_20312;
  wire [0:0] v_20313;
  wire [0:0] v_20314;
  function [0:0] mux_20314(input [0:0] sel);
    case (sel) 0: mux_20314 = 1'h0; 1: mux_20314 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20315;
  function [0:0] mux_20315(input [0:0] sel);
    case (sel) 0: mux_20315 = 1'h0; 1: mux_20315 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20316;
  wire [0:0] v_20317;
  wire [0:0] v_20318;
  wire [0:0] v_20319;
  wire [0:0] v_20320;
  wire [0:0] v_20321;
  wire [0:0] v_20322;
  function [0:0] mux_20322(input [0:0] sel);
    case (sel) 0: mux_20322 = 1'h0; 1: mux_20322 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20323;
  function [0:0] mux_20323(input [0:0] sel);
    case (sel) 0: mux_20323 = 1'h0; 1: mux_20323 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20324;
  wire [0:0] v_20325;
  wire [0:0] v_20326;
  wire [0:0] v_20327;
  function [0:0] mux_20327(input [0:0] sel);
    case (sel) 0: mux_20327 = 1'h0; 1: mux_20327 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20328;
  function [0:0] mux_20328(input [0:0] sel);
    case (sel) 0: mux_20328 = 1'h0; 1: mux_20328 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20329;
  wire [0:0] v_20330;
  wire [0:0] v_20331;
  wire [0:0] v_20332;
  wire [0:0] v_20333;
  wire [0:0] v_20334;
  function [0:0] mux_20334(input [0:0] sel);
    case (sel) 0: mux_20334 = 1'h0; 1: mux_20334 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20335;
  wire [0:0] v_20336;
  wire [0:0] v_20337;
  wire [0:0] v_20338;
  wire [0:0] v_20339;
  function [0:0] mux_20339(input [0:0] sel);
    case (sel) 0: mux_20339 = 1'h0; 1: mux_20339 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20340;
  wire [0:0] v_20341;
  wire [0:0] v_20342;
  wire [0:0] v_20343;
  function [0:0] mux_20343(input [0:0] sel);
    case (sel) 0: mux_20343 = 1'h0; 1: mux_20343 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20344;
  function [0:0] mux_20344(input [0:0] sel);
    case (sel) 0: mux_20344 = 1'h0; 1: mux_20344 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_20345 = 1'h0;
  wire [0:0] v_20346;
  wire [0:0] v_20347;
  wire [0:0] act_20348;
  wire [0:0] v_20349;
  wire [0:0] v_20350;
  wire [0:0] v_20351;
  reg [0:0] v_20352 = 1'h0;
  wire [0:0] v_20353;
  wire [0:0] v_20354;
  wire [0:0] act_20355;
  wire [0:0] v_20356;
  wire [0:0] v_20357;
  wire [0:0] v_20358;
  wire [0:0] vin0_consume_en_20359;
  wire [0:0] vout_canPeek_20359;
  wire [7:0] vout_peek_20359;
  wire [0:0] v_20360;
  wire [0:0] v_20361;
  function [0:0] mux_20361(input [0:0] sel);
    case (sel) 0: mux_20361 = 1'h0; 1: mux_20361 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20362;
  wire [0:0] v_20363;
  wire [0:0] v_20364;
  wire [0:0] v_20365;
  wire [0:0] v_20366;
  function [0:0] mux_20366(input [0:0] sel);
    case (sel) 0: mux_20366 = 1'h0; 1: mux_20366 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20367;
  wire [0:0] vin0_consume_en_20368;
  wire [0:0] vout_canPeek_20368;
  wire [7:0] vout_peek_20368;
  wire [0:0] v_20369;
  wire [0:0] v_20370;
  function [0:0] mux_20370(input [0:0] sel);
    case (sel) 0: mux_20370 = 1'h0; 1: mux_20370 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20371;
  function [0:0] mux_20371(input [0:0] sel);
    case (sel) 0: mux_20371 = 1'h0; 1: mux_20371 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20372;
  wire [0:0] v_20373;
  wire [0:0] v_20374;
  wire [0:0] v_20375;
  wire [0:0] v_20376;
  wire [0:0] v_20377;
  wire [0:0] v_20378;
  function [0:0] mux_20378(input [0:0] sel);
    case (sel) 0: mux_20378 = 1'h0; 1: mux_20378 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20379;
  wire [0:0] v_20380;
  wire [0:0] v_20381;
  wire [0:0] v_20382;
  wire [0:0] v_20383;
  function [0:0] mux_20383(input [0:0] sel);
    case (sel) 0: mux_20383 = 1'h0; 1: mux_20383 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20384;
  wire [0:0] v_20385;
  wire [0:0] v_20386;
  wire [0:0] v_20387;
  function [0:0] mux_20387(input [0:0] sel);
    case (sel) 0: mux_20387 = 1'h0; 1: mux_20387 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20388;
  function [0:0] mux_20388(input [0:0] sel);
    case (sel) 0: mux_20388 = 1'h0; 1: mux_20388 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_20389 = 1'h0;
  wire [0:0] v_20390;
  wire [0:0] v_20391;
  wire [0:0] act_20392;
  wire [0:0] v_20393;
  wire [0:0] v_20394;
  wire [0:0] v_20395;
  wire [0:0] vin0_consume_en_20396;
  wire [0:0] vout_canPeek_20396;
  wire [7:0] vout_peek_20396;
  wire [0:0] v_20397;
  wire [0:0] v_20398;
  function [0:0] mux_20398(input [0:0] sel);
    case (sel) 0: mux_20398 = 1'h0; 1: mux_20398 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20399;
  wire [0:0] v_20400;
  wire [0:0] v_20401;
  wire [0:0] v_20402;
  wire [0:0] v_20403;
  function [0:0] mux_20403(input [0:0] sel);
    case (sel) 0: mux_20403 = 1'h0; 1: mux_20403 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20404;
  wire [0:0] vin0_consume_en_20405;
  wire [0:0] vout_canPeek_20405;
  wire [7:0] vout_peek_20405;
  wire [0:0] v_20406;
  wire [0:0] v_20407;
  function [0:0] mux_20407(input [0:0] sel);
    case (sel) 0: mux_20407 = 1'h0; 1: mux_20407 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20408;
  function [0:0] mux_20408(input [0:0] sel);
    case (sel) 0: mux_20408 = 1'h0; 1: mux_20408 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20409;
  wire [0:0] v_20410;
  wire [0:0] v_20411;
  wire [0:0] v_20412;
  wire [0:0] v_20413;
  wire [0:0] v_20414;
  wire [0:0] v_20415;
  function [0:0] mux_20415(input [0:0] sel);
    case (sel) 0: mux_20415 = 1'h0; 1: mux_20415 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20416;
  function [0:0] mux_20416(input [0:0] sel);
    case (sel) 0: mux_20416 = 1'h0; 1: mux_20416 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20417;
  wire [0:0] v_20418;
  wire [0:0] v_20419;
  wire [0:0] v_20420;
  function [0:0] mux_20420(input [0:0] sel);
    case (sel) 0: mux_20420 = 1'h0; 1: mux_20420 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20421;
  function [0:0] mux_20421(input [0:0] sel);
    case (sel) 0: mux_20421 = 1'h0; 1: mux_20421 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20422;
  wire [0:0] v_20423;
  wire [0:0] v_20424;
  wire [0:0] v_20425;
  wire [0:0] v_20426;
  wire [0:0] v_20427;
  function [0:0] mux_20427(input [0:0] sel);
    case (sel) 0: mux_20427 = 1'h0; 1: mux_20427 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20428;
  function [0:0] mux_20428(input [0:0] sel);
    case (sel) 0: mux_20428 = 1'h0; 1: mux_20428 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20429;
  wire [0:0] v_20430;
  wire [0:0] v_20431;
  wire [0:0] v_20432;
  function [0:0] mux_20432(input [0:0] sel);
    case (sel) 0: mux_20432 = 1'h0; 1: mux_20432 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20433;
  function [0:0] mux_20433(input [0:0] sel);
    case (sel) 0: mux_20433 = 1'h0; 1: mux_20433 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20434;
  wire [0:0] v_20435;
  wire [0:0] v_20436;
  wire [0:0] v_20437;
  wire [0:0] v_20438;
  wire [0:0] v_20439;
  function [0:0] mux_20439(input [0:0] sel);
    case (sel) 0: mux_20439 = 1'h0; 1: mux_20439 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20440;
  function [0:0] mux_20440(input [0:0] sel);
    case (sel) 0: mux_20440 = 1'h0; 1: mux_20440 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20441;
  wire [0:0] v_20442;
  wire [0:0] v_20443;
  wire [0:0] v_20444;
  function [0:0] mux_20444(input [0:0] sel);
    case (sel) 0: mux_20444 = 1'h0; 1: mux_20444 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20445;
  function [0:0] mux_20445(input [0:0] sel);
    case (sel) 0: mux_20445 = 1'h0; 1: mux_20445 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20446;
  wire [0:0] v_20447;
  wire [0:0] v_20448;
  wire [0:0] v_20449;
  wire [0:0] v_20450;
  wire [0:0] v_20451;
  function [0:0] mux_20451(input [0:0] sel);
    case (sel) 0: mux_20451 = 1'h0; 1: mux_20451 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20452;
  function [0:0] mux_20452(input [0:0] sel);
    case (sel) 0: mux_20452 = 1'h0; 1: mux_20452 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20453;
  wire [0:0] v_20454;
  wire [0:0] v_20455;
  wire [0:0] v_20456;
  function [0:0] mux_20456(input [0:0] sel);
    case (sel) 0: mux_20456 = 1'h0; 1: mux_20456 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20457;
  function [0:0] mux_20457(input [0:0] sel);
    case (sel) 0: mux_20457 = 1'h0; 1: mux_20457 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20458;
  wire [0:0] v_20459;
  wire [0:0] v_20460;
  wire [0:0] v_20461;
  wire [0:0] v_20462;
  wire [0:0] v_20463;
  function [0:0] mux_20463(input [0:0] sel);
    case (sel) 0: mux_20463 = 1'h0; 1: mux_20463 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20464;
  function [0:0] mux_20464(input [0:0] sel);
    case (sel) 0: mux_20464 = 1'h0; 1: mux_20464 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20465;
  wire [0:0] v_20466;
  wire [0:0] v_20467;
  wire [0:0] v_20468;
  function [0:0] mux_20468(input [0:0] sel);
    case (sel) 0: mux_20468 = 1'h0; 1: mux_20468 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20469;
  function [0:0] mux_20469(input [0:0] sel);
    case (sel) 0: mux_20469 = 1'h0; 1: mux_20469 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20470;
  wire [0:0] v_20471;
  wire [0:0] v_20472;
  wire [0:0] v_20473;
  wire [0:0] v_20474;
  wire [0:0] v_20475;
  function [0:0] mux_20475(input [0:0] sel);
    case (sel) 0: mux_20475 = 1'h0; 1: mux_20475 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20476;
  wire [0:0] v_20477;
  wire [0:0] v_20478;
  wire [0:0] v_20479;
  wire [0:0] v_20480;
  function [0:0] mux_20480(input [0:0] sel);
    case (sel) 0: mux_20480 = 1'h0; 1: mux_20480 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20481;
  wire [0:0] v_20482;
  wire [0:0] v_20483;
  wire [0:0] v_20484;
  function [0:0] mux_20484(input [0:0] sel);
    case (sel) 0: mux_20484 = 1'h0; 1: mux_20484 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20485;
  function [0:0] mux_20485(input [0:0] sel);
    case (sel) 0: mux_20485 = 1'h0; 1: mux_20485 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_20486 = 1'h0;
  wire [0:0] v_20487;
  wire [0:0] v_20488;
  wire [0:0] act_20489;
  wire [0:0] v_20490;
  wire [0:0] v_20491;
  wire [0:0] v_20492;
  reg [0:0] v_20493 = 1'h0;
  wire [0:0] v_20494;
  wire [0:0] v_20495;
  wire [0:0] act_20496;
  wire [0:0] v_20497;
  wire [0:0] v_20498;
  wire [0:0] v_20499;
  reg [0:0] v_20500 = 1'h0;
  wire [0:0] v_20501;
  wire [0:0] v_20502;
  wire [0:0] act_20503;
  wire [0:0] v_20504;
  wire [0:0] v_20505;
  wire [0:0] v_20506;
  reg [0:0] v_20507 = 1'h0;
  wire [0:0] v_20508;
  wire [0:0] v_20509;
  wire [0:0] act_20510;
  wire [0:0] v_20511;
  wire [0:0] v_20512;
  wire [0:0] v_20513;
  reg [0:0] v_20514 = 1'h0;
  wire [0:0] v_20515;
  wire [0:0] v_20516;
  wire [0:0] act_20517;
  wire [0:0] v_20518;
  wire [0:0] v_20519;
  wire [0:0] v_20520;
  reg [0:0] v_20521 = 1'h0;
  wire [0:0] v_20522;
  wire [0:0] v_20523;
  wire [0:0] act_20524;
  wire [0:0] v_20525;
  wire [0:0] v_20526;
  wire [0:0] v_20527;
  wire [0:0] vin0_consume_en_20528;
  wire [0:0] vout_canPeek_20528;
  wire [7:0] vout_peek_20528;
  wire [0:0] v_20529;
  wire [0:0] v_20530;
  function [0:0] mux_20530(input [0:0] sel);
    case (sel) 0: mux_20530 = 1'h0; 1: mux_20530 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20531;
  wire [0:0] v_20532;
  wire [0:0] v_20533;
  wire [0:0] v_20534;
  wire [0:0] v_20535;
  function [0:0] mux_20535(input [0:0] sel);
    case (sel) 0: mux_20535 = 1'h0; 1: mux_20535 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20536;
  wire [0:0] vin0_consume_en_20537;
  wire [0:0] vout_canPeek_20537;
  wire [7:0] vout_peek_20537;
  wire [0:0] v_20538;
  wire [0:0] v_20539;
  function [0:0] mux_20539(input [0:0] sel);
    case (sel) 0: mux_20539 = 1'h0; 1: mux_20539 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20540;
  function [0:0] mux_20540(input [0:0] sel);
    case (sel) 0: mux_20540 = 1'h0; 1: mux_20540 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20541;
  wire [0:0] v_20542;
  wire [0:0] v_20543;
  wire [0:0] v_20544;
  wire [0:0] v_20545;
  wire [0:0] v_20546;
  wire [0:0] v_20547;
  function [0:0] mux_20547(input [0:0] sel);
    case (sel) 0: mux_20547 = 1'h0; 1: mux_20547 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20548;
  wire [0:0] v_20549;
  wire [0:0] v_20550;
  wire [0:0] v_20551;
  wire [0:0] v_20552;
  function [0:0] mux_20552(input [0:0] sel);
    case (sel) 0: mux_20552 = 1'h0; 1: mux_20552 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20553;
  wire [0:0] v_20554;
  wire [0:0] v_20555;
  wire [0:0] v_20556;
  function [0:0] mux_20556(input [0:0] sel);
    case (sel) 0: mux_20556 = 1'h0; 1: mux_20556 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20557;
  function [0:0] mux_20557(input [0:0] sel);
    case (sel) 0: mux_20557 = 1'h0; 1: mux_20557 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_20558 = 1'h0;
  wire [0:0] v_20559;
  wire [0:0] v_20560;
  wire [0:0] act_20561;
  wire [0:0] v_20562;
  wire [0:0] v_20563;
  wire [0:0] v_20564;
  wire [0:0] vin0_consume_en_20565;
  wire [0:0] vout_canPeek_20565;
  wire [7:0] vout_peek_20565;
  wire [0:0] v_20566;
  wire [0:0] v_20567;
  function [0:0] mux_20567(input [0:0] sel);
    case (sel) 0: mux_20567 = 1'h0; 1: mux_20567 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20568;
  wire [0:0] v_20569;
  wire [0:0] v_20570;
  wire [0:0] v_20571;
  wire [0:0] v_20572;
  function [0:0] mux_20572(input [0:0] sel);
    case (sel) 0: mux_20572 = 1'h0; 1: mux_20572 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20573;
  wire [0:0] vin0_consume_en_20574;
  wire [0:0] vout_canPeek_20574;
  wire [7:0] vout_peek_20574;
  wire [0:0] v_20575;
  wire [0:0] v_20576;
  function [0:0] mux_20576(input [0:0] sel);
    case (sel) 0: mux_20576 = 1'h0; 1: mux_20576 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20577;
  function [0:0] mux_20577(input [0:0] sel);
    case (sel) 0: mux_20577 = 1'h0; 1: mux_20577 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20578;
  wire [0:0] v_20579;
  wire [0:0] v_20580;
  wire [0:0] v_20581;
  wire [0:0] v_20582;
  wire [0:0] v_20583;
  wire [0:0] v_20584;
  function [0:0] mux_20584(input [0:0] sel);
    case (sel) 0: mux_20584 = 1'h0; 1: mux_20584 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20585;
  function [0:0] mux_20585(input [0:0] sel);
    case (sel) 0: mux_20585 = 1'h0; 1: mux_20585 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20586;
  wire [0:0] v_20587;
  wire [0:0] v_20588;
  wire [0:0] v_20589;
  function [0:0] mux_20589(input [0:0] sel);
    case (sel) 0: mux_20589 = 1'h0; 1: mux_20589 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20590;
  function [0:0] mux_20590(input [0:0] sel);
    case (sel) 0: mux_20590 = 1'h0; 1: mux_20590 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20591;
  wire [0:0] v_20592;
  wire [0:0] v_20593;
  wire [0:0] v_20594;
  wire [0:0] v_20595;
  wire [0:0] v_20596;
  function [0:0] mux_20596(input [0:0] sel);
    case (sel) 0: mux_20596 = 1'h0; 1: mux_20596 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20597;
  wire [0:0] v_20598;
  wire [0:0] v_20599;
  wire [0:0] v_20600;
  wire [0:0] v_20601;
  function [0:0] mux_20601(input [0:0] sel);
    case (sel) 0: mux_20601 = 1'h0; 1: mux_20601 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20602;
  wire [0:0] v_20603;
  wire [0:0] v_20604;
  wire [0:0] v_20605;
  function [0:0] mux_20605(input [0:0] sel);
    case (sel) 0: mux_20605 = 1'h0; 1: mux_20605 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20606;
  function [0:0] mux_20606(input [0:0] sel);
    case (sel) 0: mux_20606 = 1'h0; 1: mux_20606 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_20607 = 1'h0;
  wire [0:0] v_20608;
  wire [0:0] v_20609;
  wire [0:0] act_20610;
  wire [0:0] v_20611;
  wire [0:0] v_20612;
  wire [0:0] v_20613;
  reg [0:0] v_20614 = 1'h0;
  wire [0:0] v_20615;
  wire [0:0] v_20616;
  wire [0:0] act_20617;
  wire [0:0] v_20618;
  wire [0:0] v_20619;
  wire [0:0] v_20620;
  wire [0:0] vin0_consume_en_20621;
  wire [0:0] vout_canPeek_20621;
  wire [7:0] vout_peek_20621;
  wire [0:0] v_20622;
  wire [0:0] v_20623;
  function [0:0] mux_20623(input [0:0] sel);
    case (sel) 0: mux_20623 = 1'h0; 1: mux_20623 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20624;
  wire [0:0] v_20625;
  wire [0:0] v_20626;
  wire [0:0] v_20627;
  wire [0:0] v_20628;
  function [0:0] mux_20628(input [0:0] sel);
    case (sel) 0: mux_20628 = 1'h0; 1: mux_20628 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20629;
  wire [0:0] vin0_consume_en_20630;
  wire [0:0] vout_canPeek_20630;
  wire [7:0] vout_peek_20630;
  wire [0:0] v_20631;
  wire [0:0] v_20632;
  function [0:0] mux_20632(input [0:0] sel);
    case (sel) 0: mux_20632 = 1'h0; 1: mux_20632 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20633;
  function [0:0] mux_20633(input [0:0] sel);
    case (sel) 0: mux_20633 = 1'h0; 1: mux_20633 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20634;
  wire [0:0] v_20635;
  wire [0:0] v_20636;
  wire [0:0] v_20637;
  wire [0:0] v_20638;
  wire [0:0] v_20639;
  wire [0:0] v_20640;
  function [0:0] mux_20640(input [0:0] sel);
    case (sel) 0: mux_20640 = 1'h0; 1: mux_20640 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20641;
  wire [0:0] v_20642;
  wire [0:0] v_20643;
  wire [0:0] v_20644;
  wire [0:0] v_20645;
  function [0:0] mux_20645(input [0:0] sel);
    case (sel) 0: mux_20645 = 1'h0; 1: mux_20645 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20646;
  wire [0:0] v_20647;
  wire [0:0] v_20648;
  wire [0:0] v_20649;
  function [0:0] mux_20649(input [0:0] sel);
    case (sel) 0: mux_20649 = 1'h0; 1: mux_20649 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20650;
  function [0:0] mux_20650(input [0:0] sel);
    case (sel) 0: mux_20650 = 1'h0; 1: mux_20650 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_20651 = 1'h0;
  wire [0:0] v_20652;
  wire [0:0] v_20653;
  wire [0:0] act_20654;
  wire [0:0] v_20655;
  wire [0:0] v_20656;
  wire [0:0] v_20657;
  wire [0:0] vin0_consume_en_20658;
  wire [0:0] vout_canPeek_20658;
  wire [7:0] vout_peek_20658;
  wire [0:0] v_20659;
  wire [0:0] v_20660;
  function [0:0] mux_20660(input [0:0] sel);
    case (sel) 0: mux_20660 = 1'h0; 1: mux_20660 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20661;
  wire [0:0] v_20662;
  wire [0:0] v_20663;
  wire [0:0] v_20664;
  wire [0:0] v_20665;
  function [0:0] mux_20665(input [0:0] sel);
    case (sel) 0: mux_20665 = 1'h0; 1: mux_20665 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20666;
  wire [0:0] vin0_consume_en_20667;
  wire [0:0] vout_canPeek_20667;
  wire [7:0] vout_peek_20667;
  wire [0:0] v_20668;
  wire [0:0] v_20669;
  function [0:0] mux_20669(input [0:0] sel);
    case (sel) 0: mux_20669 = 1'h0; 1: mux_20669 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20670;
  function [0:0] mux_20670(input [0:0] sel);
    case (sel) 0: mux_20670 = 1'h0; 1: mux_20670 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20671;
  wire [0:0] v_20672;
  wire [0:0] v_20673;
  wire [0:0] v_20674;
  wire [0:0] v_20675;
  wire [0:0] v_20676;
  wire [0:0] v_20677;
  function [0:0] mux_20677(input [0:0] sel);
    case (sel) 0: mux_20677 = 1'h0; 1: mux_20677 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20678;
  function [0:0] mux_20678(input [0:0] sel);
    case (sel) 0: mux_20678 = 1'h0; 1: mux_20678 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20679;
  wire [0:0] v_20680;
  wire [0:0] v_20681;
  wire [0:0] v_20682;
  function [0:0] mux_20682(input [0:0] sel);
    case (sel) 0: mux_20682 = 1'h0; 1: mux_20682 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20683;
  function [0:0] mux_20683(input [0:0] sel);
    case (sel) 0: mux_20683 = 1'h0; 1: mux_20683 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20684;
  wire [0:0] v_20685;
  wire [0:0] v_20686;
  wire [0:0] v_20687;
  wire [0:0] v_20688;
  wire [0:0] v_20689;
  function [0:0] mux_20689(input [0:0] sel);
    case (sel) 0: mux_20689 = 1'h0; 1: mux_20689 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20690;
  function [0:0] mux_20690(input [0:0] sel);
    case (sel) 0: mux_20690 = 1'h0; 1: mux_20690 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20691;
  wire [0:0] v_20692;
  wire [0:0] v_20693;
  wire [0:0] v_20694;
  function [0:0] mux_20694(input [0:0] sel);
    case (sel) 0: mux_20694 = 1'h0; 1: mux_20694 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20695;
  function [0:0] mux_20695(input [0:0] sel);
    case (sel) 0: mux_20695 = 1'h0; 1: mux_20695 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20696;
  wire [0:0] v_20697;
  wire [0:0] v_20698;
  wire [0:0] v_20699;
  wire [0:0] v_20700;
  wire [0:0] v_20701;
  function [0:0] mux_20701(input [0:0] sel);
    case (sel) 0: mux_20701 = 1'h0; 1: mux_20701 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20702;
  wire [0:0] v_20703;
  wire [0:0] v_20704;
  wire [0:0] v_20705;
  wire [0:0] v_20706;
  function [0:0] mux_20706(input [0:0] sel);
    case (sel) 0: mux_20706 = 1'h0; 1: mux_20706 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20707;
  wire [0:0] v_20708;
  wire [0:0] v_20709;
  wire [0:0] v_20710;
  function [0:0] mux_20710(input [0:0] sel);
    case (sel) 0: mux_20710 = 1'h0; 1: mux_20710 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20711;
  function [0:0] mux_20711(input [0:0] sel);
    case (sel) 0: mux_20711 = 1'h0; 1: mux_20711 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_20712 = 1'h0;
  wire [0:0] v_20713;
  wire [0:0] v_20714;
  wire [0:0] act_20715;
  wire [0:0] v_20716;
  wire [0:0] v_20717;
  wire [0:0] v_20718;
  reg [0:0] v_20719 = 1'h0;
  wire [0:0] v_20720;
  wire [0:0] v_20721;
  wire [0:0] act_20722;
  wire [0:0] v_20723;
  wire [0:0] v_20724;
  wire [0:0] v_20725;
  reg [0:0] v_20726 = 1'h0;
  wire [0:0] v_20727;
  wire [0:0] v_20728;
  wire [0:0] act_20729;
  wire [0:0] v_20730;
  wire [0:0] v_20731;
  wire [0:0] v_20732;
  wire [0:0] vin0_consume_en_20733;
  wire [0:0] vout_canPeek_20733;
  wire [7:0] vout_peek_20733;
  wire [0:0] v_20734;
  wire [0:0] v_20735;
  function [0:0] mux_20735(input [0:0] sel);
    case (sel) 0: mux_20735 = 1'h0; 1: mux_20735 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20736;
  wire [0:0] v_20737;
  wire [0:0] v_20738;
  wire [0:0] v_20739;
  wire [0:0] v_20740;
  function [0:0] mux_20740(input [0:0] sel);
    case (sel) 0: mux_20740 = 1'h0; 1: mux_20740 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20741;
  wire [0:0] vin0_consume_en_20742;
  wire [0:0] vout_canPeek_20742;
  wire [7:0] vout_peek_20742;
  wire [0:0] v_20743;
  wire [0:0] v_20744;
  function [0:0] mux_20744(input [0:0] sel);
    case (sel) 0: mux_20744 = 1'h0; 1: mux_20744 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20745;
  function [0:0] mux_20745(input [0:0] sel);
    case (sel) 0: mux_20745 = 1'h0; 1: mux_20745 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20746;
  wire [0:0] v_20747;
  wire [0:0] v_20748;
  wire [0:0] v_20749;
  wire [0:0] v_20750;
  wire [0:0] v_20751;
  wire [0:0] v_20752;
  function [0:0] mux_20752(input [0:0] sel);
    case (sel) 0: mux_20752 = 1'h0; 1: mux_20752 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20753;
  wire [0:0] v_20754;
  wire [0:0] v_20755;
  wire [0:0] v_20756;
  wire [0:0] v_20757;
  function [0:0] mux_20757(input [0:0] sel);
    case (sel) 0: mux_20757 = 1'h0; 1: mux_20757 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20758;
  wire [0:0] v_20759;
  wire [0:0] v_20760;
  wire [0:0] v_20761;
  function [0:0] mux_20761(input [0:0] sel);
    case (sel) 0: mux_20761 = 1'h0; 1: mux_20761 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20762;
  function [0:0] mux_20762(input [0:0] sel);
    case (sel) 0: mux_20762 = 1'h0; 1: mux_20762 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_20763 = 1'h0;
  wire [0:0] v_20764;
  wire [0:0] v_20765;
  wire [0:0] act_20766;
  wire [0:0] v_20767;
  wire [0:0] v_20768;
  wire [0:0] v_20769;
  wire [0:0] vin0_consume_en_20770;
  wire [0:0] vout_canPeek_20770;
  wire [7:0] vout_peek_20770;
  wire [0:0] v_20771;
  wire [0:0] v_20772;
  function [0:0] mux_20772(input [0:0] sel);
    case (sel) 0: mux_20772 = 1'h0; 1: mux_20772 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20773;
  wire [0:0] v_20774;
  wire [0:0] v_20775;
  wire [0:0] v_20776;
  wire [0:0] v_20777;
  function [0:0] mux_20777(input [0:0] sel);
    case (sel) 0: mux_20777 = 1'h0; 1: mux_20777 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20778;
  wire [0:0] vin0_consume_en_20779;
  wire [0:0] vout_canPeek_20779;
  wire [7:0] vout_peek_20779;
  wire [0:0] v_20780;
  wire [0:0] v_20781;
  function [0:0] mux_20781(input [0:0] sel);
    case (sel) 0: mux_20781 = 1'h0; 1: mux_20781 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20782;
  function [0:0] mux_20782(input [0:0] sel);
    case (sel) 0: mux_20782 = 1'h0; 1: mux_20782 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20783;
  wire [0:0] v_20784;
  wire [0:0] v_20785;
  wire [0:0] v_20786;
  wire [0:0] v_20787;
  wire [0:0] v_20788;
  wire [0:0] v_20789;
  function [0:0] mux_20789(input [0:0] sel);
    case (sel) 0: mux_20789 = 1'h0; 1: mux_20789 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20790;
  function [0:0] mux_20790(input [0:0] sel);
    case (sel) 0: mux_20790 = 1'h0; 1: mux_20790 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20791;
  wire [0:0] v_20792;
  wire [0:0] v_20793;
  wire [0:0] v_20794;
  function [0:0] mux_20794(input [0:0] sel);
    case (sel) 0: mux_20794 = 1'h0; 1: mux_20794 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20795;
  function [0:0] mux_20795(input [0:0] sel);
    case (sel) 0: mux_20795 = 1'h0; 1: mux_20795 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20796;
  wire [0:0] v_20797;
  wire [0:0] v_20798;
  wire [0:0] v_20799;
  wire [0:0] v_20800;
  wire [0:0] v_20801;
  function [0:0] mux_20801(input [0:0] sel);
    case (sel) 0: mux_20801 = 1'h0; 1: mux_20801 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20802;
  wire [0:0] v_20803;
  wire [0:0] v_20804;
  wire [0:0] v_20805;
  wire [0:0] v_20806;
  function [0:0] mux_20806(input [0:0] sel);
    case (sel) 0: mux_20806 = 1'h0; 1: mux_20806 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20807;
  wire [0:0] v_20808;
  wire [0:0] v_20809;
  wire [0:0] v_20810;
  function [0:0] mux_20810(input [0:0] sel);
    case (sel) 0: mux_20810 = 1'h0; 1: mux_20810 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20811;
  function [0:0] mux_20811(input [0:0] sel);
    case (sel) 0: mux_20811 = 1'h0; 1: mux_20811 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_20812 = 1'h0;
  wire [0:0] v_20813;
  wire [0:0] v_20814;
  wire [0:0] act_20815;
  wire [0:0] v_20816;
  wire [0:0] v_20817;
  wire [0:0] v_20818;
  reg [0:0] v_20819 = 1'h0;
  wire [0:0] v_20820;
  wire [0:0] v_20821;
  wire [0:0] act_20822;
  wire [0:0] v_20823;
  wire [0:0] v_20824;
  wire [0:0] v_20825;
  wire [0:0] vin0_consume_en_20826;
  wire [0:0] vout_canPeek_20826;
  wire [7:0] vout_peek_20826;
  wire [0:0] v_20827;
  wire [0:0] v_20828;
  function [0:0] mux_20828(input [0:0] sel);
    case (sel) 0: mux_20828 = 1'h0; 1: mux_20828 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20829;
  wire [0:0] v_20830;
  wire [0:0] v_20831;
  wire [0:0] v_20832;
  wire [0:0] v_20833;
  function [0:0] mux_20833(input [0:0] sel);
    case (sel) 0: mux_20833 = 1'h0; 1: mux_20833 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20834;
  wire [0:0] vin0_consume_en_20835;
  wire [0:0] vout_canPeek_20835;
  wire [7:0] vout_peek_20835;
  wire [0:0] v_20836;
  wire [0:0] v_20837;
  function [0:0] mux_20837(input [0:0] sel);
    case (sel) 0: mux_20837 = 1'h0; 1: mux_20837 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20838;
  function [0:0] mux_20838(input [0:0] sel);
    case (sel) 0: mux_20838 = 1'h0; 1: mux_20838 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20839;
  wire [0:0] v_20840;
  wire [0:0] v_20841;
  wire [0:0] v_20842;
  wire [0:0] v_20843;
  wire [0:0] v_20844;
  wire [0:0] v_20845;
  function [0:0] mux_20845(input [0:0] sel);
    case (sel) 0: mux_20845 = 1'h0; 1: mux_20845 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20846;
  wire [0:0] v_20847;
  wire [0:0] v_20848;
  wire [0:0] v_20849;
  wire [0:0] v_20850;
  function [0:0] mux_20850(input [0:0] sel);
    case (sel) 0: mux_20850 = 1'h0; 1: mux_20850 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20851;
  wire [0:0] v_20852;
  wire [0:0] v_20853;
  wire [0:0] v_20854;
  function [0:0] mux_20854(input [0:0] sel);
    case (sel) 0: mux_20854 = 1'h0; 1: mux_20854 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20855;
  function [0:0] mux_20855(input [0:0] sel);
    case (sel) 0: mux_20855 = 1'h0; 1: mux_20855 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_20856 = 1'h0;
  wire [0:0] v_20857;
  wire [0:0] v_20858;
  wire [0:0] act_20859;
  wire [0:0] v_20860;
  wire [0:0] v_20861;
  wire [0:0] v_20862;
  wire [0:0] vin0_consume_en_20863;
  wire [0:0] vout_canPeek_20863;
  wire [7:0] vout_peek_20863;
  wire [0:0] v_20864;
  wire [0:0] v_20865;
  function [0:0] mux_20865(input [0:0] sel);
    case (sel) 0: mux_20865 = 1'h0; 1: mux_20865 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20866;
  wire [0:0] v_20867;
  wire [0:0] v_20868;
  wire [0:0] v_20869;
  wire [0:0] v_20870;
  function [0:0] mux_20870(input [0:0] sel);
    case (sel) 0: mux_20870 = 1'h0; 1: mux_20870 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20871;
  wire [0:0] vin0_consume_en_20872;
  wire [0:0] vout_canPeek_20872;
  wire [7:0] vout_peek_20872;
  wire [0:0] v_20873;
  wire [0:0] v_20874;
  function [0:0] mux_20874(input [0:0] sel);
    case (sel) 0: mux_20874 = 1'h0; 1: mux_20874 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20875;
  function [0:0] mux_20875(input [0:0] sel);
    case (sel) 0: mux_20875 = 1'h0; 1: mux_20875 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20876;
  wire [0:0] v_20877;
  wire [0:0] v_20878;
  wire [0:0] v_20879;
  wire [0:0] v_20880;
  wire [0:0] v_20881;
  wire [0:0] v_20882;
  function [0:0] mux_20882(input [0:0] sel);
    case (sel) 0: mux_20882 = 1'h0; 1: mux_20882 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20883;
  function [0:0] mux_20883(input [0:0] sel);
    case (sel) 0: mux_20883 = 1'h0; 1: mux_20883 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20884;
  wire [0:0] v_20885;
  wire [0:0] v_20886;
  wire [0:0] v_20887;
  function [0:0] mux_20887(input [0:0] sel);
    case (sel) 0: mux_20887 = 1'h0; 1: mux_20887 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20888;
  function [0:0] mux_20888(input [0:0] sel);
    case (sel) 0: mux_20888 = 1'h0; 1: mux_20888 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20889;
  wire [0:0] v_20890;
  wire [0:0] v_20891;
  wire [0:0] v_20892;
  wire [0:0] v_20893;
  wire [0:0] v_20894;
  function [0:0] mux_20894(input [0:0] sel);
    case (sel) 0: mux_20894 = 1'h0; 1: mux_20894 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20895;
  function [0:0] mux_20895(input [0:0] sel);
    case (sel) 0: mux_20895 = 1'h0; 1: mux_20895 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20896;
  wire [0:0] v_20897;
  wire [0:0] v_20898;
  wire [0:0] v_20899;
  function [0:0] mux_20899(input [0:0] sel);
    case (sel) 0: mux_20899 = 1'h0; 1: mux_20899 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20900;
  function [0:0] mux_20900(input [0:0] sel);
    case (sel) 0: mux_20900 = 1'h0; 1: mux_20900 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20901;
  wire [0:0] v_20902;
  wire [0:0] v_20903;
  wire [0:0] v_20904;
  wire [0:0] v_20905;
  wire [0:0] v_20906;
  function [0:0] mux_20906(input [0:0] sel);
    case (sel) 0: mux_20906 = 1'h0; 1: mux_20906 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20907;
  function [0:0] mux_20907(input [0:0] sel);
    case (sel) 0: mux_20907 = 1'h0; 1: mux_20907 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20908;
  wire [0:0] v_20909;
  wire [0:0] v_20910;
  wire [0:0] v_20911;
  function [0:0] mux_20911(input [0:0] sel);
    case (sel) 0: mux_20911 = 1'h0; 1: mux_20911 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20912;
  function [0:0] mux_20912(input [0:0] sel);
    case (sel) 0: mux_20912 = 1'h0; 1: mux_20912 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20913;
  wire [0:0] v_20914;
  wire [0:0] v_20915;
  wire [0:0] v_20916;
  wire [0:0] v_20917;
  wire [0:0] v_20918;
  function [0:0] mux_20918(input [0:0] sel);
    case (sel) 0: mux_20918 = 1'h0; 1: mux_20918 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20919;
  wire [0:0] v_20920;
  wire [0:0] v_20921;
  wire [0:0] v_20922;
  wire [0:0] v_20923;
  function [0:0] mux_20923(input [0:0] sel);
    case (sel) 0: mux_20923 = 1'h0; 1: mux_20923 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20924;
  wire [0:0] v_20925;
  wire [0:0] v_20926;
  wire [0:0] v_20927;
  function [0:0] mux_20927(input [0:0] sel);
    case (sel) 0: mux_20927 = 1'h0; 1: mux_20927 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20928;
  function [0:0] mux_20928(input [0:0] sel);
    case (sel) 0: mux_20928 = 1'h0; 1: mux_20928 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_20929 = 1'h0;
  wire [0:0] v_20930;
  wire [0:0] v_20931;
  wire [0:0] act_20932;
  wire [0:0] v_20933;
  wire [0:0] v_20934;
  wire [0:0] v_20935;
  reg [0:0] v_20936 = 1'h0;
  wire [0:0] v_20937;
  wire [0:0] v_20938;
  wire [0:0] act_20939;
  wire [0:0] v_20940;
  wire [0:0] v_20941;
  wire [0:0] v_20942;
  reg [0:0] v_20943 = 1'h0;
  wire [0:0] v_20944;
  wire [0:0] v_20945;
  wire [0:0] act_20946;
  wire [0:0] v_20947;
  wire [0:0] v_20948;
  wire [0:0] v_20949;
  reg [0:0] v_20950 = 1'h0;
  wire [0:0] v_20951;
  wire [0:0] v_20952;
  wire [0:0] act_20953;
  wire [0:0] v_20954;
  wire [0:0] v_20955;
  wire [0:0] v_20956;
  wire [0:0] vin0_consume_en_20957;
  wire [0:0] vout_canPeek_20957;
  wire [7:0] vout_peek_20957;
  wire [0:0] v_20958;
  wire [0:0] v_20959;
  function [0:0] mux_20959(input [0:0] sel);
    case (sel) 0: mux_20959 = 1'h0; 1: mux_20959 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20960;
  wire [0:0] v_20961;
  wire [0:0] v_20962;
  wire [0:0] v_20963;
  wire [0:0] v_20964;
  function [0:0] mux_20964(input [0:0] sel);
    case (sel) 0: mux_20964 = 1'h0; 1: mux_20964 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20965;
  wire [0:0] vin0_consume_en_20966;
  wire [0:0] vout_canPeek_20966;
  wire [7:0] vout_peek_20966;
  wire [0:0] v_20967;
  wire [0:0] v_20968;
  function [0:0] mux_20968(input [0:0] sel);
    case (sel) 0: mux_20968 = 1'h0; 1: mux_20968 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20969;
  function [0:0] mux_20969(input [0:0] sel);
    case (sel) 0: mux_20969 = 1'h0; 1: mux_20969 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20970;
  wire [0:0] v_20971;
  wire [0:0] v_20972;
  wire [0:0] v_20973;
  wire [0:0] v_20974;
  wire [0:0] v_20975;
  wire [0:0] v_20976;
  function [0:0] mux_20976(input [0:0] sel);
    case (sel) 0: mux_20976 = 1'h0; 1: mux_20976 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20977;
  wire [0:0] v_20978;
  wire [0:0] v_20979;
  wire [0:0] v_20980;
  wire [0:0] v_20981;
  function [0:0] mux_20981(input [0:0] sel);
    case (sel) 0: mux_20981 = 1'h0; 1: mux_20981 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_20982;
  wire [0:0] v_20983;
  wire [0:0] v_20984;
  wire [0:0] v_20985;
  function [0:0] mux_20985(input [0:0] sel);
    case (sel) 0: mux_20985 = 1'h0; 1: mux_20985 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20986;
  function [0:0] mux_20986(input [0:0] sel);
    case (sel) 0: mux_20986 = 1'h0; 1: mux_20986 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_20987 = 1'h0;
  wire [0:0] v_20988;
  wire [0:0] v_20989;
  wire [0:0] act_20990;
  wire [0:0] v_20991;
  wire [0:0] v_20992;
  wire [0:0] v_20993;
  wire [0:0] vin0_consume_en_20994;
  wire [0:0] vout_canPeek_20994;
  wire [7:0] vout_peek_20994;
  wire [0:0] v_20995;
  wire [0:0] v_20996;
  function [0:0] mux_20996(input [0:0] sel);
    case (sel) 0: mux_20996 = 1'h0; 1: mux_20996 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_20997;
  wire [0:0] v_20998;
  wire [0:0] v_20999;
  wire [0:0] v_21000;
  wire [0:0] v_21001;
  function [0:0] mux_21001(input [0:0] sel);
    case (sel) 0: mux_21001 = 1'h0; 1: mux_21001 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21002;
  wire [0:0] vin0_consume_en_21003;
  wire [0:0] vout_canPeek_21003;
  wire [7:0] vout_peek_21003;
  wire [0:0] v_21004;
  wire [0:0] v_21005;
  function [0:0] mux_21005(input [0:0] sel);
    case (sel) 0: mux_21005 = 1'h0; 1: mux_21005 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21006;
  function [0:0] mux_21006(input [0:0] sel);
    case (sel) 0: mux_21006 = 1'h0; 1: mux_21006 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21007;
  wire [0:0] v_21008;
  wire [0:0] v_21009;
  wire [0:0] v_21010;
  wire [0:0] v_21011;
  wire [0:0] v_21012;
  wire [0:0] v_21013;
  function [0:0] mux_21013(input [0:0] sel);
    case (sel) 0: mux_21013 = 1'h0; 1: mux_21013 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21014;
  function [0:0] mux_21014(input [0:0] sel);
    case (sel) 0: mux_21014 = 1'h0; 1: mux_21014 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21015;
  wire [0:0] v_21016;
  wire [0:0] v_21017;
  wire [0:0] v_21018;
  function [0:0] mux_21018(input [0:0] sel);
    case (sel) 0: mux_21018 = 1'h0; 1: mux_21018 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21019;
  function [0:0] mux_21019(input [0:0] sel);
    case (sel) 0: mux_21019 = 1'h0; 1: mux_21019 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21020;
  wire [0:0] v_21021;
  wire [0:0] v_21022;
  wire [0:0] v_21023;
  wire [0:0] v_21024;
  wire [0:0] v_21025;
  function [0:0] mux_21025(input [0:0] sel);
    case (sel) 0: mux_21025 = 1'h0; 1: mux_21025 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21026;
  wire [0:0] v_21027;
  wire [0:0] v_21028;
  wire [0:0] v_21029;
  wire [0:0] v_21030;
  function [0:0] mux_21030(input [0:0] sel);
    case (sel) 0: mux_21030 = 1'h0; 1: mux_21030 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21031;
  wire [0:0] v_21032;
  wire [0:0] v_21033;
  wire [0:0] v_21034;
  function [0:0] mux_21034(input [0:0] sel);
    case (sel) 0: mux_21034 = 1'h0; 1: mux_21034 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21035;
  function [0:0] mux_21035(input [0:0] sel);
    case (sel) 0: mux_21035 = 1'h0; 1: mux_21035 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_21036 = 1'h0;
  wire [0:0] v_21037;
  wire [0:0] v_21038;
  wire [0:0] act_21039;
  wire [0:0] v_21040;
  wire [0:0] v_21041;
  wire [0:0] v_21042;
  reg [0:0] v_21043 = 1'h0;
  wire [0:0] v_21044;
  wire [0:0] v_21045;
  wire [0:0] act_21046;
  wire [0:0] v_21047;
  wire [0:0] v_21048;
  wire [0:0] v_21049;
  wire [0:0] vin0_consume_en_21050;
  wire [0:0] vout_canPeek_21050;
  wire [7:0] vout_peek_21050;
  wire [0:0] v_21051;
  wire [0:0] v_21052;
  function [0:0] mux_21052(input [0:0] sel);
    case (sel) 0: mux_21052 = 1'h0; 1: mux_21052 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21053;
  wire [0:0] v_21054;
  wire [0:0] v_21055;
  wire [0:0] v_21056;
  wire [0:0] v_21057;
  function [0:0] mux_21057(input [0:0] sel);
    case (sel) 0: mux_21057 = 1'h0; 1: mux_21057 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21058;
  wire [0:0] vin0_consume_en_21059;
  wire [0:0] vout_canPeek_21059;
  wire [7:0] vout_peek_21059;
  wire [0:0] v_21060;
  wire [0:0] v_21061;
  function [0:0] mux_21061(input [0:0] sel);
    case (sel) 0: mux_21061 = 1'h0; 1: mux_21061 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21062;
  function [0:0] mux_21062(input [0:0] sel);
    case (sel) 0: mux_21062 = 1'h0; 1: mux_21062 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21063;
  wire [0:0] v_21064;
  wire [0:0] v_21065;
  wire [0:0] v_21066;
  wire [0:0] v_21067;
  wire [0:0] v_21068;
  wire [0:0] v_21069;
  function [0:0] mux_21069(input [0:0] sel);
    case (sel) 0: mux_21069 = 1'h0; 1: mux_21069 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21070;
  wire [0:0] v_21071;
  wire [0:0] v_21072;
  wire [0:0] v_21073;
  wire [0:0] v_21074;
  function [0:0] mux_21074(input [0:0] sel);
    case (sel) 0: mux_21074 = 1'h0; 1: mux_21074 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21075;
  wire [0:0] v_21076;
  wire [0:0] v_21077;
  wire [0:0] v_21078;
  function [0:0] mux_21078(input [0:0] sel);
    case (sel) 0: mux_21078 = 1'h0; 1: mux_21078 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21079;
  function [0:0] mux_21079(input [0:0] sel);
    case (sel) 0: mux_21079 = 1'h0; 1: mux_21079 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_21080 = 1'h0;
  wire [0:0] v_21081;
  wire [0:0] v_21082;
  wire [0:0] act_21083;
  wire [0:0] v_21084;
  wire [0:0] v_21085;
  wire [0:0] v_21086;
  wire [0:0] vin0_consume_en_21087;
  wire [0:0] vout_canPeek_21087;
  wire [7:0] vout_peek_21087;
  wire [0:0] v_21088;
  wire [0:0] v_21089;
  function [0:0] mux_21089(input [0:0] sel);
    case (sel) 0: mux_21089 = 1'h0; 1: mux_21089 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21090;
  wire [0:0] v_21091;
  wire [0:0] v_21092;
  wire [0:0] v_21093;
  wire [0:0] v_21094;
  function [0:0] mux_21094(input [0:0] sel);
    case (sel) 0: mux_21094 = 1'h0; 1: mux_21094 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21095;
  wire [0:0] vin0_consume_en_21096;
  wire [0:0] vout_canPeek_21096;
  wire [7:0] vout_peek_21096;
  wire [0:0] v_21097;
  wire [0:0] v_21098;
  function [0:0] mux_21098(input [0:0] sel);
    case (sel) 0: mux_21098 = 1'h0; 1: mux_21098 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21099;
  function [0:0] mux_21099(input [0:0] sel);
    case (sel) 0: mux_21099 = 1'h0; 1: mux_21099 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21100;
  wire [0:0] v_21101;
  wire [0:0] v_21102;
  wire [0:0] v_21103;
  wire [0:0] v_21104;
  wire [0:0] v_21105;
  wire [0:0] v_21106;
  function [0:0] mux_21106(input [0:0] sel);
    case (sel) 0: mux_21106 = 1'h0; 1: mux_21106 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21107;
  function [0:0] mux_21107(input [0:0] sel);
    case (sel) 0: mux_21107 = 1'h0; 1: mux_21107 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21108;
  wire [0:0] v_21109;
  wire [0:0] v_21110;
  wire [0:0] v_21111;
  function [0:0] mux_21111(input [0:0] sel);
    case (sel) 0: mux_21111 = 1'h0; 1: mux_21111 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21112;
  function [0:0] mux_21112(input [0:0] sel);
    case (sel) 0: mux_21112 = 1'h0; 1: mux_21112 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21113;
  wire [0:0] v_21114;
  wire [0:0] v_21115;
  wire [0:0] v_21116;
  wire [0:0] v_21117;
  wire [0:0] v_21118;
  function [0:0] mux_21118(input [0:0] sel);
    case (sel) 0: mux_21118 = 1'h0; 1: mux_21118 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21119;
  function [0:0] mux_21119(input [0:0] sel);
    case (sel) 0: mux_21119 = 1'h0; 1: mux_21119 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21120;
  wire [0:0] v_21121;
  wire [0:0] v_21122;
  wire [0:0] v_21123;
  function [0:0] mux_21123(input [0:0] sel);
    case (sel) 0: mux_21123 = 1'h0; 1: mux_21123 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21124;
  function [0:0] mux_21124(input [0:0] sel);
    case (sel) 0: mux_21124 = 1'h0; 1: mux_21124 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21125;
  wire [0:0] v_21126;
  wire [0:0] v_21127;
  wire [0:0] v_21128;
  wire [0:0] v_21129;
  wire [0:0] v_21130;
  function [0:0] mux_21130(input [0:0] sel);
    case (sel) 0: mux_21130 = 1'h0; 1: mux_21130 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21131;
  wire [0:0] v_21132;
  wire [0:0] v_21133;
  wire [0:0] v_21134;
  wire [0:0] v_21135;
  function [0:0] mux_21135(input [0:0] sel);
    case (sel) 0: mux_21135 = 1'h0; 1: mux_21135 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21136;
  wire [0:0] v_21137;
  wire [0:0] v_21138;
  wire [0:0] v_21139;
  function [0:0] mux_21139(input [0:0] sel);
    case (sel) 0: mux_21139 = 1'h0; 1: mux_21139 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21140;
  function [0:0] mux_21140(input [0:0] sel);
    case (sel) 0: mux_21140 = 1'h0; 1: mux_21140 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_21141 = 1'h0;
  wire [0:0] v_21142;
  wire [0:0] v_21143;
  wire [0:0] act_21144;
  wire [0:0] v_21145;
  wire [0:0] v_21146;
  wire [0:0] v_21147;
  reg [0:0] v_21148 = 1'h0;
  wire [0:0] v_21149;
  wire [0:0] v_21150;
  wire [0:0] act_21151;
  wire [0:0] v_21152;
  wire [0:0] v_21153;
  wire [0:0] v_21154;
  reg [0:0] v_21155 = 1'h0;
  wire [0:0] v_21156;
  wire [0:0] v_21157;
  wire [0:0] act_21158;
  wire [0:0] v_21159;
  wire [0:0] v_21160;
  wire [0:0] v_21161;
  wire [0:0] vin0_consume_en_21162;
  wire [0:0] vout_canPeek_21162;
  wire [7:0] vout_peek_21162;
  wire [0:0] v_21163;
  wire [0:0] v_21164;
  function [0:0] mux_21164(input [0:0] sel);
    case (sel) 0: mux_21164 = 1'h0; 1: mux_21164 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21165;
  wire [0:0] v_21166;
  wire [0:0] v_21167;
  wire [0:0] v_21168;
  wire [0:0] v_21169;
  function [0:0] mux_21169(input [0:0] sel);
    case (sel) 0: mux_21169 = 1'h0; 1: mux_21169 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21170;
  wire [0:0] vin0_consume_en_21171;
  wire [0:0] vout_canPeek_21171;
  wire [7:0] vout_peek_21171;
  wire [0:0] v_21172;
  wire [0:0] v_21173;
  function [0:0] mux_21173(input [0:0] sel);
    case (sel) 0: mux_21173 = 1'h0; 1: mux_21173 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21174;
  function [0:0] mux_21174(input [0:0] sel);
    case (sel) 0: mux_21174 = 1'h0; 1: mux_21174 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21175;
  wire [0:0] v_21176;
  wire [0:0] v_21177;
  wire [0:0] v_21178;
  wire [0:0] v_21179;
  wire [0:0] v_21180;
  wire [0:0] v_21181;
  function [0:0] mux_21181(input [0:0] sel);
    case (sel) 0: mux_21181 = 1'h0; 1: mux_21181 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21182;
  wire [0:0] v_21183;
  wire [0:0] v_21184;
  wire [0:0] v_21185;
  wire [0:0] v_21186;
  function [0:0] mux_21186(input [0:0] sel);
    case (sel) 0: mux_21186 = 1'h0; 1: mux_21186 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21187;
  wire [0:0] v_21188;
  wire [0:0] v_21189;
  wire [0:0] v_21190;
  function [0:0] mux_21190(input [0:0] sel);
    case (sel) 0: mux_21190 = 1'h0; 1: mux_21190 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21191;
  function [0:0] mux_21191(input [0:0] sel);
    case (sel) 0: mux_21191 = 1'h0; 1: mux_21191 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_21192 = 1'h0;
  wire [0:0] v_21193;
  wire [0:0] v_21194;
  wire [0:0] act_21195;
  wire [0:0] v_21196;
  wire [0:0] v_21197;
  wire [0:0] v_21198;
  wire [0:0] vin0_consume_en_21199;
  wire [0:0] vout_canPeek_21199;
  wire [7:0] vout_peek_21199;
  wire [0:0] v_21200;
  wire [0:0] v_21201;
  function [0:0] mux_21201(input [0:0] sel);
    case (sel) 0: mux_21201 = 1'h0; 1: mux_21201 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21202;
  wire [0:0] v_21203;
  wire [0:0] v_21204;
  wire [0:0] v_21205;
  wire [0:0] v_21206;
  function [0:0] mux_21206(input [0:0] sel);
    case (sel) 0: mux_21206 = 1'h0; 1: mux_21206 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21207;
  wire [0:0] vin0_consume_en_21208;
  wire [0:0] vout_canPeek_21208;
  wire [7:0] vout_peek_21208;
  wire [0:0] v_21209;
  wire [0:0] v_21210;
  function [0:0] mux_21210(input [0:0] sel);
    case (sel) 0: mux_21210 = 1'h0; 1: mux_21210 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21211;
  function [0:0] mux_21211(input [0:0] sel);
    case (sel) 0: mux_21211 = 1'h0; 1: mux_21211 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21212;
  wire [0:0] v_21213;
  wire [0:0] v_21214;
  wire [0:0] v_21215;
  wire [0:0] v_21216;
  wire [0:0] v_21217;
  wire [0:0] v_21218;
  function [0:0] mux_21218(input [0:0] sel);
    case (sel) 0: mux_21218 = 1'h0; 1: mux_21218 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21219;
  function [0:0] mux_21219(input [0:0] sel);
    case (sel) 0: mux_21219 = 1'h0; 1: mux_21219 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21220;
  wire [0:0] v_21221;
  wire [0:0] v_21222;
  wire [0:0] v_21223;
  function [0:0] mux_21223(input [0:0] sel);
    case (sel) 0: mux_21223 = 1'h0; 1: mux_21223 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21224;
  function [0:0] mux_21224(input [0:0] sel);
    case (sel) 0: mux_21224 = 1'h0; 1: mux_21224 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21225;
  wire [0:0] v_21226;
  wire [0:0] v_21227;
  wire [0:0] v_21228;
  wire [0:0] v_21229;
  wire [0:0] v_21230;
  function [0:0] mux_21230(input [0:0] sel);
    case (sel) 0: mux_21230 = 1'h0; 1: mux_21230 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21231;
  wire [0:0] v_21232;
  wire [0:0] v_21233;
  wire [0:0] v_21234;
  wire [0:0] v_21235;
  function [0:0] mux_21235(input [0:0] sel);
    case (sel) 0: mux_21235 = 1'h0; 1: mux_21235 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21236;
  wire [0:0] v_21237;
  wire [0:0] v_21238;
  wire [0:0] v_21239;
  function [0:0] mux_21239(input [0:0] sel);
    case (sel) 0: mux_21239 = 1'h0; 1: mux_21239 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21240;
  function [0:0] mux_21240(input [0:0] sel);
    case (sel) 0: mux_21240 = 1'h0; 1: mux_21240 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_21241 = 1'h0;
  wire [0:0] v_21242;
  wire [0:0] v_21243;
  wire [0:0] act_21244;
  wire [0:0] v_21245;
  wire [0:0] v_21246;
  wire [0:0] v_21247;
  reg [0:0] v_21248 = 1'h0;
  wire [0:0] v_21249;
  wire [0:0] v_21250;
  wire [0:0] act_21251;
  wire [0:0] v_21252;
  wire [0:0] v_21253;
  wire [0:0] v_21254;
  wire [0:0] vin0_consume_en_21255;
  wire [0:0] vout_canPeek_21255;
  wire [7:0] vout_peek_21255;
  wire [0:0] v_21256;
  wire [0:0] v_21257;
  function [0:0] mux_21257(input [0:0] sel);
    case (sel) 0: mux_21257 = 1'h0; 1: mux_21257 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21258;
  wire [0:0] v_21259;
  wire [0:0] v_21260;
  wire [0:0] v_21261;
  wire [0:0] v_21262;
  function [0:0] mux_21262(input [0:0] sel);
    case (sel) 0: mux_21262 = 1'h0; 1: mux_21262 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21263;
  wire [0:0] vin0_consume_en_21264;
  wire [0:0] vout_canPeek_21264;
  wire [7:0] vout_peek_21264;
  wire [0:0] v_21265;
  wire [0:0] v_21266;
  function [0:0] mux_21266(input [0:0] sel);
    case (sel) 0: mux_21266 = 1'h0; 1: mux_21266 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21267;
  function [0:0] mux_21267(input [0:0] sel);
    case (sel) 0: mux_21267 = 1'h0; 1: mux_21267 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21268;
  wire [0:0] v_21269;
  wire [0:0] v_21270;
  wire [0:0] v_21271;
  wire [0:0] v_21272;
  wire [0:0] v_21273;
  wire [0:0] v_21274;
  function [0:0] mux_21274(input [0:0] sel);
    case (sel) 0: mux_21274 = 1'h0; 1: mux_21274 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21275;
  wire [0:0] v_21276;
  wire [0:0] v_21277;
  wire [0:0] v_21278;
  wire [0:0] v_21279;
  function [0:0] mux_21279(input [0:0] sel);
    case (sel) 0: mux_21279 = 1'h0; 1: mux_21279 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21280;
  wire [0:0] v_21281;
  wire [0:0] v_21282;
  wire [0:0] v_21283;
  function [0:0] mux_21283(input [0:0] sel);
    case (sel) 0: mux_21283 = 1'h0; 1: mux_21283 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21284;
  function [0:0] mux_21284(input [0:0] sel);
    case (sel) 0: mux_21284 = 1'h0; 1: mux_21284 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_21285 = 1'h0;
  wire [0:0] v_21286;
  wire [0:0] v_21287;
  wire [0:0] act_21288;
  wire [0:0] v_21289;
  wire [0:0] v_21290;
  wire [0:0] v_21291;
  wire [0:0] vin0_consume_en_21292;
  wire [0:0] vout_canPeek_21292;
  wire [7:0] vout_peek_21292;
  wire [0:0] v_21293;
  wire [0:0] v_21294;
  function [0:0] mux_21294(input [0:0] sel);
    case (sel) 0: mux_21294 = 1'h0; 1: mux_21294 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21295;
  wire [0:0] v_21296;
  wire [0:0] v_21297;
  wire [0:0] v_21298;
  wire [0:0] v_21299;
  function [0:0] mux_21299(input [0:0] sel);
    case (sel) 0: mux_21299 = 1'h0; 1: mux_21299 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21300;
  wire [0:0] vin0_consume_en_21301;
  wire [0:0] vout_canPeek_21301;
  wire [7:0] vout_peek_21301;
  wire [0:0] v_21302;
  wire [0:0] v_21303;
  function [0:0] mux_21303(input [0:0] sel);
    case (sel) 0: mux_21303 = 1'h0; 1: mux_21303 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21304;
  function [0:0] mux_21304(input [0:0] sel);
    case (sel) 0: mux_21304 = 1'h0; 1: mux_21304 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21305;
  wire [0:0] v_21306;
  wire [0:0] v_21307;
  wire [0:0] v_21308;
  wire [0:0] v_21309;
  wire [0:0] v_21310;
  wire [0:0] v_21311;
  function [0:0] mux_21311(input [0:0] sel);
    case (sel) 0: mux_21311 = 1'h0; 1: mux_21311 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21312;
  function [0:0] mux_21312(input [0:0] sel);
    case (sel) 0: mux_21312 = 1'h0; 1: mux_21312 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21313;
  wire [0:0] v_21314;
  wire [0:0] v_21315;
  wire [0:0] v_21316;
  function [0:0] mux_21316(input [0:0] sel);
    case (sel) 0: mux_21316 = 1'h0; 1: mux_21316 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21317;
  function [0:0] mux_21317(input [0:0] sel);
    case (sel) 0: mux_21317 = 1'h0; 1: mux_21317 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21318;
  wire [0:0] v_21319;
  wire [0:0] v_21320;
  wire [0:0] v_21321;
  wire [0:0] v_21322;
  wire [0:0] v_21323;
  function [0:0] mux_21323(input [0:0] sel);
    case (sel) 0: mux_21323 = 1'h0; 1: mux_21323 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21324;
  function [0:0] mux_21324(input [0:0] sel);
    case (sel) 0: mux_21324 = 1'h0; 1: mux_21324 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21325;
  wire [0:0] v_21326;
  wire [0:0] v_21327;
  wire [0:0] v_21328;
  function [0:0] mux_21328(input [0:0] sel);
    case (sel) 0: mux_21328 = 1'h0; 1: mux_21328 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21329;
  function [0:0] mux_21329(input [0:0] sel);
    case (sel) 0: mux_21329 = 1'h0; 1: mux_21329 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21330;
  wire [0:0] v_21331;
  wire [0:0] v_21332;
  wire [0:0] v_21333;
  wire [0:0] v_21334;
  wire [0:0] v_21335;
  function [0:0] mux_21335(input [0:0] sel);
    case (sel) 0: mux_21335 = 1'h0; 1: mux_21335 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21336;
  function [0:0] mux_21336(input [0:0] sel);
    case (sel) 0: mux_21336 = 1'h0; 1: mux_21336 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21337;
  wire [0:0] v_21338;
  wire [0:0] v_21339;
  wire [0:0] v_21340;
  function [0:0] mux_21340(input [0:0] sel);
    case (sel) 0: mux_21340 = 1'h0; 1: mux_21340 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21341;
  function [0:0] mux_21341(input [0:0] sel);
    case (sel) 0: mux_21341 = 1'h0; 1: mux_21341 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21342;
  wire [0:0] v_21343;
  wire [0:0] v_21344;
  wire [0:0] v_21345;
  wire [0:0] v_21346;
  wire [0:0] v_21347;
  function [0:0] mux_21347(input [0:0] sel);
    case (sel) 0: mux_21347 = 1'h0; 1: mux_21347 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21348;
  function [0:0] mux_21348(input [0:0] sel);
    case (sel) 0: mux_21348 = 1'h0; 1: mux_21348 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21349;
  wire [0:0] v_21350;
  wire [0:0] v_21351;
  wire [0:0] v_21352;
  function [0:0] mux_21352(input [0:0] sel);
    case (sel) 0: mux_21352 = 1'h0; 1: mux_21352 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21353;
  function [0:0] mux_21353(input [0:0] sel);
    case (sel) 0: mux_21353 = 1'h0; 1: mux_21353 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21354;
  wire [0:0] v_21355;
  wire [0:0] v_21356;
  wire [0:0] v_21357;
  wire [0:0] v_21358;
  wire [0:0] v_21359;
  function [0:0] mux_21359(input [0:0] sel);
    case (sel) 0: mux_21359 = 1'h0; 1: mux_21359 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21360;
  wire [0:0] v_21361;
  wire [0:0] v_21362;
  wire [0:0] v_21363;
  wire [0:0] v_21364;
  function [0:0] mux_21364(input [0:0] sel);
    case (sel) 0: mux_21364 = 1'h0; 1: mux_21364 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21365;
  wire [0:0] v_21366;
  wire [0:0] v_21367;
  wire [0:0] v_21368;
  function [0:0] mux_21368(input [0:0] sel);
    case (sel) 0: mux_21368 = 1'h0; 1: mux_21368 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21369;
  function [0:0] mux_21369(input [0:0] sel);
    case (sel) 0: mux_21369 = 1'h0; 1: mux_21369 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_21370 = 1'h0;
  wire [0:0] v_21371;
  wire [0:0] v_21372;
  wire [0:0] act_21373;
  wire [0:0] v_21374;
  wire [0:0] v_21375;
  wire [0:0] v_21376;
  reg [0:0] v_21377 = 1'h0;
  wire [0:0] v_21378;
  wire [0:0] v_21379;
  wire [0:0] act_21380;
  wire [0:0] v_21381;
  wire [0:0] v_21382;
  wire [0:0] v_21383;
  reg [0:0] v_21384 = 1'h0;
  wire [0:0] v_21385;
  wire [0:0] v_21386;
  wire [0:0] act_21387;
  wire [0:0] v_21388;
  wire [0:0] v_21389;
  wire [0:0] v_21390;
  reg [0:0] v_21391 = 1'h0;
  wire [0:0] v_21392;
  wire [0:0] v_21393;
  wire [0:0] act_21394;
  wire [0:0] v_21395;
  wire [0:0] v_21396;
  wire [0:0] v_21397;
  reg [0:0] v_21398 = 1'h0;
  wire [0:0] v_21399;
  wire [0:0] v_21400;
  wire [0:0] act_21401;
  wire [0:0] v_21402;
  wire [0:0] v_21403;
  wire [0:0] v_21404;
  wire [0:0] vin0_consume_en_21405;
  wire [0:0] vout_canPeek_21405;
  wire [7:0] vout_peek_21405;
  wire [0:0] v_21406;
  wire [0:0] v_21407;
  function [0:0] mux_21407(input [0:0] sel);
    case (sel) 0: mux_21407 = 1'h0; 1: mux_21407 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21408;
  wire [0:0] v_21409;
  wire [0:0] v_21410;
  wire [0:0] v_21411;
  wire [0:0] v_21412;
  function [0:0] mux_21412(input [0:0] sel);
    case (sel) 0: mux_21412 = 1'h0; 1: mux_21412 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21413;
  wire [0:0] vin0_consume_en_21414;
  wire [0:0] vout_canPeek_21414;
  wire [7:0] vout_peek_21414;
  wire [0:0] v_21415;
  wire [0:0] v_21416;
  function [0:0] mux_21416(input [0:0] sel);
    case (sel) 0: mux_21416 = 1'h0; 1: mux_21416 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21417;
  function [0:0] mux_21417(input [0:0] sel);
    case (sel) 0: mux_21417 = 1'h0; 1: mux_21417 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21418;
  wire [0:0] v_21419;
  wire [0:0] v_21420;
  wire [0:0] v_21421;
  wire [0:0] v_21422;
  wire [0:0] v_21423;
  wire [0:0] v_21424;
  function [0:0] mux_21424(input [0:0] sel);
    case (sel) 0: mux_21424 = 1'h0; 1: mux_21424 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21425;
  wire [0:0] v_21426;
  wire [0:0] v_21427;
  wire [0:0] v_21428;
  wire [0:0] v_21429;
  function [0:0] mux_21429(input [0:0] sel);
    case (sel) 0: mux_21429 = 1'h0; 1: mux_21429 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21430;
  wire [0:0] v_21431;
  wire [0:0] v_21432;
  wire [0:0] v_21433;
  function [0:0] mux_21433(input [0:0] sel);
    case (sel) 0: mux_21433 = 1'h0; 1: mux_21433 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21434;
  function [0:0] mux_21434(input [0:0] sel);
    case (sel) 0: mux_21434 = 1'h0; 1: mux_21434 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_21435 = 1'h0;
  wire [0:0] v_21436;
  wire [0:0] v_21437;
  wire [0:0] act_21438;
  wire [0:0] v_21439;
  wire [0:0] v_21440;
  wire [0:0] v_21441;
  wire [0:0] vin0_consume_en_21442;
  wire [0:0] vout_canPeek_21442;
  wire [7:0] vout_peek_21442;
  wire [0:0] v_21443;
  wire [0:0] v_21444;
  function [0:0] mux_21444(input [0:0] sel);
    case (sel) 0: mux_21444 = 1'h0; 1: mux_21444 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21445;
  wire [0:0] v_21446;
  wire [0:0] v_21447;
  wire [0:0] v_21448;
  wire [0:0] v_21449;
  function [0:0] mux_21449(input [0:0] sel);
    case (sel) 0: mux_21449 = 1'h0; 1: mux_21449 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21450;
  wire [0:0] vin0_consume_en_21451;
  wire [0:0] vout_canPeek_21451;
  wire [7:0] vout_peek_21451;
  wire [0:0] v_21452;
  wire [0:0] v_21453;
  function [0:0] mux_21453(input [0:0] sel);
    case (sel) 0: mux_21453 = 1'h0; 1: mux_21453 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21454;
  function [0:0] mux_21454(input [0:0] sel);
    case (sel) 0: mux_21454 = 1'h0; 1: mux_21454 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21455;
  wire [0:0] v_21456;
  wire [0:0] v_21457;
  wire [0:0] v_21458;
  wire [0:0] v_21459;
  wire [0:0] v_21460;
  wire [0:0] v_21461;
  function [0:0] mux_21461(input [0:0] sel);
    case (sel) 0: mux_21461 = 1'h0; 1: mux_21461 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21462;
  function [0:0] mux_21462(input [0:0] sel);
    case (sel) 0: mux_21462 = 1'h0; 1: mux_21462 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21463;
  wire [0:0] v_21464;
  wire [0:0] v_21465;
  wire [0:0] v_21466;
  function [0:0] mux_21466(input [0:0] sel);
    case (sel) 0: mux_21466 = 1'h0; 1: mux_21466 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21467;
  function [0:0] mux_21467(input [0:0] sel);
    case (sel) 0: mux_21467 = 1'h0; 1: mux_21467 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21468;
  wire [0:0] v_21469;
  wire [0:0] v_21470;
  wire [0:0] v_21471;
  wire [0:0] v_21472;
  wire [0:0] v_21473;
  function [0:0] mux_21473(input [0:0] sel);
    case (sel) 0: mux_21473 = 1'h0; 1: mux_21473 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21474;
  wire [0:0] v_21475;
  wire [0:0] v_21476;
  wire [0:0] v_21477;
  wire [0:0] v_21478;
  function [0:0] mux_21478(input [0:0] sel);
    case (sel) 0: mux_21478 = 1'h0; 1: mux_21478 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21479;
  wire [0:0] v_21480;
  wire [0:0] v_21481;
  wire [0:0] v_21482;
  function [0:0] mux_21482(input [0:0] sel);
    case (sel) 0: mux_21482 = 1'h0; 1: mux_21482 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21483;
  function [0:0] mux_21483(input [0:0] sel);
    case (sel) 0: mux_21483 = 1'h0; 1: mux_21483 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_21484 = 1'h0;
  wire [0:0] v_21485;
  wire [0:0] v_21486;
  wire [0:0] act_21487;
  wire [0:0] v_21488;
  wire [0:0] v_21489;
  wire [0:0] v_21490;
  reg [0:0] v_21491 = 1'h0;
  wire [0:0] v_21492;
  wire [0:0] v_21493;
  wire [0:0] act_21494;
  wire [0:0] v_21495;
  wire [0:0] v_21496;
  wire [0:0] v_21497;
  wire [0:0] vin0_consume_en_21498;
  wire [0:0] vout_canPeek_21498;
  wire [7:0] vout_peek_21498;
  wire [0:0] v_21499;
  wire [0:0] v_21500;
  function [0:0] mux_21500(input [0:0] sel);
    case (sel) 0: mux_21500 = 1'h0; 1: mux_21500 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21501;
  wire [0:0] v_21502;
  wire [0:0] v_21503;
  wire [0:0] v_21504;
  wire [0:0] v_21505;
  function [0:0] mux_21505(input [0:0] sel);
    case (sel) 0: mux_21505 = 1'h0; 1: mux_21505 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21506;
  wire [0:0] vin0_consume_en_21507;
  wire [0:0] vout_canPeek_21507;
  wire [7:0] vout_peek_21507;
  wire [0:0] v_21508;
  wire [0:0] v_21509;
  function [0:0] mux_21509(input [0:0] sel);
    case (sel) 0: mux_21509 = 1'h0; 1: mux_21509 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21510;
  function [0:0] mux_21510(input [0:0] sel);
    case (sel) 0: mux_21510 = 1'h0; 1: mux_21510 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21511;
  wire [0:0] v_21512;
  wire [0:0] v_21513;
  wire [0:0] v_21514;
  wire [0:0] v_21515;
  wire [0:0] v_21516;
  wire [0:0] v_21517;
  function [0:0] mux_21517(input [0:0] sel);
    case (sel) 0: mux_21517 = 1'h0; 1: mux_21517 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21518;
  wire [0:0] v_21519;
  wire [0:0] v_21520;
  wire [0:0] v_21521;
  wire [0:0] v_21522;
  function [0:0] mux_21522(input [0:0] sel);
    case (sel) 0: mux_21522 = 1'h0; 1: mux_21522 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21523;
  wire [0:0] v_21524;
  wire [0:0] v_21525;
  wire [0:0] v_21526;
  function [0:0] mux_21526(input [0:0] sel);
    case (sel) 0: mux_21526 = 1'h0; 1: mux_21526 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21527;
  function [0:0] mux_21527(input [0:0] sel);
    case (sel) 0: mux_21527 = 1'h0; 1: mux_21527 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_21528 = 1'h0;
  wire [0:0] v_21529;
  wire [0:0] v_21530;
  wire [0:0] act_21531;
  wire [0:0] v_21532;
  wire [0:0] v_21533;
  wire [0:0] v_21534;
  wire [0:0] vin0_consume_en_21535;
  wire [0:0] vout_canPeek_21535;
  wire [7:0] vout_peek_21535;
  wire [0:0] v_21536;
  wire [0:0] v_21537;
  function [0:0] mux_21537(input [0:0] sel);
    case (sel) 0: mux_21537 = 1'h0; 1: mux_21537 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21538;
  wire [0:0] v_21539;
  wire [0:0] v_21540;
  wire [0:0] v_21541;
  wire [0:0] v_21542;
  function [0:0] mux_21542(input [0:0] sel);
    case (sel) 0: mux_21542 = 1'h0; 1: mux_21542 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21543;
  wire [0:0] vin0_consume_en_21544;
  wire [0:0] vout_canPeek_21544;
  wire [7:0] vout_peek_21544;
  wire [0:0] v_21545;
  wire [0:0] v_21546;
  function [0:0] mux_21546(input [0:0] sel);
    case (sel) 0: mux_21546 = 1'h0; 1: mux_21546 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21547;
  function [0:0] mux_21547(input [0:0] sel);
    case (sel) 0: mux_21547 = 1'h0; 1: mux_21547 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21548;
  wire [0:0] v_21549;
  wire [0:0] v_21550;
  wire [0:0] v_21551;
  wire [0:0] v_21552;
  wire [0:0] v_21553;
  wire [0:0] v_21554;
  function [0:0] mux_21554(input [0:0] sel);
    case (sel) 0: mux_21554 = 1'h0; 1: mux_21554 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21555;
  function [0:0] mux_21555(input [0:0] sel);
    case (sel) 0: mux_21555 = 1'h0; 1: mux_21555 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21556;
  wire [0:0] v_21557;
  wire [0:0] v_21558;
  wire [0:0] v_21559;
  function [0:0] mux_21559(input [0:0] sel);
    case (sel) 0: mux_21559 = 1'h0; 1: mux_21559 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21560;
  function [0:0] mux_21560(input [0:0] sel);
    case (sel) 0: mux_21560 = 1'h0; 1: mux_21560 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21561;
  wire [0:0] v_21562;
  wire [0:0] v_21563;
  wire [0:0] v_21564;
  wire [0:0] v_21565;
  wire [0:0] v_21566;
  function [0:0] mux_21566(input [0:0] sel);
    case (sel) 0: mux_21566 = 1'h0; 1: mux_21566 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21567;
  function [0:0] mux_21567(input [0:0] sel);
    case (sel) 0: mux_21567 = 1'h0; 1: mux_21567 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21568;
  wire [0:0] v_21569;
  wire [0:0] v_21570;
  wire [0:0] v_21571;
  function [0:0] mux_21571(input [0:0] sel);
    case (sel) 0: mux_21571 = 1'h0; 1: mux_21571 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21572;
  function [0:0] mux_21572(input [0:0] sel);
    case (sel) 0: mux_21572 = 1'h0; 1: mux_21572 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21573;
  wire [0:0] v_21574;
  wire [0:0] v_21575;
  wire [0:0] v_21576;
  wire [0:0] v_21577;
  wire [0:0] v_21578;
  function [0:0] mux_21578(input [0:0] sel);
    case (sel) 0: mux_21578 = 1'h0; 1: mux_21578 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21579;
  wire [0:0] v_21580;
  wire [0:0] v_21581;
  wire [0:0] v_21582;
  wire [0:0] v_21583;
  function [0:0] mux_21583(input [0:0] sel);
    case (sel) 0: mux_21583 = 1'h0; 1: mux_21583 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21584;
  wire [0:0] v_21585;
  wire [0:0] v_21586;
  wire [0:0] v_21587;
  function [0:0] mux_21587(input [0:0] sel);
    case (sel) 0: mux_21587 = 1'h0; 1: mux_21587 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21588;
  function [0:0] mux_21588(input [0:0] sel);
    case (sel) 0: mux_21588 = 1'h0; 1: mux_21588 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_21589 = 1'h0;
  wire [0:0] v_21590;
  wire [0:0] v_21591;
  wire [0:0] act_21592;
  wire [0:0] v_21593;
  wire [0:0] v_21594;
  wire [0:0] v_21595;
  reg [0:0] v_21596 = 1'h0;
  wire [0:0] v_21597;
  wire [0:0] v_21598;
  wire [0:0] act_21599;
  wire [0:0] v_21600;
  wire [0:0] v_21601;
  wire [0:0] v_21602;
  reg [0:0] v_21603 = 1'h0;
  wire [0:0] v_21604;
  wire [0:0] v_21605;
  wire [0:0] act_21606;
  wire [0:0] v_21607;
  wire [0:0] v_21608;
  wire [0:0] v_21609;
  wire [0:0] vin0_consume_en_21610;
  wire [0:0] vout_canPeek_21610;
  wire [7:0] vout_peek_21610;
  wire [0:0] v_21611;
  wire [0:0] v_21612;
  function [0:0] mux_21612(input [0:0] sel);
    case (sel) 0: mux_21612 = 1'h0; 1: mux_21612 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21613;
  wire [0:0] v_21614;
  wire [0:0] v_21615;
  wire [0:0] v_21616;
  wire [0:0] v_21617;
  function [0:0] mux_21617(input [0:0] sel);
    case (sel) 0: mux_21617 = 1'h0; 1: mux_21617 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21618;
  wire [0:0] vin0_consume_en_21619;
  wire [0:0] vout_canPeek_21619;
  wire [7:0] vout_peek_21619;
  wire [0:0] v_21620;
  wire [0:0] v_21621;
  function [0:0] mux_21621(input [0:0] sel);
    case (sel) 0: mux_21621 = 1'h0; 1: mux_21621 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21622;
  function [0:0] mux_21622(input [0:0] sel);
    case (sel) 0: mux_21622 = 1'h0; 1: mux_21622 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21623;
  wire [0:0] v_21624;
  wire [0:0] v_21625;
  wire [0:0] v_21626;
  wire [0:0] v_21627;
  wire [0:0] v_21628;
  wire [0:0] v_21629;
  function [0:0] mux_21629(input [0:0] sel);
    case (sel) 0: mux_21629 = 1'h0; 1: mux_21629 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21630;
  wire [0:0] v_21631;
  wire [0:0] v_21632;
  wire [0:0] v_21633;
  wire [0:0] v_21634;
  function [0:0] mux_21634(input [0:0] sel);
    case (sel) 0: mux_21634 = 1'h0; 1: mux_21634 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21635;
  wire [0:0] v_21636;
  wire [0:0] v_21637;
  wire [0:0] v_21638;
  function [0:0] mux_21638(input [0:0] sel);
    case (sel) 0: mux_21638 = 1'h0; 1: mux_21638 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21639;
  function [0:0] mux_21639(input [0:0] sel);
    case (sel) 0: mux_21639 = 1'h0; 1: mux_21639 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_21640 = 1'h0;
  wire [0:0] v_21641;
  wire [0:0] v_21642;
  wire [0:0] act_21643;
  wire [0:0] v_21644;
  wire [0:0] v_21645;
  wire [0:0] v_21646;
  wire [0:0] vin0_consume_en_21647;
  wire [0:0] vout_canPeek_21647;
  wire [7:0] vout_peek_21647;
  wire [0:0] v_21648;
  wire [0:0] v_21649;
  function [0:0] mux_21649(input [0:0] sel);
    case (sel) 0: mux_21649 = 1'h0; 1: mux_21649 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21650;
  wire [0:0] v_21651;
  wire [0:0] v_21652;
  wire [0:0] v_21653;
  wire [0:0] v_21654;
  function [0:0] mux_21654(input [0:0] sel);
    case (sel) 0: mux_21654 = 1'h0; 1: mux_21654 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21655;
  wire [0:0] vin0_consume_en_21656;
  wire [0:0] vout_canPeek_21656;
  wire [7:0] vout_peek_21656;
  wire [0:0] v_21657;
  wire [0:0] v_21658;
  function [0:0] mux_21658(input [0:0] sel);
    case (sel) 0: mux_21658 = 1'h0; 1: mux_21658 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21659;
  function [0:0] mux_21659(input [0:0] sel);
    case (sel) 0: mux_21659 = 1'h0; 1: mux_21659 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21660;
  wire [0:0] v_21661;
  wire [0:0] v_21662;
  wire [0:0] v_21663;
  wire [0:0] v_21664;
  wire [0:0] v_21665;
  wire [0:0] v_21666;
  function [0:0] mux_21666(input [0:0] sel);
    case (sel) 0: mux_21666 = 1'h0; 1: mux_21666 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21667;
  function [0:0] mux_21667(input [0:0] sel);
    case (sel) 0: mux_21667 = 1'h0; 1: mux_21667 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21668;
  wire [0:0] v_21669;
  wire [0:0] v_21670;
  wire [0:0] v_21671;
  function [0:0] mux_21671(input [0:0] sel);
    case (sel) 0: mux_21671 = 1'h0; 1: mux_21671 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21672;
  function [0:0] mux_21672(input [0:0] sel);
    case (sel) 0: mux_21672 = 1'h0; 1: mux_21672 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21673;
  wire [0:0] v_21674;
  wire [0:0] v_21675;
  wire [0:0] v_21676;
  wire [0:0] v_21677;
  wire [0:0] v_21678;
  function [0:0] mux_21678(input [0:0] sel);
    case (sel) 0: mux_21678 = 1'h0; 1: mux_21678 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21679;
  wire [0:0] v_21680;
  wire [0:0] v_21681;
  wire [0:0] v_21682;
  wire [0:0] v_21683;
  function [0:0] mux_21683(input [0:0] sel);
    case (sel) 0: mux_21683 = 1'h0; 1: mux_21683 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21684;
  wire [0:0] v_21685;
  wire [0:0] v_21686;
  wire [0:0] v_21687;
  function [0:0] mux_21687(input [0:0] sel);
    case (sel) 0: mux_21687 = 1'h0; 1: mux_21687 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21688;
  function [0:0] mux_21688(input [0:0] sel);
    case (sel) 0: mux_21688 = 1'h0; 1: mux_21688 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_21689 = 1'h0;
  wire [0:0] v_21690;
  wire [0:0] v_21691;
  wire [0:0] act_21692;
  wire [0:0] v_21693;
  wire [0:0] v_21694;
  wire [0:0] v_21695;
  reg [0:0] v_21696 = 1'h0;
  wire [0:0] v_21697;
  wire [0:0] v_21698;
  wire [0:0] act_21699;
  wire [0:0] v_21700;
  wire [0:0] v_21701;
  wire [0:0] v_21702;
  wire [0:0] vin0_consume_en_21703;
  wire [0:0] vout_canPeek_21703;
  wire [7:0] vout_peek_21703;
  wire [0:0] v_21704;
  wire [0:0] v_21705;
  function [0:0] mux_21705(input [0:0] sel);
    case (sel) 0: mux_21705 = 1'h0; 1: mux_21705 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21706;
  wire [0:0] v_21707;
  wire [0:0] v_21708;
  wire [0:0] v_21709;
  wire [0:0] v_21710;
  function [0:0] mux_21710(input [0:0] sel);
    case (sel) 0: mux_21710 = 1'h0; 1: mux_21710 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21711;
  wire [0:0] vin0_consume_en_21712;
  wire [0:0] vout_canPeek_21712;
  wire [7:0] vout_peek_21712;
  wire [0:0] v_21713;
  wire [0:0] v_21714;
  function [0:0] mux_21714(input [0:0] sel);
    case (sel) 0: mux_21714 = 1'h0; 1: mux_21714 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21715;
  function [0:0] mux_21715(input [0:0] sel);
    case (sel) 0: mux_21715 = 1'h0; 1: mux_21715 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21716;
  wire [0:0] v_21717;
  wire [0:0] v_21718;
  wire [0:0] v_21719;
  wire [0:0] v_21720;
  wire [0:0] v_21721;
  wire [0:0] v_21722;
  function [0:0] mux_21722(input [0:0] sel);
    case (sel) 0: mux_21722 = 1'h0; 1: mux_21722 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21723;
  wire [0:0] v_21724;
  wire [0:0] v_21725;
  wire [0:0] v_21726;
  wire [0:0] v_21727;
  function [0:0] mux_21727(input [0:0] sel);
    case (sel) 0: mux_21727 = 1'h0; 1: mux_21727 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21728;
  wire [0:0] v_21729;
  wire [0:0] v_21730;
  wire [0:0] v_21731;
  function [0:0] mux_21731(input [0:0] sel);
    case (sel) 0: mux_21731 = 1'h0; 1: mux_21731 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21732;
  function [0:0] mux_21732(input [0:0] sel);
    case (sel) 0: mux_21732 = 1'h0; 1: mux_21732 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_21733 = 1'h0;
  wire [0:0] v_21734;
  wire [0:0] v_21735;
  wire [0:0] act_21736;
  wire [0:0] v_21737;
  wire [0:0] v_21738;
  wire [0:0] v_21739;
  wire [0:0] vin0_consume_en_21740;
  wire [0:0] vout_canPeek_21740;
  wire [7:0] vout_peek_21740;
  wire [0:0] v_21741;
  wire [0:0] v_21742;
  function [0:0] mux_21742(input [0:0] sel);
    case (sel) 0: mux_21742 = 1'h0; 1: mux_21742 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21743;
  wire [0:0] v_21744;
  wire [0:0] v_21745;
  wire [0:0] v_21746;
  wire [0:0] v_21747;
  function [0:0] mux_21747(input [0:0] sel);
    case (sel) 0: mux_21747 = 1'h0; 1: mux_21747 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21748;
  wire [0:0] vin0_consume_en_21749;
  wire [0:0] vout_canPeek_21749;
  wire [7:0] vout_peek_21749;
  wire [0:0] v_21750;
  wire [0:0] v_21751;
  function [0:0] mux_21751(input [0:0] sel);
    case (sel) 0: mux_21751 = 1'h0; 1: mux_21751 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21752;
  function [0:0] mux_21752(input [0:0] sel);
    case (sel) 0: mux_21752 = 1'h0; 1: mux_21752 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21753;
  wire [0:0] v_21754;
  wire [0:0] v_21755;
  wire [0:0] v_21756;
  wire [0:0] v_21757;
  wire [0:0] v_21758;
  wire [0:0] v_21759;
  function [0:0] mux_21759(input [0:0] sel);
    case (sel) 0: mux_21759 = 1'h0; 1: mux_21759 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21760;
  function [0:0] mux_21760(input [0:0] sel);
    case (sel) 0: mux_21760 = 1'h0; 1: mux_21760 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21761;
  wire [0:0] v_21762;
  wire [0:0] v_21763;
  wire [0:0] v_21764;
  function [0:0] mux_21764(input [0:0] sel);
    case (sel) 0: mux_21764 = 1'h0; 1: mux_21764 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21765;
  function [0:0] mux_21765(input [0:0] sel);
    case (sel) 0: mux_21765 = 1'h0; 1: mux_21765 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21766;
  wire [0:0] v_21767;
  wire [0:0] v_21768;
  wire [0:0] v_21769;
  wire [0:0] v_21770;
  wire [0:0] v_21771;
  function [0:0] mux_21771(input [0:0] sel);
    case (sel) 0: mux_21771 = 1'h0; 1: mux_21771 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21772;
  function [0:0] mux_21772(input [0:0] sel);
    case (sel) 0: mux_21772 = 1'h0; 1: mux_21772 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21773;
  wire [0:0] v_21774;
  wire [0:0] v_21775;
  wire [0:0] v_21776;
  function [0:0] mux_21776(input [0:0] sel);
    case (sel) 0: mux_21776 = 1'h0; 1: mux_21776 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21777;
  function [0:0] mux_21777(input [0:0] sel);
    case (sel) 0: mux_21777 = 1'h0; 1: mux_21777 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21778;
  wire [0:0] v_21779;
  wire [0:0] v_21780;
  wire [0:0] v_21781;
  wire [0:0] v_21782;
  wire [0:0] v_21783;
  function [0:0] mux_21783(input [0:0] sel);
    case (sel) 0: mux_21783 = 1'h0; 1: mux_21783 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21784;
  function [0:0] mux_21784(input [0:0] sel);
    case (sel) 0: mux_21784 = 1'h0; 1: mux_21784 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21785;
  wire [0:0] v_21786;
  wire [0:0] v_21787;
  wire [0:0] v_21788;
  function [0:0] mux_21788(input [0:0] sel);
    case (sel) 0: mux_21788 = 1'h0; 1: mux_21788 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21789;
  function [0:0] mux_21789(input [0:0] sel);
    case (sel) 0: mux_21789 = 1'h0; 1: mux_21789 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21790;
  wire [0:0] v_21791;
  wire [0:0] v_21792;
  wire [0:0] v_21793;
  wire [0:0] v_21794;
  wire [0:0] v_21795;
  function [0:0] mux_21795(input [0:0] sel);
    case (sel) 0: mux_21795 = 1'h0; 1: mux_21795 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21796;
  wire [0:0] v_21797;
  wire [0:0] v_21798;
  wire [0:0] v_21799;
  wire [0:0] v_21800;
  function [0:0] mux_21800(input [0:0] sel);
    case (sel) 0: mux_21800 = 1'h0; 1: mux_21800 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21801;
  wire [0:0] v_21802;
  wire [0:0] v_21803;
  wire [0:0] v_21804;
  function [0:0] mux_21804(input [0:0] sel);
    case (sel) 0: mux_21804 = 1'h0; 1: mux_21804 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21805;
  function [0:0] mux_21805(input [0:0] sel);
    case (sel) 0: mux_21805 = 1'h0; 1: mux_21805 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_21806 = 1'h0;
  wire [0:0] v_21807;
  wire [0:0] v_21808;
  wire [0:0] act_21809;
  wire [0:0] v_21810;
  wire [0:0] v_21811;
  wire [0:0] v_21812;
  reg [0:0] v_21813 = 1'h0;
  wire [0:0] v_21814;
  wire [0:0] v_21815;
  wire [0:0] act_21816;
  wire [0:0] v_21817;
  wire [0:0] v_21818;
  wire [0:0] v_21819;
  reg [0:0] v_21820 = 1'h0;
  wire [0:0] v_21821;
  wire [0:0] v_21822;
  wire [0:0] act_21823;
  wire [0:0] v_21824;
  wire [0:0] v_21825;
  wire [0:0] v_21826;
  reg [0:0] v_21827 = 1'h0;
  wire [0:0] v_21828;
  wire [0:0] v_21829;
  wire [0:0] act_21830;
  wire [0:0] v_21831;
  wire [0:0] v_21832;
  wire [0:0] v_21833;
  wire [0:0] vin0_consume_en_21834;
  wire [0:0] vout_canPeek_21834;
  wire [7:0] vout_peek_21834;
  wire [0:0] v_21835;
  wire [0:0] v_21836;
  function [0:0] mux_21836(input [0:0] sel);
    case (sel) 0: mux_21836 = 1'h0; 1: mux_21836 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21837;
  wire [0:0] v_21838;
  wire [0:0] v_21839;
  wire [0:0] v_21840;
  wire [0:0] v_21841;
  function [0:0] mux_21841(input [0:0] sel);
    case (sel) 0: mux_21841 = 1'h0; 1: mux_21841 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21842;
  wire [0:0] vin0_consume_en_21843;
  wire [0:0] vout_canPeek_21843;
  wire [7:0] vout_peek_21843;
  wire [0:0] v_21844;
  wire [0:0] v_21845;
  function [0:0] mux_21845(input [0:0] sel);
    case (sel) 0: mux_21845 = 1'h0; 1: mux_21845 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21846;
  function [0:0] mux_21846(input [0:0] sel);
    case (sel) 0: mux_21846 = 1'h0; 1: mux_21846 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21847;
  wire [0:0] v_21848;
  wire [0:0] v_21849;
  wire [0:0] v_21850;
  wire [0:0] v_21851;
  wire [0:0] v_21852;
  wire [0:0] v_21853;
  function [0:0] mux_21853(input [0:0] sel);
    case (sel) 0: mux_21853 = 1'h0; 1: mux_21853 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21854;
  wire [0:0] v_21855;
  wire [0:0] v_21856;
  wire [0:0] v_21857;
  wire [0:0] v_21858;
  function [0:0] mux_21858(input [0:0] sel);
    case (sel) 0: mux_21858 = 1'h0; 1: mux_21858 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21859;
  wire [0:0] v_21860;
  wire [0:0] v_21861;
  wire [0:0] v_21862;
  function [0:0] mux_21862(input [0:0] sel);
    case (sel) 0: mux_21862 = 1'h0; 1: mux_21862 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21863;
  function [0:0] mux_21863(input [0:0] sel);
    case (sel) 0: mux_21863 = 1'h0; 1: mux_21863 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_21864 = 1'h0;
  wire [0:0] v_21865;
  wire [0:0] v_21866;
  wire [0:0] act_21867;
  wire [0:0] v_21868;
  wire [0:0] v_21869;
  wire [0:0] v_21870;
  wire [0:0] vin0_consume_en_21871;
  wire [0:0] vout_canPeek_21871;
  wire [7:0] vout_peek_21871;
  wire [0:0] v_21872;
  wire [0:0] v_21873;
  function [0:0] mux_21873(input [0:0] sel);
    case (sel) 0: mux_21873 = 1'h0; 1: mux_21873 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21874;
  wire [0:0] v_21875;
  wire [0:0] v_21876;
  wire [0:0] v_21877;
  wire [0:0] v_21878;
  function [0:0] mux_21878(input [0:0] sel);
    case (sel) 0: mux_21878 = 1'h0; 1: mux_21878 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21879;
  wire [0:0] vin0_consume_en_21880;
  wire [0:0] vout_canPeek_21880;
  wire [7:0] vout_peek_21880;
  wire [0:0] v_21881;
  wire [0:0] v_21882;
  function [0:0] mux_21882(input [0:0] sel);
    case (sel) 0: mux_21882 = 1'h0; 1: mux_21882 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21883;
  function [0:0] mux_21883(input [0:0] sel);
    case (sel) 0: mux_21883 = 1'h0; 1: mux_21883 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21884;
  wire [0:0] v_21885;
  wire [0:0] v_21886;
  wire [0:0] v_21887;
  wire [0:0] v_21888;
  wire [0:0] v_21889;
  wire [0:0] v_21890;
  function [0:0] mux_21890(input [0:0] sel);
    case (sel) 0: mux_21890 = 1'h0; 1: mux_21890 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21891;
  function [0:0] mux_21891(input [0:0] sel);
    case (sel) 0: mux_21891 = 1'h0; 1: mux_21891 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21892;
  wire [0:0] v_21893;
  wire [0:0] v_21894;
  wire [0:0] v_21895;
  function [0:0] mux_21895(input [0:0] sel);
    case (sel) 0: mux_21895 = 1'h0; 1: mux_21895 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21896;
  function [0:0] mux_21896(input [0:0] sel);
    case (sel) 0: mux_21896 = 1'h0; 1: mux_21896 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21897;
  wire [0:0] v_21898;
  wire [0:0] v_21899;
  wire [0:0] v_21900;
  wire [0:0] v_21901;
  wire [0:0] v_21902;
  function [0:0] mux_21902(input [0:0] sel);
    case (sel) 0: mux_21902 = 1'h0; 1: mux_21902 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21903;
  wire [0:0] v_21904;
  wire [0:0] v_21905;
  wire [0:0] v_21906;
  wire [0:0] v_21907;
  function [0:0] mux_21907(input [0:0] sel);
    case (sel) 0: mux_21907 = 1'h0; 1: mux_21907 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21908;
  wire [0:0] v_21909;
  wire [0:0] v_21910;
  wire [0:0] v_21911;
  function [0:0] mux_21911(input [0:0] sel);
    case (sel) 0: mux_21911 = 1'h0; 1: mux_21911 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21912;
  function [0:0] mux_21912(input [0:0] sel);
    case (sel) 0: mux_21912 = 1'h0; 1: mux_21912 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_21913 = 1'h0;
  wire [0:0] v_21914;
  wire [0:0] v_21915;
  wire [0:0] act_21916;
  wire [0:0] v_21917;
  wire [0:0] v_21918;
  wire [0:0] v_21919;
  reg [0:0] v_21920 = 1'h0;
  wire [0:0] v_21921;
  wire [0:0] v_21922;
  wire [0:0] act_21923;
  wire [0:0] v_21924;
  wire [0:0] v_21925;
  wire [0:0] v_21926;
  wire [0:0] vin0_consume_en_21927;
  wire [0:0] vout_canPeek_21927;
  wire [7:0] vout_peek_21927;
  wire [0:0] v_21928;
  wire [0:0] v_21929;
  function [0:0] mux_21929(input [0:0] sel);
    case (sel) 0: mux_21929 = 1'h0; 1: mux_21929 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21930;
  wire [0:0] v_21931;
  wire [0:0] v_21932;
  wire [0:0] v_21933;
  wire [0:0] v_21934;
  function [0:0] mux_21934(input [0:0] sel);
    case (sel) 0: mux_21934 = 1'h0; 1: mux_21934 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21935;
  wire [0:0] vin0_consume_en_21936;
  wire [0:0] vout_canPeek_21936;
  wire [7:0] vout_peek_21936;
  wire [0:0] v_21937;
  wire [0:0] v_21938;
  function [0:0] mux_21938(input [0:0] sel);
    case (sel) 0: mux_21938 = 1'h0; 1: mux_21938 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21939;
  function [0:0] mux_21939(input [0:0] sel);
    case (sel) 0: mux_21939 = 1'h0; 1: mux_21939 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21940;
  wire [0:0] v_21941;
  wire [0:0] v_21942;
  wire [0:0] v_21943;
  wire [0:0] v_21944;
  wire [0:0] v_21945;
  wire [0:0] v_21946;
  function [0:0] mux_21946(input [0:0] sel);
    case (sel) 0: mux_21946 = 1'h0; 1: mux_21946 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21947;
  wire [0:0] v_21948;
  wire [0:0] v_21949;
  wire [0:0] v_21950;
  wire [0:0] v_21951;
  function [0:0] mux_21951(input [0:0] sel);
    case (sel) 0: mux_21951 = 1'h0; 1: mux_21951 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21952;
  wire [0:0] v_21953;
  wire [0:0] v_21954;
  wire [0:0] v_21955;
  function [0:0] mux_21955(input [0:0] sel);
    case (sel) 0: mux_21955 = 1'h0; 1: mux_21955 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21956;
  function [0:0] mux_21956(input [0:0] sel);
    case (sel) 0: mux_21956 = 1'h0; 1: mux_21956 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_21957 = 1'h0;
  wire [0:0] v_21958;
  wire [0:0] v_21959;
  wire [0:0] act_21960;
  wire [0:0] v_21961;
  wire [0:0] v_21962;
  wire [0:0] v_21963;
  wire [0:0] vin0_consume_en_21964;
  wire [0:0] vout_canPeek_21964;
  wire [7:0] vout_peek_21964;
  wire [0:0] v_21965;
  wire [0:0] v_21966;
  function [0:0] mux_21966(input [0:0] sel);
    case (sel) 0: mux_21966 = 1'h0; 1: mux_21966 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21967;
  wire [0:0] v_21968;
  wire [0:0] v_21969;
  wire [0:0] v_21970;
  wire [0:0] v_21971;
  function [0:0] mux_21971(input [0:0] sel);
    case (sel) 0: mux_21971 = 1'h0; 1: mux_21971 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21972;
  wire [0:0] vin0_consume_en_21973;
  wire [0:0] vout_canPeek_21973;
  wire [7:0] vout_peek_21973;
  wire [0:0] v_21974;
  wire [0:0] v_21975;
  function [0:0] mux_21975(input [0:0] sel);
    case (sel) 0: mux_21975 = 1'h0; 1: mux_21975 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21976;
  function [0:0] mux_21976(input [0:0] sel);
    case (sel) 0: mux_21976 = 1'h0; 1: mux_21976 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21977;
  wire [0:0] v_21978;
  wire [0:0] v_21979;
  wire [0:0] v_21980;
  wire [0:0] v_21981;
  wire [0:0] v_21982;
  wire [0:0] v_21983;
  function [0:0] mux_21983(input [0:0] sel);
    case (sel) 0: mux_21983 = 1'h0; 1: mux_21983 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21984;
  function [0:0] mux_21984(input [0:0] sel);
    case (sel) 0: mux_21984 = 1'h0; 1: mux_21984 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21985;
  wire [0:0] v_21986;
  wire [0:0] v_21987;
  wire [0:0] v_21988;
  function [0:0] mux_21988(input [0:0] sel);
    case (sel) 0: mux_21988 = 1'h0; 1: mux_21988 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21989;
  function [0:0] mux_21989(input [0:0] sel);
    case (sel) 0: mux_21989 = 1'h0; 1: mux_21989 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21990;
  wire [0:0] v_21991;
  wire [0:0] v_21992;
  wire [0:0] v_21993;
  wire [0:0] v_21994;
  wire [0:0] v_21995;
  function [0:0] mux_21995(input [0:0] sel);
    case (sel) 0: mux_21995 = 1'h0; 1: mux_21995 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_21996;
  function [0:0] mux_21996(input [0:0] sel);
    case (sel) 0: mux_21996 = 1'h0; 1: mux_21996 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_21997;
  wire [0:0] v_21998;
  wire [0:0] v_21999;
  wire [0:0] v_22000;
  function [0:0] mux_22000(input [0:0] sel);
    case (sel) 0: mux_22000 = 1'h0; 1: mux_22000 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22001;
  function [0:0] mux_22001(input [0:0] sel);
    case (sel) 0: mux_22001 = 1'h0; 1: mux_22001 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22002;
  wire [0:0] v_22003;
  wire [0:0] v_22004;
  wire [0:0] v_22005;
  wire [0:0] v_22006;
  wire [0:0] v_22007;
  function [0:0] mux_22007(input [0:0] sel);
    case (sel) 0: mux_22007 = 1'h0; 1: mux_22007 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22008;
  wire [0:0] v_22009;
  wire [0:0] v_22010;
  wire [0:0] v_22011;
  wire [0:0] v_22012;
  function [0:0] mux_22012(input [0:0] sel);
    case (sel) 0: mux_22012 = 1'h0; 1: mux_22012 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22013;
  wire [0:0] v_22014;
  wire [0:0] v_22015;
  wire [0:0] v_22016;
  function [0:0] mux_22016(input [0:0] sel);
    case (sel) 0: mux_22016 = 1'h0; 1: mux_22016 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22017;
  function [0:0] mux_22017(input [0:0] sel);
    case (sel) 0: mux_22017 = 1'h0; 1: mux_22017 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_22018 = 1'h0;
  wire [0:0] v_22019;
  wire [0:0] v_22020;
  wire [0:0] act_22021;
  wire [0:0] v_22022;
  wire [0:0] v_22023;
  wire [0:0] v_22024;
  reg [0:0] v_22025 = 1'h0;
  wire [0:0] v_22026;
  wire [0:0] v_22027;
  wire [0:0] act_22028;
  wire [0:0] v_22029;
  wire [0:0] v_22030;
  wire [0:0] v_22031;
  reg [0:0] v_22032 = 1'h0;
  wire [0:0] v_22033;
  wire [0:0] v_22034;
  wire [0:0] act_22035;
  wire [0:0] v_22036;
  wire [0:0] v_22037;
  wire [0:0] v_22038;
  wire [0:0] vin0_consume_en_22039;
  wire [0:0] vout_canPeek_22039;
  wire [7:0] vout_peek_22039;
  wire [0:0] v_22040;
  wire [0:0] v_22041;
  function [0:0] mux_22041(input [0:0] sel);
    case (sel) 0: mux_22041 = 1'h0; 1: mux_22041 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22042;
  wire [0:0] v_22043;
  wire [0:0] v_22044;
  wire [0:0] v_22045;
  wire [0:0] v_22046;
  function [0:0] mux_22046(input [0:0] sel);
    case (sel) 0: mux_22046 = 1'h0; 1: mux_22046 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22047;
  wire [0:0] vin0_consume_en_22048;
  wire [0:0] vout_canPeek_22048;
  wire [7:0] vout_peek_22048;
  wire [0:0] v_22049;
  wire [0:0] v_22050;
  function [0:0] mux_22050(input [0:0] sel);
    case (sel) 0: mux_22050 = 1'h0; 1: mux_22050 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22051;
  function [0:0] mux_22051(input [0:0] sel);
    case (sel) 0: mux_22051 = 1'h0; 1: mux_22051 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22052;
  wire [0:0] v_22053;
  wire [0:0] v_22054;
  wire [0:0] v_22055;
  wire [0:0] v_22056;
  wire [0:0] v_22057;
  wire [0:0] v_22058;
  function [0:0] mux_22058(input [0:0] sel);
    case (sel) 0: mux_22058 = 1'h0; 1: mux_22058 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22059;
  wire [0:0] v_22060;
  wire [0:0] v_22061;
  wire [0:0] v_22062;
  wire [0:0] v_22063;
  function [0:0] mux_22063(input [0:0] sel);
    case (sel) 0: mux_22063 = 1'h0; 1: mux_22063 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22064;
  wire [0:0] v_22065;
  wire [0:0] v_22066;
  wire [0:0] v_22067;
  function [0:0] mux_22067(input [0:0] sel);
    case (sel) 0: mux_22067 = 1'h0; 1: mux_22067 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22068;
  function [0:0] mux_22068(input [0:0] sel);
    case (sel) 0: mux_22068 = 1'h0; 1: mux_22068 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_22069 = 1'h0;
  wire [0:0] v_22070;
  wire [0:0] v_22071;
  wire [0:0] act_22072;
  wire [0:0] v_22073;
  wire [0:0] v_22074;
  wire [0:0] v_22075;
  wire [0:0] vin0_consume_en_22076;
  wire [0:0] vout_canPeek_22076;
  wire [7:0] vout_peek_22076;
  wire [0:0] v_22077;
  wire [0:0] v_22078;
  function [0:0] mux_22078(input [0:0] sel);
    case (sel) 0: mux_22078 = 1'h0; 1: mux_22078 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22079;
  wire [0:0] v_22080;
  wire [0:0] v_22081;
  wire [0:0] v_22082;
  wire [0:0] v_22083;
  function [0:0] mux_22083(input [0:0] sel);
    case (sel) 0: mux_22083 = 1'h0; 1: mux_22083 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22084;
  wire [0:0] vin0_consume_en_22085;
  wire [0:0] vout_canPeek_22085;
  wire [7:0] vout_peek_22085;
  wire [0:0] v_22086;
  wire [0:0] v_22087;
  function [0:0] mux_22087(input [0:0] sel);
    case (sel) 0: mux_22087 = 1'h0; 1: mux_22087 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22088;
  function [0:0] mux_22088(input [0:0] sel);
    case (sel) 0: mux_22088 = 1'h0; 1: mux_22088 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22089;
  wire [0:0] v_22090;
  wire [0:0] v_22091;
  wire [0:0] v_22092;
  wire [0:0] v_22093;
  wire [0:0] v_22094;
  wire [0:0] v_22095;
  function [0:0] mux_22095(input [0:0] sel);
    case (sel) 0: mux_22095 = 1'h0; 1: mux_22095 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22096;
  function [0:0] mux_22096(input [0:0] sel);
    case (sel) 0: mux_22096 = 1'h0; 1: mux_22096 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22097;
  wire [0:0] v_22098;
  wire [0:0] v_22099;
  wire [0:0] v_22100;
  function [0:0] mux_22100(input [0:0] sel);
    case (sel) 0: mux_22100 = 1'h0; 1: mux_22100 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22101;
  function [0:0] mux_22101(input [0:0] sel);
    case (sel) 0: mux_22101 = 1'h0; 1: mux_22101 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22102;
  wire [0:0] v_22103;
  wire [0:0] v_22104;
  wire [0:0] v_22105;
  wire [0:0] v_22106;
  wire [0:0] v_22107;
  function [0:0] mux_22107(input [0:0] sel);
    case (sel) 0: mux_22107 = 1'h0; 1: mux_22107 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22108;
  wire [0:0] v_22109;
  wire [0:0] v_22110;
  wire [0:0] v_22111;
  wire [0:0] v_22112;
  function [0:0] mux_22112(input [0:0] sel);
    case (sel) 0: mux_22112 = 1'h0; 1: mux_22112 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22113;
  wire [0:0] v_22114;
  wire [0:0] v_22115;
  wire [0:0] v_22116;
  function [0:0] mux_22116(input [0:0] sel);
    case (sel) 0: mux_22116 = 1'h0; 1: mux_22116 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22117;
  function [0:0] mux_22117(input [0:0] sel);
    case (sel) 0: mux_22117 = 1'h0; 1: mux_22117 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_22118 = 1'h0;
  wire [0:0] v_22119;
  wire [0:0] v_22120;
  wire [0:0] act_22121;
  wire [0:0] v_22122;
  wire [0:0] v_22123;
  wire [0:0] v_22124;
  reg [0:0] v_22125 = 1'h0;
  wire [0:0] v_22126;
  wire [0:0] v_22127;
  wire [0:0] act_22128;
  wire [0:0] v_22129;
  wire [0:0] v_22130;
  wire [0:0] v_22131;
  wire [0:0] vin0_consume_en_22132;
  wire [0:0] vout_canPeek_22132;
  wire [7:0] vout_peek_22132;
  wire [0:0] v_22133;
  wire [0:0] v_22134;
  function [0:0] mux_22134(input [0:0] sel);
    case (sel) 0: mux_22134 = 1'h0; 1: mux_22134 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22135;
  wire [0:0] v_22136;
  wire [0:0] v_22137;
  wire [0:0] v_22138;
  wire [0:0] v_22139;
  function [0:0] mux_22139(input [0:0] sel);
    case (sel) 0: mux_22139 = 1'h0; 1: mux_22139 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22140;
  wire [0:0] vin0_consume_en_22141;
  wire [0:0] vout_canPeek_22141;
  wire [7:0] vout_peek_22141;
  wire [0:0] v_22142;
  wire [0:0] v_22143;
  function [0:0] mux_22143(input [0:0] sel);
    case (sel) 0: mux_22143 = 1'h0; 1: mux_22143 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22144;
  function [0:0] mux_22144(input [0:0] sel);
    case (sel) 0: mux_22144 = 1'h0; 1: mux_22144 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22145;
  wire [0:0] v_22146;
  wire [0:0] v_22147;
  wire [0:0] v_22148;
  wire [0:0] v_22149;
  wire [0:0] v_22150;
  wire [0:0] v_22151;
  function [0:0] mux_22151(input [0:0] sel);
    case (sel) 0: mux_22151 = 1'h0; 1: mux_22151 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22152;
  wire [0:0] v_22153;
  wire [0:0] v_22154;
  wire [0:0] v_22155;
  wire [0:0] v_22156;
  function [0:0] mux_22156(input [0:0] sel);
    case (sel) 0: mux_22156 = 1'h0; 1: mux_22156 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22157;
  wire [0:0] v_22158;
  wire [0:0] v_22159;
  wire [0:0] v_22160;
  function [0:0] mux_22160(input [0:0] sel);
    case (sel) 0: mux_22160 = 1'h0; 1: mux_22160 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22161;
  function [0:0] mux_22161(input [0:0] sel);
    case (sel) 0: mux_22161 = 1'h0; 1: mux_22161 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_22162 = 1'h0;
  wire [0:0] v_22163;
  wire [0:0] v_22164;
  wire [0:0] act_22165;
  wire [0:0] v_22166;
  wire [0:0] v_22167;
  wire [0:0] v_22168;
  wire [0:0] vin0_consume_en_22169;
  wire [0:0] vout_canPeek_22169;
  wire [7:0] vout_peek_22169;
  wire [0:0] v_22170;
  wire [0:0] v_22171;
  function [0:0] mux_22171(input [0:0] sel);
    case (sel) 0: mux_22171 = 1'h0; 1: mux_22171 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22172;
  wire [0:0] v_22173;
  wire [0:0] v_22174;
  wire [0:0] v_22175;
  wire [0:0] v_22176;
  function [0:0] mux_22176(input [0:0] sel);
    case (sel) 0: mux_22176 = 1'h0; 1: mux_22176 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22177;
  wire [0:0] vin0_consume_en_22178;
  wire [0:0] vout_canPeek_22178;
  wire [7:0] vout_peek_22178;
  wire [0:0] v_22179;
  wire [0:0] v_22180;
  function [0:0] mux_22180(input [0:0] sel);
    case (sel) 0: mux_22180 = 1'h0; 1: mux_22180 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22181;
  function [0:0] mux_22181(input [0:0] sel);
    case (sel) 0: mux_22181 = 1'h0; 1: mux_22181 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22182;
  wire [0:0] v_22183;
  wire [0:0] v_22184;
  wire [0:0] v_22185;
  wire [0:0] v_22186;
  wire [0:0] v_22187;
  wire [0:0] v_22188;
  function [0:0] mux_22188(input [0:0] sel);
    case (sel) 0: mux_22188 = 1'h0; 1: mux_22188 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22189;
  function [0:0] mux_22189(input [0:0] sel);
    case (sel) 0: mux_22189 = 1'h0; 1: mux_22189 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22190;
  wire [0:0] v_22191;
  wire [0:0] v_22192;
  wire [0:0] v_22193;
  function [0:0] mux_22193(input [0:0] sel);
    case (sel) 0: mux_22193 = 1'h0; 1: mux_22193 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22194;
  function [0:0] mux_22194(input [0:0] sel);
    case (sel) 0: mux_22194 = 1'h0; 1: mux_22194 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22195;
  wire [0:0] v_22196;
  wire [0:0] v_22197;
  wire [0:0] v_22198;
  wire [0:0] v_22199;
  wire [0:0] v_22200;
  function [0:0] mux_22200(input [0:0] sel);
    case (sel) 0: mux_22200 = 1'h0; 1: mux_22200 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22201;
  function [0:0] mux_22201(input [0:0] sel);
    case (sel) 0: mux_22201 = 1'h0; 1: mux_22201 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22202;
  wire [0:0] v_22203;
  wire [0:0] v_22204;
  wire [0:0] v_22205;
  function [0:0] mux_22205(input [0:0] sel);
    case (sel) 0: mux_22205 = 1'h0; 1: mux_22205 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22206;
  function [0:0] mux_22206(input [0:0] sel);
    case (sel) 0: mux_22206 = 1'h0; 1: mux_22206 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22207;
  wire [0:0] v_22208;
  wire [0:0] v_22209;
  wire [0:0] v_22210;
  wire [0:0] v_22211;
  wire [0:0] v_22212;
  function [0:0] mux_22212(input [0:0] sel);
    case (sel) 0: mux_22212 = 1'h0; 1: mux_22212 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22213;
  function [0:0] mux_22213(input [0:0] sel);
    case (sel) 0: mux_22213 = 1'h0; 1: mux_22213 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22214;
  wire [0:0] v_22215;
  wire [0:0] v_22216;
  wire [0:0] v_22217;
  function [0:0] mux_22217(input [0:0] sel);
    case (sel) 0: mux_22217 = 1'h0; 1: mux_22217 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22218;
  function [0:0] mux_22218(input [0:0] sel);
    case (sel) 0: mux_22218 = 1'h0; 1: mux_22218 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22219;
  wire [0:0] v_22220;
  wire [0:0] v_22221;
  wire [0:0] v_22222;
  wire [0:0] v_22223;
  wire [0:0] v_22224;
  function [0:0] mux_22224(input [0:0] sel);
    case (sel) 0: mux_22224 = 1'h0; 1: mux_22224 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22225;
  function [0:0] mux_22225(input [0:0] sel);
    case (sel) 0: mux_22225 = 1'h0; 1: mux_22225 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22226;
  wire [0:0] v_22227;
  wire [0:0] v_22228;
  wire [0:0] v_22229;
  function [0:0] mux_22229(input [0:0] sel);
    case (sel) 0: mux_22229 = 1'h0; 1: mux_22229 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22230;
  function [0:0] mux_22230(input [0:0] sel);
    case (sel) 0: mux_22230 = 1'h0; 1: mux_22230 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22231;
  wire [0:0] v_22232;
  wire [0:0] v_22233;
  wire [0:0] v_22234;
  wire [0:0] v_22235;
  wire [0:0] v_22236;
  function [0:0] mux_22236(input [0:0] sel);
    case (sel) 0: mux_22236 = 1'h0; 1: mux_22236 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22237;
  function [0:0] mux_22237(input [0:0] sel);
    case (sel) 0: mux_22237 = 1'h0; 1: mux_22237 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22238;
  wire [0:0] v_22239;
  wire [0:0] v_22240;
  wire [0:0] v_22241;
  function [0:0] mux_22241(input [0:0] sel);
    case (sel) 0: mux_22241 = 1'h0; 1: mux_22241 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22242;
  function [0:0] mux_22242(input [0:0] sel);
    case (sel) 0: mux_22242 = 1'h0; 1: mux_22242 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22243;
  wire [0:0] v_22244;
  wire [0:0] v_22245;
  wire [0:0] v_22246;
  wire [0:0] v_22247;
  wire [0:0] v_22248;
  function [0:0] mux_22248(input [0:0] sel);
    case (sel) 0: mux_22248 = 1'h0; 1: mux_22248 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22249;
  function [0:0] mux_22249(input [0:0] sel);
    case (sel) 0: mux_22249 = 1'h0; 1: mux_22249 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22250;
  wire [0:0] v_22251;
  wire [0:0] v_22252;
  wire [0:0] v_22253;
  function [0:0] mux_22253(input [0:0] sel);
    case (sel) 0: mux_22253 = 1'h0; 1: mux_22253 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22254;
  function [0:0] mux_22254(input [0:0] sel);
    case (sel) 0: mux_22254 = 1'h0; 1: mux_22254 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22255;
  wire [0:0] v_22256;
  wire [0:0] v_22257;
  wire [0:0] v_22258;
  wire [0:0] v_22259;
  wire [0:0] v_22260;
  function [0:0] mux_22260(input [0:0] sel);
    case (sel) 0: mux_22260 = 1'h0; 1: mux_22260 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22261;
  function [0:0] mux_22261(input [0:0] sel);
    case (sel) 0: mux_22261 = 1'h0; 1: mux_22261 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22262;
  wire [0:0] v_22263;
  wire [0:0] v_22264;
  wire [0:0] v_22265;
  function [0:0] mux_22265(input [0:0] sel);
    case (sel) 0: mux_22265 = 1'h0; 1: mux_22265 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22266;
  function [0:0] mux_22266(input [0:0] sel);
    case (sel) 0: mux_22266 = 1'h0; 1: mux_22266 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22267;
  wire [0:0] v_22268;
  wire [0:0] v_22269;
  wire [0:0] v_22270;
  wire [0:0] v_22271;
  wire [0:0] v_22272;
  function [0:0] mux_22272(input [0:0] sel);
    case (sel) 0: mux_22272 = 1'h0; 1: mux_22272 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22273;
  function [0:0] mux_22273(input [0:0] sel);
    case (sel) 0: mux_22273 = 1'h0; 1: mux_22273 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22274;
  wire [0:0] v_22275;
  wire [0:0] v_22276;
  wire [0:0] v_22277;
  function [0:0] mux_22277(input [0:0] sel);
    case (sel) 0: mux_22277 = 1'h0; 1: mux_22277 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22278;
  function [0:0] mux_22278(input [0:0] sel);
    case (sel) 0: mux_22278 = 1'h0; 1: mux_22278 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22279;
  wire [0:0] v_22280;
  wire [0:0] v_22281;
  wire [0:0] v_22282;
  wire [0:0] v_22283;
  wire [0:0] v_22284;
  function [0:0] mux_22284(input [0:0] sel);
    case (sel) 0: mux_22284 = 1'h0; 1: mux_22284 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22285;
  function [0:0] mux_22285(input [0:0] sel);
    case (sel) 0: mux_22285 = 1'h0; 1: mux_22285 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22286;
  wire [0:0] v_22287;
  wire [0:0] v_22288;
  wire [0:0] v_22289;
  function [0:0] mux_22289(input [0:0] sel);
    case (sel) 0: mux_22289 = 1'h0; 1: mux_22289 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22290;
  function [0:0] mux_22290(input [0:0] sel);
    case (sel) 0: mux_22290 = 1'h0; 1: mux_22290 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22291;
  wire [0:0] v_22292;
  wire [0:0] v_22293;
  wire [0:0] v_22294;
  wire [0:0] v_22295;
  wire [0:0] v_22296;
  function [0:0] mux_22296(input [0:0] sel);
    case (sel) 0: mux_22296 = 1'h0; 1: mux_22296 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22297;
  wire [0:0] v_22298;
  wire [0:0] v_22299;
  function [0:0] mux_22299(input [0:0] sel);
    case (sel) 0: mux_22299 = 1'h0; 1: mux_22299 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22300;
  wire [0:0] v_22301;
  wire [0:0] v_22302;
  wire [0:0] v_22303;
  function [0:0] mux_22303(input [0:0] sel);
    case (sel) 0: mux_22303 = 1'h0; 1: mux_22303 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22304;
  function [0:0] mux_22304(input [0:0] sel);
    case (sel) 0: mux_22304 = 1'h0; 1: mux_22304 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22305;
  function [0:0] mux_22305(input [0:0] sel);
    case (sel) 0: mux_22305 = 1'h0; 1: mux_22305 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22306;
  wire [0:0] v_22307;
  wire [0:0] v_22308;
  wire [0:0] v_22309;
  function [0:0] mux_22309(input [0:0] sel);
    case (sel) 0: mux_22309 = 1'h0; 1: mux_22309 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22310;
  function [0:0] mux_22310(input [0:0] sel);
    case (sel) 0: mux_22310 = 1'h0; 1: mux_22310 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22311;
  function [0:0] mux_22311(input [0:0] sel);
    case (sel) 0: mux_22311 = 1'h0; 1: mux_22311 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22312;
  wire [0:0] v_22313;
  wire [0:0] v_22314;
  wire [0:0] v_22315;
  function [0:0] mux_22315(input [0:0] sel);
    case (sel) 0: mux_22315 = 1'h0; 1: mux_22315 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22316;
  function [0:0] mux_22316(input [0:0] sel);
    case (sel) 0: mux_22316 = 1'h0; 1: mux_22316 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22317;
  function [0:0] mux_22317(input [0:0] sel);
    case (sel) 0: mux_22317 = 1'h0; 1: mux_22317 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22318;
  wire [0:0] v_22319;
  wire [0:0] v_22320;
  wire [0:0] v_22321;
  function [0:0] mux_22321(input [0:0] sel);
    case (sel) 0: mux_22321 = 1'h0; 1: mux_22321 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22322;
  function [0:0] mux_22322(input [0:0] sel);
    case (sel) 0: mux_22322 = 1'h0; 1: mux_22322 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22323;
  function [0:0] mux_22323(input [0:0] sel);
    case (sel) 0: mux_22323 = 1'h0; 1: mux_22323 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22324;
  wire [0:0] v_22325;
  wire [0:0] v_22326;
  wire [0:0] v_22327;
  function [0:0] mux_22327(input [0:0] sel);
    case (sel) 0: mux_22327 = 1'h0; 1: mux_22327 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22328;
  function [0:0] mux_22328(input [0:0] sel);
    case (sel) 0: mux_22328 = 1'h0; 1: mux_22328 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22329;
  function [0:0] mux_22329(input [0:0] sel);
    case (sel) 0: mux_22329 = 1'h0; 1: mux_22329 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22330;
  wire [0:0] v_22331;
  wire [0:0] v_22332;
  wire [0:0] v_22333;
  function [0:0] mux_22333(input [0:0] sel);
    case (sel) 0: mux_22333 = 1'h0; 1: mux_22333 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22334;
  function [0:0] mux_22334(input [0:0] sel);
    case (sel) 0: mux_22334 = 1'h0; 1: mux_22334 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22335;
  function [0:0] mux_22335(input [0:0] sel);
    case (sel) 0: mux_22335 = 1'h0; 1: mux_22335 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22336;
  wire [0:0] v_22337;
  wire [0:0] v_22338;
  wire [0:0] v_22339;
  function [0:0] mux_22339(input [0:0] sel);
    case (sel) 0: mux_22339 = 1'h0; 1: mux_22339 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22340;
  function [0:0] mux_22340(input [0:0] sel);
    case (sel) 0: mux_22340 = 1'h0; 1: mux_22340 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22341;
  function [0:0] mux_22341(input [0:0] sel);
    case (sel) 0: mux_22341 = 1'h0; 1: mux_22341 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22342;
  wire [0:0] v_22343;
  wire [0:0] v_22344;
  wire [0:0] v_22345;
  function [0:0] mux_22345(input [0:0] sel);
    case (sel) 0: mux_22345 = 1'h0; 1: mux_22345 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22346;
  function [0:0] mux_22346(input [0:0] sel);
    case (sel) 0: mux_22346 = 1'h0; 1: mux_22346 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22347;
  function [0:0] mux_22347(input [0:0] sel);
    case (sel) 0: mux_22347 = 1'h0; 1: mux_22347 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22348;
  wire [0:0] v_22349;
  wire [0:0] v_22350;
  wire [0:0] v_22351;
  function [0:0] mux_22351(input [0:0] sel);
    case (sel) 0: mux_22351 = 1'h0; 1: mux_22351 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22352;
  function [0:0] mux_22352(input [0:0] sel);
    case (sel) 0: mux_22352 = 1'h0; 1: mux_22352 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22353;
  function [0:0] mux_22353(input [0:0] sel);
    case (sel) 0: mux_22353 = 1'h0; 1: mux_22353 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22354;
  wire [0:0] v_22355;
  wire [0:0] v_22356;
  wire [0:0] v_22357;
  function [0:0] mux_22357(input [0:0] sel);
    case (sel) 0: mux_22357 = 1'h0; 1: mux_22357 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22358;
  function [0:0] mux_22358(input [0:0] sel);
    case (sel) 0: mux_22358 = 1'h0; 1: mux_22358 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22359;
  function [0:0] mux_22359(input [0:0] sel);
    case (sel) 0: mux_22359 = 1'h0; 1: mux_22359 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22360;
  wire [0:0] v_22361;
  wire [0:0] v_22362;
  wire [0:0] v_22363;
  function [0:0] mux_22363(input [0:0] sel);
    case (sel) 0: mux_22363 = 1'h0; 1: mux_22363 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22364;
  function [0:0] mux_22364(input [0:0] sel);
    case (sel) 0: mux_22364 = 1'h0; 1: mux_22364 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22365;
  function [0:0] mux_22365(input [0:0] sel);
    case (sel) 0: mux_22365 = 1'h0; 1: mux_22365 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22366;
  wire [0:0] v_22367;
  wire [0:0] v_22368;
  wire [0:0] v_22369;
  function [0:0] mux_22369(input [0:0] sel);
    case (sel) 0: mux_22369 = 1'h0; 1: mux_22369 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22370;
  function [0:0] mux_22370(input [0:0] sel);
    case (sel) 0: mux_22370 = 1'h0; 1: mux_22370 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22371;
  function [0:0] mux_22371(input [0:0] sel);
    case (sel) 0: mux_22371 = 1'h0; 1: mux_22371 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22372;
  wire [0:0] v_22373;
  wire [0:0] v_22374;
  wire [0:0] v_22375;
  function [0:0] mux_22375(input [0:0] sel);
    case (sel) 0: mux_22375 = 1'h0; 1: mux_22375 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22376;
  function [0:0] mux_22376(input [0:0] sel);
    case (sel) 0: mux_22376 = 1'h0; 1: mux_22376 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22377;
  function [0:0] mux_22377(input [0:0] sel);
    case (sel) 0: mux_22377 = 1'h0; 1: mux_22377 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22378;
  wire [0:0] v_22380;
  function [0:0] mux_22380(input [0:0] sel);
    case (sel) 0: mux_22380 = 1'h0; 1: mux_22380 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_22381;
  reg [7:0] v_22384 = 8'h0;
  wire [7:0] v_22385;
  wire [7:0] v_22386;
  function [7:0] mux_22386(input [0:0] sel);
    case (sel) 0: mux_22386 = 8'h0; 1: mux_22386 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22387;
  wire [7:0] v_22388;
  wire [7:0] v_22389;
  function [7:0] mux_22389(input [0:0] sel);
    case (sel) 0: mux_22389 = 8'h0; 1: mux_22389 = v_22390;
    endcase
  endfunction
  reg [7:0] v_22390 = 8'h0;
  wire [7:0] v_22391;
  wire [7:0] v_22392;
  function [7:0] mux_22392(input [0:0] sel);
    case (sel) 0: mux_22392 = 8'h0; 1: mux_22392 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22393;
  wire [7:0] v_22394;
  wire [7:0] v_22395;
  function [7:0] mux_22395(input [0:0] sel);
    case (sel) 0: mux_22395 = 8'h0; 1: mux_22395 = v_22396;
    endcase
  endfunction
  reg [7:0] v_22396 = 8'h0;
  wire [7:0] v_22397;
  wire [7:0] v_22398;
  function [7:0] mux_22398(input [0:0] sel);
    case (sel) 0: mux_22398 = 8'h0; 1: mux_22398 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22399;
  wire [7:0] v_22400;
  wire [7:0] v_22401;
  function [7:0] mux_22401(input [0:0] sel);
    case (sel) 0: mux_22401 = 8'h0; 1: mux_22401 = v_22402;
    endcase
  endfunction
  reg [7:0] v_22402 = 8'h0;
  wire [7:0] v_22403;
  wire [7:0] v_22404;
  function [7:0] mux_22404(input [0:0] sel);
    case (sel) 0: mux_22404 = 8'h0; 1: mux_22404 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22405;
  wire [7:0] v_22406;
  wire [7:0] v_22407;
  function [7:0] mux_22407(input [0:0] sel);
    case (sel) 0: mux_22407 = 8'h0; 1: mux_22407 = v_22408;
    endcase
  endfunction
  reg [7:0] v_22408 = 8'h0;
  wire [7:0] v_22409;
  wire [7:0] v_22410;
  function [7:0] mux_22410(input [0:0] sel);
    case (sel) 0: mux_22410 = 8'h0; 1: mux_22410 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22411;
  wire [7:0] v_22412;
  wire [7:0] v_22413;
  function [7:0] mux_22413(input [0:0] sel);
    case (sel) 0: mux_22413 = 8'h0; 1: mux_22413 = v_22414;
    endcase
  endfunction
  reg [7:0] v_22414 = 8'h0;
  wire [7:0] v_22415;
  wire [7:0] v_22416;
  function [7:0] mux_22416(input [0:0] sel);
    case (sel) 0: mux_22416 = 8'h0; 1: mux_22416 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22417;
  wire [7:0] v_22418;
  wire [7:0] v_22419;
  function [7:0] mux_22419(input [0:0] sel);
    case (sel) 0: mux_22419 = 8'h0; 1: mux_22419 = v_22420;
    endcase
  endfunction
  reg [7:0] v_22420 = 8'h0;
  wire [7:0] v_22421;
  wire [7:0] v_22422;
  function [7:0] mux_22422(input [0:0] sel);
    case (sel) 0: mux_22422 = 8'h0; 1: mux_22422 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22423;
  wire [7:0] v_22424;
  wire [7:0] v_22425;
  function [7:0] mux_22425(input [0:0] sel);
    case (sel) 0: mux_22425 = 8'h0; 1: mux_22425 = v_22426;
    endcase
  endfunction
  reg [7:0] v_22426 = 8'h0;
  wire [7:0] v_22427;
  wire [7:0] v_22428;
  function [7:0] mux_22428(input [0:0] sel);
    case (sel) 0: mux_22428 = 8'h0; 1: mux_22428 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22429;
  wire [7:0] v_22430;
  wire [7:0] v_22431;
  function [7:0] mux_22431(input [0:0] sel);
    case (sel) 0: mux_22431 = 8'h0; 1: mux_22431 = v_22432;
    endcase
  endfunction
  reg [7:0] v_22432 = 8'h0;
  wire [7:0] v_22433;
  wire [7:0] v_22434;
  function [7:0] mux_22434(input [0:0] sel);
    case (sel) 0: mux_22434 = 8'h0; 1: mux_22434 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22435;
  wire [7:0] v_22436;
  wire [7:0] v_22437;
  function [7:0] mux_22437(input [0:0] sel);
    case (sel) 0: mux_22437 = 8'h0; 1: mux_22437 = v_22438;
    endcase
  endfunction
  reg [7:0] v_22438 = 8'h0;
  wire [7:0] v_22439;
  wire [7:0] v_22440;
  function [7:0] mux_22440(input [0:0] sel);
    case (sel) 0: mux_22440 = 8'h0; 1: mux_22440 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22441;
  wire [7:0] v_22442;
  wire [7:0] v_22443;
  function [7:0] mux_22443(input [0:0] sel);
    case (sel) 0: mux_22443 = 8'h0; 1: mux_22443 = vout_peek_22178;
    endcase
  endfunction
  wire [7:0] v_22444;
  function [7:0] mux_22444(input [0:0] sel);
    case (sel) 0: mux_22444 = 8'h0; 1: mux_22444 = vout_peek_22169;
    endcase
  endfunction
  wire [7:0] v_22445;
  function [7:0] mux_22445(input [0:0] sel);
    case (sel) 0: mux_22445 = 8'h0; 1: mux_22445 = v_22446;
    endcase
  endfunction
  reg [7:0] v_22446 = 8'h0;
  wire [7:0] v_22447;
  wire [7:0] v_22448;
  function [7:0] mux_22448(input [0:0] sel);
    case (sel) 0: mux_22448 = 8'h0; 1: mux_22448 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22449;
  wire [7:0] v_22450;
  wire [7:0] v_22451;
  function [7:0] mux_22451(input [0:0] sel);
    case (sel) 0: mux_22451 = 8'h0; 1: mux_22451 = vout_peek_22141;
    endcase
  endfunction
  wire [7:0] v_22452;
  function [7:0] mux_22452(input [0:0] sel);
    case (sel) 0: mux_22452 = 8'h0; 1: mux_22452 = vout_peek_22132;
    endcase
  endfunction
  wire [7:0] v_22453;
  function [7:0] mux_22453(input [0:0] sel);
    case (sel) 0: mux_22453 = 8'h0; 1: mux_22453 = v_22454;
    endcase
  endfunction
  reg [7:0] v_22454 = 8'h0;
  wire [7:0] v_22455;
  wire [7:0] v_22456;
  function [7:0] mux_22456(input [0:0] sel);
    case (sel) 0: mux_22456 = 8'h0; 1: mux_22456 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22457;
  wire [7:0] v_22458;
  wire [7:0] v_22459;
  function [7:0] mux_22459(input [0:0] sel);
    case (sel) 0: mux_22459 = 8'h0; 1: mux_22459 = v_22460;
    endcase
  endfunction
  reg [7:0] v_22460 = 8'h0;
  wire [7:0] v_22461;
  wire [7:0] v_22462;
  function [7:0] mux_22462(input [0:0] sel);
    case (sel) 0: mux_22462 = 8'h0; 1: mux_22462 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22463;
  wire [7:0] v_22464;
  wire [7:0] v_22465;
  function [7:0] mux_22465(input [0:0] sel);
    case (sel) 0: mux_22465 = 8'h0; 1: mux_22465 = vout_peek_22085;
    endcase
  endfunction
  wire [7:0] v_22466;
  function [7:0] mux_22466(input [0:0] sel);
    case (sel) 0: mux_22466 = 8'h0; 1: mux_22466 = vout_peek_22076;
    endcase
  endfunction
  wire [7:0] v_22467;
  function [7:0] mux_22467(input [0:0] sel);
    case (sel) 0: mux_22467 = 8'h0; 1: mux_22467 = v_22468;
    endcase
  endfunction
  reg [7:0] v_22468 = 8'h0;
  wire [7:0] v_22469;
  wire [7:0] v_22470;
  function [7:0] mux_22470(input [0:0] sel);
    case (sel) 0: mux_22470 = 8'h0; 1: mux_22470 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22471;
  wire [7:0] v_22472;
  wire [7:0] v_22473;
  function [7:0] mux_22473(input [0:0] sel);
    case (sel) 0: mux_22473 = 8'h0; 1: mux_22473 = vout_peek_22048;
    endcase
  endfunction
  wire [7:0] v_22474;
  function [7:0] mux_22474(input [0:0] sel);
    case (sel) 0: mux_22474 = 8'h0; 1: mux_22474 = vout_peek_22039;
    endcase
  endfunction
  wire [7:0] v_22475;
  function [7:0] mux_22475(input [0:0] sel);
    case (sel) 0: mux_22475 = 8'h0; 1: mux_22475 = v_22476;
    endcase
  endfunction
  reg [7:0] v_22476 = 8'h0;
  wire [7:0] v_22477;
  wire [7:0] v_22478;
  function [7:0] mux_22478(input [0:0] sel);
    case (sel) 0: mux_22478 = 8'h0; 1: mux_22478 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22479;
  wire [7:0] v_22480;
  wire [7:0] v_22481;
  function [7:0] mux_22481(input [0:0] sel);
    case (sel) 0: mux_22481 = 8'h0; 1: mux_22481 = v_22482;
    endcase
  endfunction
  reg [7:0] v_22482 = 8'h0;
  wire [7:0] v_22483;
  wire [7:0] v_22484;
  function [7:0] mux_22484(input [0:0] sel);
    case (sel) 0: mux_22484 = 8'h0; 1: mux_22484 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22485;
  wire [7:0] v_22486;
  wire [7:0] v_22487;
  function [7:0] mux_22487(input [0:0] sel);
    case (sel) 0: mux_22487 = 8'h0; 1: mux_22487 = v_22488;
    endcase
  endfunction
  reg [7:0] v_22488 = 8'h0;
  wire [7:0] v_22489;
  wire [7:0] v_22490;
  function [7:0] mux_22490(input [0:0] sel);
    case (sel) 0: mux_22490 = 8'h0; 1: mux_22490 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22491;
  wire [7:0] v_22492;
  wire [7:0] v_22493;
  function [7:0] mux_22493(input [0:0] sel);
    case (sel) 0: mux_22493 = 8'h0; 1: mux_22493 = vout_peek_21973;
    endcase
  endfunction
  wire [7:0] v_22494;
  function [7:0] mux_22494(input [0:0] sel);
    case (sel) 0: mux_22494 = 8'h0; 1: mux_22494 = vout_peek_21964;
    endcase
  endfunction
  wire [7:0] v_22495;
  function [7:0] mux_22495(input [0:0] sel);
    case (sel) 0: mux_22495 = 8'h0; 1: mux_22495 = v_22496;
    endcase
  endfunction
  reg [7:0] v_22496 = 8'h0;
  wire [7:0] v_22497;
  wire [7:0] v_22498;
  function [7:0] mux_22498(input [0:0] sel);
    case (sel) 0: mux_22498 = 8'h0; 1: mux_22498 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22499;
  wire [7:0] v_22500;
  wire [7:0] v_22501;
  function [7:0] mux_22501(input [0:0] sel);
    case (sel) 0: mux_22501 = 8'h0; 1: mux_22501 = vout_peek_21936;
    endcase
  endfunction
  wire [7:0] v_22502;
  function [7:0] mux_22502(input [0:0] sel);
    case (sel) 0: mux_22502 = 8'h0; 1: mux_22502 = vout_peek_21927;
    endcase
  endfunction
  wire [7:0] v_22503;
  function [7:0] mux_22503(input [0:0] sel);
    case (sel) 0: mux_22503 = 8'h0; 1: mux_22503 = v_22504;
    endcase
  endfunction
  reg [7:0] v_22504 = 8'h0;
  wire [7:0] v_22505;
  wire [7:0] v_22506;
  function [7:0] mux_22506(input [0:0] sel);
    case (sel) 0: mux_22506 = 8'h0; 1: mux_22506 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22507;
  wire [7:0] v_22508;
  wire [7:0] v_22509;
  function [7:0] mux_22509(input [0:0] sel);
    case (sel) 0: mux_22509 = 8'h0; 1: mux_22509 = v_22510;
    endcase
  endfunction
  reg [7:0] v_22510 = 8'h0;
  wire [7:0] v_22511;
  wire [7:0] v_22512;
  function [7:0] mux_22512(input [0:0] sel);
    case (sel) 0: mux_22512 = 8'h0; 1: mux_22512 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22513;
  wire [7:0] v_22514;
  wire [7:0] v_22515;
  function [7:0] mux_22515(input [0:0] sel);
    case (sel) 0: mux_22515 = 8'h0; 1: mux_22515 = vout_peek_21880;
    endcase
  endfunction
  wire [7:0] v_22516;
  function [7:0] mux_22516(input [0:0] sel);
    case (sel) 0: mux_22516 = 8'h0; 1: mux_22516 = vout_peek_21871;
    endcase
  endfunction
  wire [7:0] v_22517;
  function [7:0] mux_22517(input [0:0] sel);
    case (sel) 0: mux_22517 = 8'h0; 1: mux_22517 = v_22518;
    endcase
  endfunction
  reg [7:0] v_22518 = 8'h0;
  wire [7:0] v_22519;
  wire [7:0] v_22520;
  function [7:0] mux_22520(input [0:0] sel);
    case (sel) 0: mux_22520 = 8'h0; 1: mux_22520 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22521;
  wire [7:0] v_22522;
  wire [7:0] v_22523;
  function [7:0] mux_22523(input [0:0] sel);
    case (sel) 0: mux_22523 = 8'h0; 1: mux_22523 = vout_peek_21843;
    endcase
  endfunction
  wire [7:0] v_22524;
  function [7:0] mux_22524(input [0:0] sel);
    case (sel) 0: mux_22524 = 8'h0; 1: mux_22524 = vout_peek_21834;
    endcase
  endfunction
  wire [7:0] v_22525;
  function [7:0] mux_22525(input [0:0] sel);
    case (sel) 0: mux_22525 = 8'h0; 1: mux_22525 = v_22526;
    endcase
  endfunction
  reg [7:0] v_22526 = 8'h0;
  wire [7:0] v_22527;
  wire [7:0] v_22528;
  function [7:0] mux_22528(input [0:0] sel);
    case (sel) 0: mux_22528 = 8'h0; 1: mux_22528 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22529;
  wire [7:0] v_22530;
  wire [7:0] v_22531;
  function [7:0] mux_22531(input [0:0] sel);
    case (sel) 0: mux_22531 = 8'h0; 1: mux_22531 = v_22532;
    endcase
  endfunction
  reg [7:0] v_22532 = 8'h0;
  wire [7:0] v_22533;
  wire [7:0] v_22534;
  function [7:0] mux_22534(input [0:0] sel);
    case (sel) 0: mux_22534 = 8'h0; 1: mux_22534 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22535;
  wire [7:0] v_22536;
  wire [7:0] v_22537;
  function [7:0] mux_22537(input [0:0] sel);
    case (sel) 0: mux_22537 = 8'h0; 1: mux_22537 = v_22538;
    endcase
  endfunction
  reg [7:0] v_22538 = 8'h0;
  wire [7:0] v_22539;
  wire [7:0] v_22540;
  function [7:0] mux_22540(input [0:0] sel);
    case (sel) 0: mux_22540 = 8'h0; 1: mux_22540 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22541;
  wire [7:0] v_22542;
  wire [7:0] v_22543;
  function [7:0] mux_22543(input [0:0] sel);
    case (sel) 0: mux_22543 = 8'h0; 1: mux_22543 = v_22544;
    endcase
  endfunction
  reg [7:0] v_22544 = 8'h0;
  wire [7:0] v_22545;
  wire [7:0] v_22546;
  function [7:0] mux_22546(input [0:0] sel);
    case (sel) 0: mux_22546 = 8'h0; 1: mux_22546 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22547;
  wire [7:0] v_22548;
  wire [7:0] v_22549;
  function [7:0] mux_22549(input [0:0] sel);
    case (sel) 0: mux_22549 = 8'h0; 1: mux_22549 = vout_peek_21749;
    endcase
  endfunction
  wire [7:0] v_22550;
  function [7:0] mux_22550(input [0:0] sel);
    case (sel) 0: mux_22550 = 8'h0; 1: mux_22550 = vout_peek_21740;
    endcase
  endfunction
  wire [7:0] v_22551;
  function [7:0] mux_22551(input [0:0] sel);
    case (sel) 0: mux_22551 = 8'h0; 1: mux_22551 = v_22552;
    endcase
  endfunction
  reg [7:0] v_22552 = 8'h0;
  wire [7:0] v_22553;
  wire [7:0] v_22554;
  function [7:0] mux_22554(input [0:0] sel);
    case (sel) 0: mux_22554 = 8'h0; 1: mux_22554 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22555;
  wire [7:0] v_22556;
  wire [7:0] v_22557;
  function [7:0] mux_22557(input [0:0] sel);
    case (sel) 0: mux_22557 = 8'h0; 1: mux_22557 = vout_peek_21712;
    endcase
  endfunction
  wire [7:0] v_22558;
  function [7:0] mux_22558(input [0:0] sel);
    case (sel) 0: mux_22558 = 8'h0; 1: mux_22558 = vout_peek_21703;
    endcase
  endfunction
  wire [7:0] v_22559;
  function [7:0] mux_22559(input [0:0] sel);
    case (sel) 0: mux_22559 = 8'h0; 1: mux_22559 = v_22560;
    endcase
  endfunction
  reg [7:0] v_22560 = 8'h0;
  wire [7:0] v_22561;
  wire [7:0] v_22562;
  function [7:0] mux_22562(input [0:0] sel);
    case (sel) 0: mux_22562 = 8'h0; 1: mux_22562 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22563;
  wire [7:0] v_22564;
  wire [7:0] v_22565;
  function [7:0] mux_22565(input [0:0] sel);
    case (sel) 0: mux_22565 = 8'h0; 1: mux_22565 = v_22566;
    endcase
  endfunction
  reg [7:0] v_22566 = 8'h0;
  wire [7:0] v_22567;
  wire [7:0] v_22568;
  function [7:0] mux_22568(input [0:0] sel);
    case (sel) 0: mux_22568 = 8'h0; 1: mux_22568 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22569;
  wire [7:0] v_22570;
  wire [7:0] v_22571;
  function [7:0] mux_22571(input [0:0] sel);
    case (sel) 0: mux_22571 = 8'h0; 1: mux_22571 = vout_peek_21656;
    endcase
  endfunction
  wire [7:0] v_22572;
  function [7:0] mux_22572(input [0:0] sel);
    case (sel) 0: mux_22572 = 8'h0; 1: mux_22572 = vout_peek_21647;
    endcase
  endfunction
  wire [7:0] v_22573;
  function [7:0] mux_22573(input [0:0] sel);
    case (sel) 0: mux_22573 = 8'h0; 1: mux_22573 = v_22574;
    endcase
  endfunction
  reg [7:0] v_22574 = 8'h0;
  wire [7:0] v_22575;
  wire [7:0] v_22576;
  function [7:0] mux_22576(input [0:0] sel);
    case (sel) 0: mux_22576 = 8'h0; 1: mux_22576 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22577;
  wire [7:0] v_22578;
  wire [7:0] v_22579;
  function [7:0] mux_22579(input [0:0] sel);
    case (sel) 0: mux_22579 = 8'h0; 1: mux_22579 = vout_peek_21619;
    endcase
  endfunction
  wire [7:0] v_22580;
  function [7:0] mux_22580(input [0:0] sel);
    case (sel) 0: mux_22580 = 8'h0; 1: mux_22580 = vout_peek_21610;
    endcase
  endfunction
  wire [7:0] v_22581;
  function [7:0] mux_22581(input [0:0] sel);
    case (sel) 0: mux_22581 = 8'h0; 1: mux_22581 = v_22582;
    endcase
  endfunction
  reg [7:0] v_22582 = 8'h0;
  wire [7:0] v_22583;
  wire [7:0] v_22584;
  function [7:0] mux_22584(input [0:0] sel);
    case (sel) 0: mux_22584 = 8'h0; 1: mux_22584 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22585;
  wire [7:0] v_22586;
  wire [7:0] v_22587;
  function [7:0] mux_22587(input [0:0] sel);
    case (sel) 0: mux_22587 = 8'h0; 1: mux_22587 = v_22588;
    endcase
  endfunction
  reg [7:0] v_22588 = 8'h0;
  wire [7:0] v_22589;
  wire [7:0] v_22590;
  function [7:0] mux_22590(input [0:0] sel);
    case (sel) 0: mux_22590 = 8'h0; 1: mux_22590 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22591;
  wire [7:0] v_22592;
  wire [7:0] v_22593;
  function [7:0] mux_22593(input [0:0] sel);
    case (sel) 0: mux_22593 = 8'h0; 1: mux_22593 = v_22594;
    endcase
  endfunction
  reg [7:0] v_22594 = 8'h0;
  wire [7:0] v_22595;
  wire [7:0] v_22596;
  function [7:0] mux_22596(input [0:0] sel);
    case (sel) 0: mux_22596 = 8'h0; 1: mux_22596 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22597;
  wire [7:0] v_22598;
  wire [7:0] v_22599;
  function [7:0] mux_22599(input [0:0] sel);
    case (sel) 0: mux_22599 = 8'h0; 1: mux_22599 = vout_peek_21544;
    endcase
  endfunction
  wire [7:0] v_22600;
  function [7:0] mux_22600(input [0:0] sel);
    case (sel) 0: mux_22600 = 8'h0; 1: mux_22600 = vout_peek_21535;
    endcase
  endfunction
  wire [7:0] v_22601;
  function [7:0] mux_22601(input [0:0] sel);
    case (sel) 0: mux_22601 = 8'h0; 1: mux_22601 = v_22602;
    endcase
  endfunction
  reg [7:0] v_22602 = 8'h0;
  wire [7:0] v_22603;
  wire [7:0] v_22604;
  function [7:0] mux_22604(input [0:0] sel);
    case (sel) 0: mux_22604 = 8'h0; 1: mux_22604 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22605;
  wire [7:0] v_22606;
  wire [7:0] v_22607;
  function [7:0] mux_22607(input [0:0] sel);
    case (sel) 0: mux_22607 = 8'h0; 1: mux_22607 = vout_peek_21507;
    endcase
  endfunction
  wire [7:0] v_22608;
  function [7:0] mux_22608(input [0:0] sel);
    case (sel) 0: mux_22608 = 8'h0; 1: mux_22608 = vout_peek_21498;
    endcase
  endfunction
  wire [7:0] v_22609;
  function [7:0] mux_22609(input [0:0] sel);
    case (sel) 0: mux_22609 = 8'h0; 1: mux_22609 = v_22610;
    endcase
  endfunction
  reg [7:0] v_22610 = 8'h0;
  wire [7:0] v_22611;
  wire [7:0] v_22612;
  function [7:0] mux_22612(input [0:0] sel);
    case (sel) 0: mux_22612 = 8'h0; 1: mux_22612 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22613;
  wire [7:0] v_22614;
  wire [7:0] v_22615;
  function [7:0] mux_22615(input [0:0] sel);
    case (sel) 0: mux_22615 = 8'h0; 1: mux_22615 = v_22616;
    endcase
  endfunction
  reg [7:0] v_22616 = 8'h0;
  wire [7:0] v_22617;
  wire [7:0] v_22618;
  function [7:0] mux_22618(input [0:0] sel);
    case (sel) 0: mux_22618 = 8'h0; 1: mux_22618 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22619;
  wire [7:0] v_22620;
  wire [7:0] v_22621;
  function [7:0] mux_22621(input [0:0] sel);
    case (sel) 0: mux_22621 = 8'h0; 1: mux_22621 = vout_peek_21451;
    endcase
  endfunction
  wire [7:0] v_22622;
  function [7:0] mux_22622(input [0:0] sel);
    case (sel) 0: mux_22622 = 8'h0; 1: mux_22622 = vout_peek_21442;
    endcase
  endfunction
  wire [7:0] v_22623;
  function [7:0] mux_22623(input [0:0] sel);
    case (sel) 0: mux_22623 = 8'h0; 1: mux_22623 = v_22624;
    endcase
  endfunction
  reg [7:0] v_22624 = 8'h0;
  wire [7:0] v_22625;
  wire [7:0] v_22626;
  function [7:0] mux_22626(input [0:0] sel);
    case (sel) 0: mux_22626 = 8'h0; 1: mux_22626 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22627;
  wire [7:0] v_22628;
  wire [7:0] v_22629;
  function [7:0] mux_22629(input [0:0] sel);
    case (sel) 0: mux_22629 = 8'h0; 1: mux_22629 = vout_peek_21414;
    endcase
  endfunction
  wire [7:0] v_22630;
  function [7:0] mux_22630(input [0:0] sel);
    case (sel) 0: mux_22630 = 8'h0; 1: mux_22630 = vout_peek_21405;
    endcase
  endfunction
  wire [7:0] v_22631;
  function [7:0] mux_22631(input [0:0] sel);
    case (sel) 0: mux_22631 = 8'h0; 1: mux_22631 = v_22632;
    endcase
  endfunction
  reg [7:0] v_22632 = 8'h0;
  wire [7:0] v_22633;
  wire [7:0] v_22634;
  function [7:0] mux_22634(input [0:0] sel);
    case (sel) 0: mux_22634 = 8'h0; 1: mux_22634 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22635;
  wire [7:0] v_22636;
  wire [7:0] v_22637;
  function [7:0] mux_22637(input [0:0] sel);
    case (sel) 0: mux_22637 = 8'h0; 1: mux_22637 = v_22638;
    endcase
  endfunction
  reg [7:0] v_22638 = 8'h0;
  wire [7:0] v_22639;
  wire [7:0] v_22640;
  function [7:0] mux_22640(input [0:0] sel);
    case (sel) 0: mux_22640 = 8'h0; 1: mux_22640 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22641;
  wire [7:0] v_22642;
  wire [7:0] v_22643;
  function [7:0] mux_22643(input [0:0] sel);
    case (sel) 0: mux_22643 = 8'h0; 1: mux_22643 = v_22644;
    endcase
  endfunction
  reg [7:0] v_22644 = 8'h0;
  wire [7:0] v_22645;
  wire [7:0] v_22646;
  function [7:0] mux_22646(input [0:0] sel);
    case (sel) 0: mux_22646 = 8'h0; 1: mux_22646 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22647;
  wire [7:0] v_22648;
  wire [7:0] v_22649;
  function [7:0] mux_22649(input [0:0] sel);
    case (sel) 0: mux_22649 = 8'h0; 1: mux_22649 = v_22650;
    endcase
  endfunction
  reg [7:0] v_22650 = 8'h0;
  wire [7:0] v_22651;
  wire [7:0] v_22652;
  function [7:0] mux_22652(input [0:0] sel);
    case (sel) 0: mux_22652 = 8'h0; 1: mux_22652 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22653;
  wire [7:0] v_22654;
  wire [7:0] v_22655;
  function [7:0] mux_22655(input [0:0] sel);
    case (sel) 0: mux_22655 = 8'h0; 1: mux_22655 = v_22656;
    endcase
  endfunction
  reg [7:0] v_22656 = 8'h0;
  wire [7:0] v_22657;
  wire [7:0] v_22658;
  function [7:0] mux_22658(input [0:0] sel);
    case (sel) 0: mux_22658 = 8'h0; 1: mux_22658 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22659;
  wire [7:0] v_22660;
  wire [7:0] v_22661;
  function [7:0] mux_22661(input [0:0] sel);
    case (sel) 0: mux_22661 = 8'h0; 1: mux_22661 = vout_peek_21301;
    endcase
  endfunction
  wire [7:0] v_22662;
  function [7:0] mux_22662(input [0:0] sel);
    case (sel) 0: mux_22662 = 8'h0; 1: mux_22662 = vout_peek_21292;
    endcase
  endfunction
  wire [7:0] v_22663;
  function [7:0] mux_22663(input [0:0] sel);
    case (sel) 0: mux_22663 = 8'h0; 1: mux_22663 = v_22664;
    endcase
  endfunction
  reg [7:0] v_22664 = 8'h0;
  wire [7:0] v_22665;
  wire [7:0] v_22666;
  function [7:0] mux_22666(input [0:0] sel);
    case (sel) 0: mux_22666 = 8'h0; 1: mux_22666 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22667;
  wire [7:0] v_22668;
  wire [7:0] v_22669;
  function [7:0] mux_22669(input [0:0] sel);
    case (sel) 0: mux_22669 = 8'h0; 1: mux_22669 = vout_peek_21264;
    endcase
  endfunction
  wire [7:0] v_22670;
  function [7:0] mux_22670(input [0:0] sel);
    case (sel) 0: mux_22670 = 8'h0; 1: mux_22670 = vout_peek_21255;
    endcase
  endfunction
  wire [7:0] v_22671;
  function [7:0] mux_22671(input [0:0] sel);
    case (sel) 0: mux_22671 = 8'h0; 1: mux_22671 = v_22672;
    endcase
  endfunction
  reg [7:0] v_22672 = 8'h0;
  wire [7:0] v_22673;
  wire [7:0] v_22674;
  function [7:0] mux_22674(input [0:0] sel);
    case (sel) 0: mux_22674 = 8'h0; 1: mux_22674 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22675;
  wire [7:0] v_22676;
  wire [7:0] v_22677;
  function [7:0] mux_22677(input [0:0] sel);
    case (sel) 0: mux_22677 = 8'h0; 1: mux_22677 = v_22678;
    endcase
  endfunction
  reg [7:0] v_22678 = 8'h0;
  wire [7:0] v_22679;
  wire [7:0] v_22680;
  function [7:0] mux_22680(input [0:0] sel);
    case (sel) 0: mux_22680 = 8'h0; 1: mux_22680 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22681;
  wire [7:0] v_22682;
  wire [7:0] v_22683;
  function [7:0] mux_22683(input [0:0] sel);
    case (sel) 0: mux_22683 = 8'h0; 1: mux_22683 = vout_peek_21208;
    endcase
  endfunction
  wire [7:0] v_22684;
  function [7:0] mux_22684(input [0:0] sel);
    case (sel) 0: mux_22684 = 8'h0; 1: mux_22684 = vout_peek_21199;
    endcase
  endfunction
  wire [7:0] v_22685;
  function [7:0] mux_22685(input [0:0] sel);
    case (sel) 0: mux_22685 = 8'h0; 1: mux_22685 = v_22686;
    endcase
  endfunction
  reg [7:0] v_22686 = 8'h0;
  wire [7:0] v_22687;
  wire [7:0] v_22688;
  function [7:0] mux_22688(input [0:0] sel);
    case (sel) 0: mux_22688 = 8'h0; 1: mux_22688 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22689;
  wire [7:0] v_22690;
  wire [7:0] v_22691;
  function [7:0] mux_22691(input [0:0] sel);
    case (sel) 0: mux_22691 = 8'h0; 1: mux_22691 = vout_peek_21171;
    endcase
  endfunction
  wire [7:0] v_22692;
  function [7:0] mux_22692(input [0:0] sel);
    case (sel) 0: mux_22692 = 8'h0; 1: mux_22692 = vout_peek_21162;
    endcase
  endfunction
  wire [7:0] v_22693;
  function [7:0] mux_22693(input [0:0] sel);
    case (sel) 0: mux_22693 = 8'h0; 1: mux_22693 = v_22694;
    endcase
  endfunction
  reg [7:0] v_22694 = 8'h0;
  wire [7:0] v_22695;
  wire [7:0] v_22696;
  function [7:0] mux_22696(input [0:0] sel);
    case (sel) 0: mux_22696 = 8'h0; 1: mux_22696 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22697;
  wire [7:0] v_22698;
  wire [7:0] v_22699;
  function [7:0] mux_22699(input [0:0] sel);
    case (sel) 0: mux_22699 = 8'h0; 1: mux_22699 = v_22700;
    endcase
  endfunction
  reg [7:0] v_22700 = 8'h0;
  wire [7:0] v_22701;
  wire [7:0] v_22702;
  function [7:0] mux_22702(input [0:0] sel);
    case (sel) 0: mux_22702 = 8'h0; 1: mux_22702 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22703;
  wire [7:0] v_22704;
  wire [7:0] v_22705;
  function [7:0] mux_22705(input [0:0] sel);
    case (sel) 0: mux_22705 = 8'h0; 1: mux_22705 = v_22706;
    endcase
  endfunction
  reg [7:0] v_22706 = 8'h0;
  wire [7:0] v_22707;
  wire [7:0] v_22708;
  function [7:0] mux_22708(input [0:0] sel);
    case (sel) 0: mux_22708 = 8'h0; 1: mux_22708 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22709;
  wire [7:0] v_22710;
  wire [7:0] v_22711;
  function [7:0] mux_22711(input [0:0] sel);
    case (sel) 0: mux_22711 = 8'h0; 1: mux_22711 = vout_peek_21096;
    endcase
  endfunction
  wire [7:0] v_22712;
  function [7:0] mux_22712(input [0:0] sel);
    case (sel) 0: mux_22712 = 8'h0; 1: mux_22712 = vout_peek_21087;
    endcase
  endfunction
  wire [7:0] v_22713;
  function [7:0] mux_22713(input [0:0] sel);
    case (sel) 0: mux_22713 = 8'h0; 1: mux_22713 = v_22714;
    endcase
  endfunction
  reg [7:0] v_22714 = 8'h0;
  wire [7:0] v_22715;
  wire [7:0] v_22716;
  function [7:0] mux_22716(input [0:0] sel);
    case (sel) 0: mux_22716 = 8'h0; 1: mux_22716 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22717;
  wire [7:0] v_22718;
  wire [7:0] v_22719;
  function [7:0] mux_22719(input [0:0] sel);
    case (sel) 0: mux_22719 = 8'h0; 1: mux_22719 = vout_peek_21059;
    endcase
  endfunction
  wire [7:0] v_22720;
  function [7:0] mux_22720(input [0:0] sel);
    case (sel) 0: mux_22720 = 8'h0; 1: mux_22720 = vout_peek_21050;
    endcase
  endfunction
  wire [7:0] v_22721;
  function [7:0] mux_22721(input [0:0] sel);
    case (sel) 0: mux_22721 = 8'h0; 1: mux_22721 = v_22722;
    endcase
  endfunction
  reg [7:0] v_22722 = 8'h0;
  wire [7:0] v_22723;
  wire [7:0] v_22724;
  function [7:0] mux_22724(input [0:0] sel);
    case (sel) 0: mux_22724 = 8'h0; 1: mux_22724 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22725;
  wire [7:0] v_22726;
  wire [7:0] v_22727;
  function [7:0] mux_22727(input [0:0] sel);
    case (sel) 0: mux_22727 = 8'h0; 1: mux_22727 = v_22728;
    endcase
  endfunction
  reg [7:0] v_22728 = 8'h0;
  wire [7:0] v_22729;
  wire [7:0] v_22730;
  function [7:0] mux_22730(input [0:0] sel);
    case (sel) 0: mux_22730 = 8'h0; 1: mux_22730 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22731;
  wire [7:0] v_22732;
  wire [7:0] v_22733;
  function [7:0] mux_22733(input [0:0] sel);
    case (sel) 0: mux_22733 = 8'h0; 1: mux_22733 = vout_peek_21003;
    endcase
  endfunction
  wire [7:0] v_22734;
  function [7:0] mux_22734(input [0:0] sel);
    case (sel) 0: mux_22734 = 8'h0; 1: mux_22734 = vout_peek_20994;
    endcase
  endfunction
  wire [7:0] v_22735;
  function [7:0] mux_22735(input [0:0] sel);
    case (sel) 0: mux_22735 = 8'h0; 1: mux_22735 = v_22736;
    endcase
  endfunction
  reg [7:0] v_22736 = 8'h0;
  wire [7:0] v_22737;
  wire [7:0] v_22738;
  function [7:0] mux_22738(input [0:0] sel);
    case (sel) 0: mux_22738 = 8'h0; 1: mux_22738 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22739;
  wire [7:0] v_22740;
  wire [7:0] v_22741;
  function [7:0] mux_22741(input [0:0] sel);
    case (sel) 0: mux_22741 = 8'h0; 1: mux_22741 = vout_peek_20966;
    endcase
  endfunction
  wire [7:0] v_22742;
  function [7:0] mux_22742(input [0:0] sel);
    case (sel) 0: mux_22742 = 8'h0; 1: mux_22742 = vout_peek_20957;
    endcase
  endfunction
  wire [7:0] v_22743;
  function [7:0] mux_22743(input [0:0] sel);
    case (sel) 0: mux_22743 = 8'h0; 1: mux_22743 = v_22744;
    endcase
  endfunction
  reg [7:0] v_22744 = 8'h0;
  wire [7:0] v_22745;
  wire [7:0] v_22746;
  function [7:0] mux_22746(input [0:0] sel);
    case (sel) 0: mux_22746 = 8'h0; 1: mux_22746 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22747;
  wire [7:0] v_22748;
  wire [7:0] v_22749;
  function [7:0] mux_22749(input [0:0] sel);
    case (sel) 0: mux_22749 = 8'h0; 1: mux_22749 = v_22750;
    endcase
  endfunction
  reg [7:0] v_22750 = 8'h0;
  wire [7:0] v_22751;
  wire [7:0] v_22752;
  function [7:0] mux_22752(input [0:0] sel);
    case (sel) 0: mux_22752 = 8'h0; 1: mux_22752 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22753;
  wire [7:0] v_22754;
  wire [7:0] v_22755;
  function [7:0] mux_22755(input [0:0] sel);
    case (sel) 0: mux_22755 = 8'h0; 1: mux_22755 = v_22756;
    endcase
  endfunction
  reg [7:0] v_22756 = 8'h0;
  wire [7:0] v_22757;
  wire [7:0] v_22758;
  function [7:0] mux_22758(input [0:0] sel);
    case (sel) 0: mux_22758 = 8'h0; 1: mux_22758 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22759;
  wire [7:0] v_22760;
  wire [7:0] v_22761;
  function [7:0] mux_22761(input [0:0] sel);
    case (sel) 0: mux_22761 = 8'h0; 1: mux_22761 = v_22762;
    endcase
  endfunction
  reg [7:0] v_22762 = 8'h0;
  wire [7:0] v_22763;
  wire [7:0] v_22764;
  function [7:0] mux_22764(input [0:0] sel);
    case (sel) 0: mux_22764 = 8'h0; 1: mux_22764 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22765;
  wire [7:0] v_22766;
  wire [7:0] v_22767;
  function [7:0] mux_22767(input [0:0] sel);
    case (sel) 0: mux_22767 = 8'h0; 1: mux_22767 = vout_peek_20872;
    endcase
  endfunction
  wire [7:0] v_22768;
  function [7:0] mux_22768(input [0:0] sel);
    case (sel) 0: mux_22768 = 8'h0; 1: mux_22768 = vout_peek_20863;
    endcase
  endfunction
  wire [7:0] v_22769;
  function [7:0] mux_22769(input [0:0] sel);
    case (sel) 0: mux_22769 = 8'h0; 1: mux_22769 = v_22770;
    endcase
  endfunction
  reg [7:0] v_22770 = 8'h0;
  wire [7:0] v_22771;
  wire [7:0] v_22772;
  function [7:0] mux_22772(input [0:0] sel);
    case (sel) 0: mux_22772 = 8'h0; 1: mux_22772 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22773;
  wire [7:0] v_22774;
  wire [7:0] v_22775;
  function [7:0] mux_22775(input [0:0] sel);
    case (sel) 0: mux_22775 = 8'h0; 1: mux_22775 = vout_peek_20835;
    endcase
  endfunction
  wire [7:0] v_22776;
  function [7:0] mux_22776(input [0:0] sel);
    case (sel) 0: mux_22776 = 8'h0; 1: mux_22776 = vout_peek_20826;
    endcase
  endfunction
  wire [7:0] v_22777;
  function [7:0] mux_22777(input [0:0] sel);
    case (sel) 0: mux_22777 = 8'h0; 1: mux_22777 = v_22778;
    endcase
  endfunction
  reg [7:0] v_22778 = 8'h0;
  wire [7:0] v_22779;
  wire [7:0] v_22780;
  function [7:0] mux_22780(input [0:0] sel);
    case (sel) 0: mux_22780 = 8'h0; 1: mux_22780 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22781;
  wire [7:0] v_22782;
  wire [7:0] v_22783;
  function [7:0] mux_22783(input [0:0] sel);
    case (sel) 0: mux_22783 = 8'h0; 1: mux_22783 = v_22784;
    endcase
  endfunction
  reg [7:0] v_22784 = 8'h0;
  wire [7:0] v_22785;
  wire [7:0] v_22786;
  function [7:0] mux_22786(input [0:0] sel);
    case (sel) 0: mux_22786 = 8'h0; 1: mux_22786 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22787;
  wire [7:0] v_22788;
  wire [7:0] v_22789;
  function [7:0] mux_22789(input [0:0] sel);
    case (sel) 0: mux_22789 = 8'h0; 1: mux_22789 = vout_peek_20779;
    endcase
  endfunction
  wire [7:0] v_22790;
  function [7:0] mux_22790(input [0:0] sel);
    case (sel) 0: mux_22790 = 8'h0; 1: mux_22790 = vout_peek_20770;
    endcase
  endfunction
  wire [7:0] v_22791;
  function [7:0] mux_22791(input [0:0] sel);
    case (sel) 0: mux_22791 = 8'h0; 1: mux_22791 = v_22792;
    endcase
  endfunction
  reg [7:0] v_22792 = 8'h0;
  wire [7:0] v_22793;
  wire [7:0] v_22794;
  function [7:0] mux_22794(input [0:0] sel);
    case (sel) 0: mux_22794 = 8'h0; 1: mux_22794 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22795;
  wire [7:0] v_22796;
  wire [7:0] v_22797;
  function [7:0] mux_22797(input [0:0] sel);
    case (sel) 0: mux_22797 = 8'h0; 1: mux_22797 = vout_peek_20742;
    endcase
  endfunction
  wire [7:0] v_22798;
  function [7:0] mux_22798(input [0:0] sel);
    case (sel) 0: mux_22798 = 8'h0; 1: mux_22798 = vout_peek_20733;
    endcase
  endfunction
  wire [7:0] v_22799;
  function [7:0] mux_22799(input [0:0] sel);
    case (sel) 0: mux_22799 = 8'h0; 1: mux_22799 = v_22800;
    endcase
  endfunction
  reg [7:0] v_22800 = 8'h0;
  wire [7:0] v_22801;
  wire [7:0] v_22802;
  function [7:0] mux_22802(input [0:0] sel);
    case (sel) 0: mux_22802 = 8'h0; 1: mux_22802 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22803;
  wire [7:0] v_22804;
  wire [7:0] v_22805;
  function [7:0] mux_22805(input [0:0] sel);
    case (sel) 0: mux_22805 = 8'h0; 1: mux_22805 = v_22806;
    endcase
  endfunction
  reg [7:0] v_22806 = 8'h0;
  wire [7:0] v_22807;
  wire [7:0] v_22808;
  function [7:0] mux_22808(input [0:0] sel);
    case (sel) 0: mux_22808 = 8'h0; 1: mux_22808 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22809;
  wire [7:0] v_22810;
  wire [7:0] v_22811;
  function [7:0] mux_22811(input [0:0] sel);
    case (sel) 0: mux_22811 = 8'h0; 1: mux_22811 = v_22812;
    endcase
  endfunction
  reg [7:0] v_22812 = 8'h0;
  wire [7:0] v_22813;
  wire [7:0] v_22814;
  function [7:0] mux_22814(input [0:0] sel);
    case (sel) 0: mux_22814 = 8'h0; 1: mux_22814 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22815;
  wire [7:0] v_22816;
  wire [7:0] v_22817;
  function [7:0] mux_22817(input [0:0] sel);
    case (sel) 0: mux_22817 = 8'h0; 1: mux_22817 = vout_peek_20667;
    endcase
  endfunction
  wire [7:0] v_22818;
  function [7:0] mux_22818(input [0:0] sel);
    case (sel) 0: mux_22818 = 8'h0; 1: mux_22818 = vout_peek_20658;
    endcase
  endfunction
  wire [7:0] v_22819;
  function [7:0] mux_22819(input [0:0] sel);
    case (sel) 0: mux_22819 = 8'h0; 1: mux_22819 = v_22820;
    endcase
  endfunction
  reg [7:0] v_22820 = 8'h0;
  wire [7:0] v_22821;
  wire [7:0] v_22822;
  function [7:0] mux_22822(input [0:0] sel);
    case (sel) 0: mux_22822 = 8'h0; 1: mux_22822 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22823;
  wire [7:0] v_22824;
  wire [7:0] v_22825;
  function [7:0] mux_22825(input [0:0] sel);
    case (sel) 0: mux_22825 = 8'h0; 1: mux_22825 = vout_peek_20630;
    endcase
  endfunction
  wire [7:0] v_22826;
  function [7:0] mux_22826(input [0:0] sel);
    case (sel) 0: mux_22826 = 8'h0; 1: mux_22826 = vout_peek_20621;
    endcase
  endfunction
  wire [7:0] v_22827;
  function [7:0] mux_22827(input [0:0] sel);
    case (sel) 0: mux_22827 = 8'h0; 1: mux_22827 = v_22828;
    endcase
  endfunction
  reg [7:0] v_22828 = 8'h0;
  wire [7:0] v_22829;
  wire [7:0] v_22830;
  function [7:0] mux_22830(input [0:0] sel);
    case (sel) 0: mux_22830 = 8'h0; 1: mux_22830 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22831;
  wire [7:0] v_22832;
  wire [7:0] v_22833;
  function [7:0] mux_22833(input [0:0] sel);
    case (sel) 0: mux_22833 = 8'h0; 1: mux_22833 = v_22834;
    endcase
  endfunction
  reg [7:0] v_22834 = 8'h0;
  wire [7:0] v_22835;
  wire [7:0] v_22836;
  function [7:0] mux_22836(input [0:0] sel);
    case (sel) 0: mux_22836 = 8'h0; 1: mux_22836 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22837;
  wire [7:0] v_22838;
  wire [7:0] v_22839;
  function [7:0] mux_22839(input [0:0] sel);
    case (sel) 0: mux_22839 = 8'h0; 1: mux_22839 = vout_peek_20574;
    endcase
  endfunction
  wire [7:0] v_22840;
  function [7:0] mux_22840(input [0:0] sel);
    case (sel) 0: mux_22840 = 8'h0; 1: mux_22840 = vout_peek_20565;
    endcase
  endfunction
  wire [7:0] v_22841;
  function [7:0] mux_22841(input [0:0] sel);
    case (sel) 0: mux_22841 = 8'h0; 1: mux_22841 = v_22842;
    endcase
  endfunction
  reg [7:0] v_22842 = 8'h0;
  wire [7:0] v_22843;
  wire [7:0] v_22844;
  function [7:0] mux_22844(input [0:0] sel);
    case (sel) 0: mux_22844 = 8'h0; 1: mux_22844 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22845;
  wire [7:0] v_22846;
  wire [7:0] v_22847;
  function [7:0] mux_22847(input [0:0] sel);
    case (sel) 0: mux_22847 = 8'h0; 1: mux_22847 = vout_peek_20537;
    endcase
  endfunction
  wire [7:0] v_22848;
  function [7:0] mux_22848(input [0:0] sel);
    case (sel) 0: mux_22848 = 8'h0; 1: mux_22848 = vout_peek_20528;
    endcase
  endfunction
  wire [7:0] v_22849;
  function [7:0] mux_22849(input [0:0] sel);
    case (sel) 0: mux_22849 = 8'h0; 1: mux_22849 = v_22850;
    endcase
  endfunction
  reg [7:0] v_22850 = 8'h0;
  wire [7:0] v_22851;
  wire [7:0] v_22852;
  function [7:0] mux_22852(input [0:0] sel);
    case (sel) 0: mux_22852 = 8'h0; 1: mux_22852 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22853;
  wire [7:0] v_22854;
  wire [7:0] v_22855;
  function [7:0] mux_22855(input [0:0] sel);
    case (sel) 0: mux_22855 = 8'h0; 1: mux_22855 = v_22856;
    endcase
  endfunction
  reg [7:0] v_22856 = 8'h0;
  wire [7:0] v_22857;
  wire [7:0] v_22858;
  function [7:0] mux_22858(input [0:0] sel);
    case (sel) 0: mux_22858 = 8'h0; 1: mux_22858 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22859;
  wire [7:0] v_22860;
  wire [7:0] v_22861;
  function [7:0] mux_22861(input [0:0] sel);
    case (sel) 0: mux_22861 = 8'h0; 1: mux_22861 = v_22862;
    endcase
  endfunction
  reg [7:0] v_22862 = 8'h0;
  wire [7:0] v_22863;
  wire [7:0] v_22864;
  function [7:0] mux_22864(input [0:0] sel);
    case (sel) 0: mux_22864 = 8'h0; 1: mux_22864 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22865;
  wire [7:0] v_22866;
  wire [7:0] v_22867;
  function [7:0] mux_22867(input [0:0] sel);
    case (sel) 0: mux_22867 = 8'h0; 1: mux_22867 = v_22868;
    endcase
  endfunction
  reg [7:0] v_22868 = 8'h0;
  wire [7:0] v_22869;
  wire [7:0] v_22870;
  function [7:0] mux_22870(input [0:0] sel);
    case (sel) 0: mux_22870 = 8'h0; 1: mux_22870 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22871;
  wire [7:0] v_22872;
  wire [7:0] v_22873;
  function [7:0] mux_22873(input [0:0] sel);
    case (sel) 0: mux_22873 = 8'h0; 1: mux_22873 = v_22874;
    endcase
  endfunction
  reg [7:0] v_22874 = 8'h0;
  wire [7:0] v_22875;
  wire [7:0] v_22876;
  function [7:0] mux_22876(input [0:0] sel);
    case (sel) 0: mux_22876 = 8'h0; 1: mux_22876 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22877;
  wire [7:0] v_22878;
  wire [7:0] v_22879;
  function [7:0] mux_22879(input [0:0] sel);
    case (sel) 0: mux_22879 = 8'h0; 1: mux_22879 = v_22880;
    endcase
  endfunction
  reg [7:0] v_22880 = 8'h0;
  wire [7:0] v_22881;
  wire [7:0] v_22882;
  function [7:0] mux_22882(input [0:0] sel);
    case (sel) 0: mux_22882 = 8'h0; 1: mux_22882 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22883;
  wire [7:0] v_22884;
  wire [7:0] v_22885;
  function [7:0] mux_22885(input [0:0] sel);
    case (sel) 0: mux_22885 = 8'h0; 1: mux_22885 = vout_peek_20405;
    endcase
  endfunction
  wire [7:0] v_22886;
  function [7:0] mux_22886(input [0:0] sel);
    case (sel) 0: mux_22886 = 8'h0; 1: mux_22886 = vout_peek_20396;
    endcase
  endfunction
  wire [7:0] v_22887;
  function [7:0] mux_22887(input [0:0] sel);
    case (sel) 0: mux_22887 = 8'h0; 1: mux_22887 = v_22888;
    endcase
  endfunction
  reg [7:0] v_22888 = 8'h0;
  wire [7:0] v_22889;
  wire [7:0] v_22890;
  function [7:0] mux_22890(input [0:0] sel);
    case (sel) 0: mux_22890 = 8'h0; 1: mux_22890 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22891;
  wire [7:0] v_22892;
  wire [7:0] v_22893;
  function [7:0] mux_22893(input [0:0] sel);
    case (sel) 0: mux_22893 = 8'h0; 1: mux_22893 = vout_peek_20368;
    endcase
  endfunction
  wire [7:0] v_22894;
  function [7:0] mux_22894(input [0:0] sel);
    case (sel) 0: mux_22894 = 8'h0; 1: mux_22894 = vout_peek_20359;
    endcase
  endfunction
  wire [7:0] v_22895;
  function [7:0] mux_22895(input [0:0] sel);
    case (sel) 0: mux_22895 = 8'h0; 1: mux_22895 = v_22896;
    endcase
  endfunction
  reg [7:0] v_22896 = 8'h0;
  wire [7:0] v_22897;
  wire [7:0] v_22898;
  function [7:0] mux_22898(input [0:0] sel);
    case (sel) 0: mux_22898 = 8'h0; 1: mux_22898 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22899;
  wire [7:0] v_22900;
  wire [7:0] v_22901;
  function [7:0] mux_22901(input [0:0] sel);
    case (sel) 0: mux_22901 = 8'h0; 1: mux_22901 = v_22902;
    endcase
  endfunction
  reg [7:0] v_22902 = 8'h0;
  wire [7:0] v_22903;
  wire [7:0] v_22904;
  function [7:0] mux_22904(input [0:0] sel);
    case (sel) 0: mux_22904 = 8'h0; 1: mux_22904 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22905;
  wire [7:0] v_22906;
  wire [7:0] v_22907;
  function [7:0] mux_22907(input [0:0] sel);
    case (sel) 0: mux_22907 = 8'h0; 1: mux_22907 = vout_peek_20312;
    endcase
  endfunction
  wire [7:0] v_22908;
  function [7:0] mux_22908(input [0:0] sel);
    case (sel) 0: mux_22908 = 8'h0; 1: mux_22908 = vout_peek_20303;
    endcase
  endfunction
  wire [7:0] v_22909;
  function [7:0] mux_22909(input [0:0] sel);
    case (sel) 0: mux_22909 = 8'h0; 1: mux_22909 = v_22910;
    endcase
  endfunction
  reg [7:0] v_22910 = 8'h0;
  wire [7:0] v_22911;
  wire [7:0] v_22912;
  function [7:0] mux_22912(input [0:0] sel);
    case (sel) 0: mux_22912 = 8'h0; 1: mux_22912 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22913;
  wire [7:0] v_22914;
  wire [7:0] v_22915;
  function [7:0] mux_22915(input [0:0] sel);
    case (sel) 0: mux_22915 = 8'h0; 1: mux_22915 = vout_peek_20275;
    endcase
  endfunction
  wire [7:0] v_22916;
  function [7:0] mux_22916(input [0:0] sel);
    case (sel) 0: mux_22916 = 8'h0; 1: mux_22916 = vout_peek_20266;
    endcase
  endfunction
  wire [7:0] v_22917;
  function [7:0] mux_22917(input [0:0] sel);
    case (sel) 0: mux_22917 = 8'h0; 1: mux_22917 = v_22918;
    endcase
  endfunction
  reg [7:0] v_22918 = 8'h0;
  wire [7:0] v_22919;
  wire [7:0] v_22920;
  function [7:0] mux_22920(input [0:0] sel);
    case (sel) 0: mux_22920 = 8'h0; 1: mux_22920 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22921;
  wire [7:0] v_22922;
  wire [7:0] v_22923;
  function [7:0] mux_22923(input [0:0] sel);
    case (sel) 0: mux_22923 = 8'h0; 1: mux_22923 = v_22924;
    endcase
  endfunction
  reg [7:0] v_22924 = 8'h0;
  wire [7:0] v_22925;
  wire [7:0] v_22926;
  function [7:0] mux_22926(input [0:0] sel);
    case (sel) 0: mux_22926 = 8'h0; 1: mux_22926 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22927;
  wire [7:0] v_22928;
  wire [7:0] v_22929;
  function [7:0] mux_22929(input [0:0] sel);
    case (sel) 0: mux_22929 = 8'h0; 1: mux_22929 = v_22930;
    endcase
  endfunction
  reg [7:0] v_22930 = 8'h0;
  wire [7:0] v_22931;
  wire [7:0] v_22932;
  function [7:0] mux_22932(input [0:0] sel);
    case (sel) 0: mux_22932 = 8'h0; 1: mux_22932 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22933;
  wire [7:0] v_22934;
  wire [7:0] v_22935;
  function [7:0] mux_22935(input [0:0] sel);
    case (sel) 0: mux_22935 = 8'h0; 1: mux_22935 = vout_peek_20200;
    endcase
  endfunction
  wire [7:0] v_22936;
  function [7:0] mux_22936(input [0:0] sel);
    case (sel) 0: mux_22936 = 8'h0; 1: mux_22936 = vout_peek_20191;
    endcase
  endfunction
  wire [7:0] v_22937;
  function [7:0] mux_22937(input [0:0] sel);
    case (sel) 0: mux_22937 = 8'h0; 1: mux_22937 = v_22938;
    endcase
  endfunction
  reg [7:0] v_22938 = 8'h0;
  wire [7:0] v_22939;
  wire [7:0] v_22940;
  function [7:0] mux_22940(input [0:0] sel);
    case (sel) 0: mux_22940 = 8'h0; 1: mux_22940 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22941;
  wire [7:0] v_22942;
  wire [7:0] v_22943;
  function [7:0] mux_22943(input [0:0] sel);
    case (sel) 0: mux_22943 = 8'h0; 1: mux_22943 = vout_peek_20163;
    endcase
  endfunction
  wire [7:0] v_22944;
  function [7:0] mux_22944(input [0:0] sel);
    case (sel) 0: mux_22944 = 8'h0; 1: mux_22944 = vout_peek_20154;
    endcase
  endfunction
  wire [7:0] v_22945;
  function [7:0] mux_22945(input [0:0] sel);
    case (sel) 0: mux_22945 = 8'h0; 1: mux_22945 = v_22946;
    endcase
  endfunction
  reg [7:0] v_22946 = 8'h0;
  wire [7:0] v_22947;
  wire [7:0] v_22948;
  function [7:0] mux_22948(input [0:0] sel);
    case (sel) 0: mux_22948 = 8'h0; 1: mux_22948 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22949;
  wire [7:0] v_22950;
  wire [7:0] v_22951;
  function [7:0] mux_22951(input [0:0] sel);
    case (sel) 0: mux_22951 = 8'h0; 1: mux_22951 = v_22952;
    endcase
  endfunction
  reg [7:0] v_22952 = 8'h0;
  wire [7:0] v_22953;
  wire [7:0] v_22954;
  function [7:0] mux_22954(input [0:0] sel);
    case (sel) 0: mux_22954 = 8'h0; 1: mux_22954 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22955;
  wire [7:0] v_22956;
  wire [7:0] v_22957;
  function [7:0] mux_22957(input [0:0] sel);
    case (sel) 0: mux_22957 = 8'h0; 1: mux_22957 = vout_peek_20107;
    endcase
  endfunction
  wire [7:0] v_22958;
  function [7:0] mux_22958(input [0:0] sel);
    case (sel) 0: mux_22958 = 8'h0; 1: mux_22958 = vout_peek_20098;
    endcase
  endfunction
  wire [7:0] v_22959;
  function [7:0] mux_22959(input [0:0] sel);
    case (sel) 0: mux_22959 = 8'h0; 1: mux_22959 = v_22960;
    endcase
  endfunction
  reg [7:0] v_22960 = 8'h0;
  wire [7:0] v_22961;
  wire [7:0] v_22962;
  function [7:0] mux_22962(input [0:0] sel);
    case (sel) 0: mux_22962 = 8'h0; 1: mux_22962 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22963;
  wire [7:0] v_22964;
  wire [7:0] v_22965;
  function [7:0] mux_22965(input [0:0] sel);
    case (sel) 0: mux_22965 = 8'h0; 1: mux_22965 = vout_peek_20070;
    endcase
  endfunction
  wire [7:0] v_22966;
  function [7:0] mux_22966(input [0:0] sel);
    case (sel) 0: mux_22966 = 8'h0; 1: mux_22966 = vout_peek_20061;
    endcase
  endfunction
  wire [7:0] v_22967;
  function [7:0] mux_22967(input [0:0] sel);
    case (sel) 0: mux_22967 = 8'h0; 1: mux_22967 = v_22968;
    endcase
  endfunction
  reg [7:0] v_22968 = 8'h0;
  wire [7:0] v_22969;
  wire [7:0] v_22970;
  function [7:0] mux_22970(input [0:0] sel);
    case (sel) 0: mux_22970 = 8'h0; 1: mux_22970 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22971;
  wire [7:0] v_22972;
  wire [7:0] v_22973;
  function [7:0] mux_22973(input [0:0] sel);
    case (sel) 0: mux_22973 = 8'h0; 1: mux_22973 = v_22974;
    endcase
  endfunction
  reg [7:0] v_22974 = 8'h0;
  wire [7:0] v_22975;
  wire [7:0] v_22976;
  function [7:0] mux_22976(input [0:0] sel);
    case (sel) 0: mux_22976 = 8'h0; 1: mux_22976 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22977;
  wire [7:0] v_22978;
  wire [7:0] v_22979;
  function [7:0] mux_22979(input [0:0] sel);
    case (sel) 0: mux_22979 = 8'h0; 1: mux_22979 = v_22980;
    endcase
  endfunction
  reg [7:0] v_22980 = 8'h0;
  wire [7:0] v_22981;
  wire [7:0] v_22982;
  function [7:0] mux_22982(input [0:0] sel);
    case (sel) 0: mux_22982 = 8'h0; 1: mux_22982 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22983;
  wire [7:0] v_22984;
  wire [7:0] v_22985;
  function [7:0] mux_22985(input [0:0] sel);
    case (sel) 0: mux_22985 = 8'h0; 1: mux_22985 = v_22986;
    endcase
  endfunction
  reg [7:0] v_22986 = 8'h0;
  wire [7:0] v_22987;
  wire [7:0] v_22988;
  function [7:0] mux_22988(input [0:0] sel);
    case (sel) 0: mux_22988 = 8'h0; 1: mux_22988 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22989;
  wire [7:0] v_22990;
  wire [7:0] v_22991;
  function [7:0] mux_22991(input [0:0] sel);
    case (sel) 0: mux_22991 = 8'h0; 1: mux_22991 = vout_peek_19976;
    endcase
  endfunction
  wire [7:0] v_22992;
  function [7:0] mux_22992(input [0:0] sel);
    case (sel) 0: mux_22992 = 8'h0; 1: mux_22992 = vout_peek_19967;
    endcase
  endfunction
  wire [7:0] v_22993;
  function [7:0] mux_22993(input [0:0] sel);
    case (sel) 0: mux_22993 = 8'h0; 1: mux_22993 = v_22994;
    endcase
  endfunction
  reg [7:0] v_22994 = 8'h0;
  wire [7:0] v_22995;
  wire [7:0] v_22996;
  function [7:0] mux_22996(input [0:0] sel);
    case (sel) 0: mux_22996 = 8'h0; 1: mux_22996 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_22997;
  wire [7:0] v_22998;
  wire [7:0] v_22999;
  function [7:0] mux_22999(input [0:0] sel);
    case (sel) 0: mux_22999 = 8'h0; 1: mux_22999 = vout_peek_19939;
    endcase
  endfunction
  wire [7:0] v_23000;
  function [7:0] mux_23000(input [0:0] sel);
    case (sel) 0: mux_23000 = 8'h0; 1: mux_23000 = vout_peek_19930;
    endcase
  endfunction
  wire [7:0] v_23001;
  function [7:0] mux_23001(input [0:0] sel);
    case (sel) 0: mux_23001 = 8'h0; 1: mux_23001 = v_23002;
    endcase
  endfunction
  reg [7:0] v_23002 = 8'h0;
  wire [7:0] v_23003;
  wire [7:0] v_23004;
  function [7:0] mux_23004(input [0:0] sel);
    case (sel) 0: mux_23004 = 8'h0; 1: mux_23004 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23005;
  wire [7:0] v_23006;
  wire [7:0] v_23007;
  function [7:0] mux_23007(input [0:0] sel);
    case (sel) 0: mux_23007 = 8'h0; 1: mux_23007 = v_23008;
    endcase
  endfunction
  reg [7:0] v_23008 = 8'h0;
  wire [7:0] v_23009;
  wire [7:0] v_23010;
  function [7:0] mux_23010(input [0:0] sel);
    case (sel) 0: mux_23010 = 8'h0; 1: mux_23010 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23011;
  wire [7:0] v_23012;
  wire [7:0] v_23013;
  function [7:0] mux_23013(input [0:0] sel);
    case (sel) 0: mux_23013 = 8'h0; 1: mux_23013 = vout_peek_19883;
    endcase
  endfunction
  wire [7:0] v_23014;
  function [7:0] mux_23014(input [0:0] sel);
    case (sel) 0: mux_23014 = 8'h0; 1: mux_23014 = vout_peek_19874;
    endcase
  endfunction
  wire [7:0] v_23015;
  function [7:0] mux_23015(input [0:0] sel);
    case (sel) 0: mux_23015 = 8'h0; 1: mux_23015 = v_23016;
    endcase
  endfunction
  reg [7:0] v_23016 = 8'h0;
  wire [7:0] v_23017;
  wire [7:0] v_23018;
  function [7:0] mux_23018(input [0:0] sel);
    case (sel) 0: mux_23018 = 8'h0; 1: mux_23018 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23019;
  wire [7:0] v_23020;
  wire [7:0] v_23021;
  function [7:0] mux_23021(input [0:0] sel);
    case (sel) 0: mux_23021 = 8'h0; 1: mux_23021 = vout_peek_19846;
    endcase
  endfunction
  wire [7:0] v_23022;
  function [7:0] mux_23022(input [0:0] sel);
    case (sel) 0: mux_23022 = 8'h0; 1: mux_23022 = vout_peek_19837;
    endcase
  endfunction
  wire [7:0] v_23023;
  function [7:0] mux_23023(input [0:0] sel);
    case (sel) 0: mux_23023 = 8'h0; 1: mux_23023 = v_23024;
    endcase
  endfunction
  reg [7:0] v_23024 = 8'h0;
  wire [7:0] v_23025;
  wire [7:0] v_23026;
  function [7:0] mux_23026(input [0:0] sel);
    case (sel) 0: mux_23026 = 8'h0; 1: mux_23026 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23027;
  wire [7:0] v_23028;
  wire [7:0] v_23029;
  function [7:0] mux_23029(input [0:0] sel);
    case (sel) 0: mux_23029 = 8'h0; 1: mux_23029 = v_23030;
    endcase
  endfunction
  reg [7:0] v_23030 = 8'h0;
  wire [7:0] v_23031;
  wire [7:0] v_23032;
  function [7:0] mux_23032(input [0:0] sel);
    case (sel) 0: mux_23032 = 8'h0; 1: mux_23032 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23033;
  wire [7:0] v_23034;
  wire [7:0] v_23035;
  function [7:0] mux_23035(input [0:0] sel);
    case (sel) 0: mux_23035 = 8'h0; 1: mux_23035 = v_23036;
    endcase
  endfunction
  reg [7:0] v_23036 = 8'h0;
  wire [7:0] v_23037;
  wire [7:0] v_23038;
  function [7:0] mux_23038(input [0:0] sel);
    case (sel) 0: mux_23038 = 8'h0; 1: mux_23038 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23039;
  wire [7:0] v_23040;
  wire [7:0] v_23041;
  function [7:0] mux_23041(input [0:0] sel);
    case (sel) 0: mux_23041 = 8'h0; 1: mux_23041 = vout_peek_19771;
    endcase
  endfunction
  wire [7:0] v_23042;
  function [7:0] mux_23042(input [0:0] sel);
    case (sel) 0: mux_23042 = 8'h0; 1: mux_23042 = vout_peek_19762;
    endcase
  endfunction
  wire [7:0] v_23043;
  function [7:0] mux_23043(input [0:0] sel);
    case (sel) 0: mux_23043 = 8'h0; 1: mux_23043 = v_23044;
    endcase
  endfunction
  reg [7:0] v_23044 = 8'h0;
  wire [7:0] v_23045;
  wire [7:0] v_23046;
  function [7:0] mux_23046(input [0:0] sel);
    case (sel) 0: mux_23046 = 8'h0; 1: mux_23046 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23047;
  wire [7:0] v_23048;
  wire [7:0] v_23049;
  function [7:0] mux_23049(input [0:0] sel);
    case (sel) 0: mux_23049 = 8'h0; 1: mux_23049 = vout_peek_19734;
    endcase
  endfunction
  wire [7:0] v_23050;
  function [7:0] mux_23050(input [0:0] sel);
    case (sel) 0: mux_23050 = 8'h0; 1: mux_23050 = vout_peek_19725;
    endcase
  endfunction
  wire [7:0] v_23051;
  function [7:0] mux_23051(input [0:0] sel);
    case (sel) 0: mux_23051 = 8'h0; 1: mux_23051 = v_23052;
    endcase
  endfunction
  reg [7:0] v_23052 = 8'h0;
  wire [7:0] v_23053;
  wire [7:0] v_23054;
  function [7:0] mux_23054(input [0:0] sel);
    case (sel) 0: mux_23054 = 8'h0; 1: mux_23054 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23055;
  wire [7:0] v_23056;
  wire [7:0] v_23057;
  function [7:0] mux_23057(input [0:0] sel);
    case (sel) 0: mux_23057 = 8'h0; 1: mux_23057 = v_23058;
    endcase
  endfunction
  reg [7:0] v_23058 = 8'h0;
  wire [7:0] v_23059;
  wire [7:0] v_23060;
  function [7:0] mux_23060(input [0:0] sel);
    case (sel) 0: mux_23060 = 8'h0; 1: mux_23060 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23061;
  wire [7:0] v_23062;
  wire [7:0] v_23063;
  function [7:0] mux_23063(input [0:0] sel);
    case (sel) 0: mux_23063 = 8'h0; 1: mux_23063 = vout_peek_19678;
    endcase
  endfunction
  wire [7:0] v_23064;
  function [7:0] mux_23064(input [0:0] sel);
    case (sel) 0: mux_23064 = 8'h0; 1: mux_23064 = vout_peek_19669;
    endcase
  endfunction
  wire [7:0] v_23065;
  function [7:0] mux_23065(input [0:0] sel);
    case (sel) 0: mux_23065 = 8'h0; 1: mux_23065 = v_23066;
    endcase
  endfunction
  reg [7:0] v_23066 = 8'h0;
  wire [7:0] v_23067;
  wire [7:0] v_23068;
  function [7:0] mux_23068(input [0:0] sel);
    case (sel) 0: mux_23068 = 8'h0; 1: mux_23068 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23069;
  wire [7:0] v_23070;
  wire [7:0] v_23071;
  function [7:0] mux_23071(input [0:0] sel);
    case (sel) 0: mux_23071 = 8'h0; 1: mux_23071 = vout_peek_19641;
    endcase
  endfunction
  wire [7:0] v_23072;
  function [7:0] mux_23072(input [0:0] sel);
    case (sel) 0: mux_23072 = 8'h0; 1: mux_23072 = vout_peek_19632;
    endcase
  endfunction
  wire [7:0] v_23073;
  function [7:0] mux_23073(input [0:0] sel);
    case (sel) 0: mux_23073 = 8'h0; 1: mux_23073 = v_23074;
    endcase
  endfunction
  reg [7:0] v_23074 = 8'h0;
  wire [7:0] v_23075;
  wire [7:0] v_23076;
  function [7:0] mux_23076(input [0:0] sel);
    case (sel) 0: mux_23076 = 8'h0; 1: mux_23076 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23077;
  wire [7:0] v_23078;
  wire [7:0] v_23079;
  function [7:0] mux_23079(input [0:0] sel);
    case (sel) 0: mux_23079 = 8'h0; 1: mux_23079 = v_23080;
    endcase
  endfunction
  reg [7:0] v_23080 = 8'h0;
  wire [7:0] v_23081;
  wire [7:0] v_23082;
  function [7:0] mux_23082(input [0:0] sel);
    case (sel) 0: mux_23082 = 8'h0; 1: mux_23082 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23083;
  wire [7:0] v_23084;
  wire [7:0] v_23085;
  function [7:0] mux_23085(input [0:0] sel);
    case (sel) 0: mux_23085 = 8'h0; 1: mux_23085 = v_23086;
    endcase
  endfunction
  reg [7:0] v_23086 = 8'h0;
  wire [7:0] v_23087;
  wire [7:0] v_23088;
  function [7:0] mux_23088(input [0:0] sel);
    case (sel) 0: mux_23088 = 8'h0; 1: mux_23088 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23089;
  wire [7:0] v_23090;
  wire [7:0] v_23091;
  function [7:0] mux_23091(input [0:0] sel);
    case (sel) 0: mux_23091 = 8'h0; 1: mux_23091 = v_23092;
    endcase
  endfunction
  reg [7:0] v_23092 = 8'h0;
  wire [7:0] v_23093;
  wire [7:0] v_23094;
  function [7:0] mux_23094(input [0:0] sel);
    case (sel) 0: mux_23094 = 8'h0; 1: mux_23094 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23095;
  wire [7:0] v_23096;
  wire [7:0] v_23097;
  function [7:0] mux_23097(input [0:0] sel);
    case (sel) 0: mux_23097 = 8'h0; 1: mux_23097 = v_23098;
    endcase
  endfunction
  reg [7:0] v_23098 = 8'h0;
  wire [7:0] v_23099;
  wire [7:0] v_23100;
  function [7:0] mux_23100(input [0:0] sel);
    case (sel) 0: mux_23100 = 8'h0; 1: mux_23100 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23101;
  wire [7:0] v_23102;
  wire [7:0] v_23103;
  function [7:0] mux_23103(input [0:0] sel);
    case (sel) 0: mux_23103 = 8'h0; 1: mux_23103 = vout_peek_19528;
    endcase
  endfunction
  wire [7:0] v_23104;
  function [7:0] mux_23104(input [0:0] sel);
    case (sel) 0: mux_23104 = 8'h0; 1: mux_23104 = vout_peek_19519;
    endcase
  endfunction
  wire [7:0] v_23105;
  function [7:0] mux_23105(input [0:0] sel);
    case (sel) 0: mux_23105 = 8'h0; 1: mux_23105 = v_23106;
    endcase
  endfunction
  reg [7:0] v_23106 = 8'h0;
  wire [7:0] v_23107;
  wire [7:0] v_23108;
  function [7:0] mux_23108(input [0:0] sel);
    case (sel) 0: mux_23108 = 8'h0; 1: mux_23108 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23109;
  wire [7:0] v_23110;
  wire [7:0] v_23111;
  function [7:0] mux_23111(input [0:0] sel);
    case (sel) 0: mux_23111 = 8'h0; 1: mux_23111 = vout_peek_19491;
    endcase
  endfunction
  wire [7:0] v_23112;
  function [7:0] mux_23112(input [0:0] sel);
    case (sel) 0: mux_23112 = 8'h0; 1: mux_23112 = vout_peek_19482;
    endcase
  endfunction
  wire [7:0] v_23113;
  function [7:0] mux_23113(input [0:0] sel);
    case (sel) 0: mux_23113 = 8'h0; 1: mux_23113 = v_23114;
    endcase
  endfunction
  reg [7:0] v_23114 = 8'h0;
  wire [7:0] v_23115;
  wire [7:0] v_23116;
  function [7:0] mux_23116(input [0:0] sel);
    case (sel) 0: mux_23116 = 8'h0; 1: mux_23116 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23117;
  wire [7:0] v_23118;
  wire [7:0] v_23119;
  function [7:0] mux_23119(input [0:0] sel);
    case (sel) 0: mux_23119 = 8'h0; 1: mux_23119 = v_23120;
    endcase
  endfunction
  reg [7:0] v_23120 = 8'h0;
  wire [7:0] v_23121;
  wire [7:0] v_23122;
  function [7:0] mux_23122(input [0:0] sel);
    case (sel) 0: mux_23122 = 8'h0; 1: mux_23122 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23123;
  wire [7:0] v_23124;
  wire [7:0] v_23125;
  function [7:0] mux_23125(input [0:0] sel);
    case (sel) 0: mux_23125 = 8'h0; 1: mux_23125 = vout_peek_19435;
    endcase
  endfunction
  wire [7:0] v_23126;
  function [7:0] mux_23126(input [0:0] sel);
    case (sel) 0: mux_23126 = 8'h0; 1: mux_23126 = vout_peek_19426;
    endcase
  endfunction
  wire [7:0] v_23127;
  function [7:0] mux_23127(input [0:0] sel);
    case (sel) 0: mux_23127 = 8'h0; 1: mux_23127 = v_23128;
    endcase
  endfunction
  reg [7:0] v_23128 = 8'h0;
  wire [7:0] v_23129;
  wire [7:0] v_23130;
  function [7:0] mux_23130(input [0:0] sel);
    case (sel) 0: mux_23130 = 8'h0; 1: mux_23130 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23131;
  wire [7:0] v_23132;
  wire [7:0] v_23133;
  function [7:0] mux_23133(input [0:0] sel);
    case (sel) 0: mux_23133 = 8'h0; 1: mux_23133 = vout_peek_19398;
    endcase
  endfunction
  wire [7:0] v_23134;
  function [7:0] mux_23134(input [0:0] sel);
    case (sel) 0: mux_23134 = 8'h0; 1: mux_23134 = vout_peek_19389;
    endcase
  endfunction
  wire [7:0] v_23135;
  function [7:0] mux_23135(input [0:0] sel);
    case (sel) 0: mux_23135 = 8'h0; 1: mux_23135 = v_23136;
    endcase
  endfunction
  reg [7:0] v_23136 = 8'h0;
  wire [7:0] v_23137;
  wire [7:0] v_23138;
  function [7:0] mux_23138(input [0:0] sel);
    case (sel) 0: mux_23138 = 8'h0; 1: mux_23138 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23139;
  wire [7:0] v_23140;
  wire [7:0] v_23141;
  function [7:0] mux_23141(input [0:0] sel);
    case (sel) 0: mux_23141 = 8'h0; 1: mux_23141 = v_23142;
    endcase
  endfunction
  reg [7:0] v_23142 = 8'h0;
  wire [7:0] v_23143;
  wire [7:0] v_23144;
  function [7:0] mux_23144(input [0:0] sel);
    case (sel) 0: mux_23144 = 8'h0; 1: mux_23144 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23145;
  wire [7:0] v_23146;
  wire [7:0] v_23147;
  function [7:0] mux_23147(input [0:0] sel);
    case (sel) 0: mux_23147 = 8'h0; 1: mux_23147 = v_23148;
    endcase
  endfunction
  reg [7:0] v_23148 = 8'h0;
  wire [7:0] v_23149;
  wire [7:0] v_23150;
  function [7:0] mux_23150(input [0:0] sel);
    case (sel) 0: mux_23150 = 8'h0; 1: mux_23150 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23151;
  wire [7:0] v_23152;
  wire [7:0] v_23153;
  function [7:0] mux_23153(input [0:0] sel);
    case (sel) 0: mux_23153 = 8'h0; 1: mux_23153 = vout_peek_19323;
    endcase
  endfunction
  wire [7:0] v_23154;
  function [7:0] mux_23154(input [0:0] sel);
    case (sel) 0: mux_23154 = 8'h0; 1: mux_23154 = vout_peek_19314;
    endcase
  endfunction
  wire [7:0] v_23155;
  function [7:0] mux_23155(input [0:0] sel);
    case (sel) 0: mux_23155 = 8'h0; 1: mux_23155 = v_23156;
    endcase
  endfunction
  reg [7:0] v_23156 = 8'h0;
  wire [7:0] v_23157;
  wire [7:0] v_23158;
  function [7:0] mux_23158(input [0:0] sel);
    case (sel) 0: mux_23158 = 8'h0; 1: mux_23158 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23159;
  wire [7:0] v_23160;
  wire [7:0] v_23161;
  function [7:0] mux_23161(input [0:0] sel);
    case (sel) 0: mux_23161 = 8'h0; 1: mux_23161 = vout_peek_19286;
    endcase
  endfunction
  wire [7:0] v_23162;
  function [7:0] mux_23162(input [0:0] sel);
    case (sel) 0: mux_23162 = 8'h0; 1: mux_23162 = vout_peek_19277;
    endcase
  endfunction
  wire [7:0] v_23163;
  function [7:0] mux_23163(input [0:0] sel);
    case (sel) 0: mux_23163 = 8'h0; 1: mux_23163 = v_23164;
    endcase
  endfunction
  reg [7:0] v_23164 = 8'h0;
  wire [7:0] v_23165;
  wire [7:0] v_23166;
  function [7:0] mux_23166(input [0:0] sel);
    case (sel) 0: mux_23166 = 8'h0; 1: mux_23166 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23167;
  wire [7:0] v_23168;
  wire [7:0] v_23169;
  function [7:0] mux_23169(input [0:0] sel);
    case (sel) 0: mux_23169 = 8'h0; 1: mux_23169 = v_23170;
    endcase
  endfunction
  reg [7:0] v_23170 = 8'h0;
  wire [7:0] v_23171;
  wire [7:0] v_23172;
  function [7:0] mux_23172(input [0:0] sel);
    case (sel) 0: mux_23172 = 8'h0; 1: mux_23172 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23173;
  wire [7:0] v_23174;
  wire [7:0] v_23175;
  function [7:0] mux_23175(input [0:0] sel);
    case (sel) 0: mux_23175 = 8'h0; 1: mux_23175 = vout_peek_19230;
    endcase
  endfunction
  wire [7:0] v_23176;
  function [7:0] mux_23176(input [0:0] sel);
    case (sel) 0: mux_23176 = 8'h0; 1: mux_23176 = vout_peek_19221;
    endcase
  endfunction
  wire [7:0] v_23177;
  function [7:0] mux_23177(input [0:0] sel);
    case (sel) 0: mux_23177 = 8'h0; 1: mux_23177 = v_23178;
    endcase
  endfunction
  reg [7:0] v_23178 = 8'h0;
  wire [7:0] v_23179;
  wire [7:0] v_23180;
  function [7:0] mux_23180(input [0:0] sel);
    case (sel) 0: mux_23180 = 8'h0; 1: mux_23180 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23181;
  wire [7:0] v_23182;
  wire [7:0] v_23183;
  function [7:0] mux_23183(input [0:0] sel);
    case (sel) 0: mux_23183 = 8'h0; 1: mux_23183 = vout_peek_19193;
    endcase
  endfunction
  wire [7:0] v_23184;
  function [7:0] mux_23184(input [0:0] sel);
    case (sel) 0: mux_23184 = 8'h0; 1: mux_23184 = vout_peek_19184;
    endcase
  endfunction
  wire [7:0] v_23185;
  function [7:0] mux_23185(input [0:0] sel);
    case (sel) 0: mux_23185 = 8'h0; 1: mux_23185 = v_23186;
    endcase
  endfunction
  reg [7:0] v_23186 = 8'h0;
  wire [7:0] v_23187;
  wire [7:0] v_23188;
  function [7:0] mux_23188(input [0:0] sel);
    case (sel) 0: mux_23188 = 8'h0; 1: mux_23188 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23189;
  wire [7:0] v_23190;
  wire [7:0] v_23191;
  function [7:0] mux_23191(input [0:0] sel);
    case (sel) 0: mux_23191 = 8'h0; 1: mux_23191 = v_23192;
    endcase
  endfunction
  reg [7:0] v_23192 = 8'h0;
  wire [7:0] v_23193;
  wire [7:0] v_23194;
  function [7:0] mux_23194(input [0:0] sel);
    case (sel) 0: mux_23194 = 8'h0; 1: mux_23194 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23195;
  wire [7:0] v_23196;
  wire [7:0] v_23197;
  function [7:0] mux_23197(input [0:0] sel);
    case (sel) 0: mux_23197 = 8'h0; 1: mux_23197 = v_23198;
    endcase
  endfunction
  reg [7:0] v_23198 = 8'h0;
  wire [7:0] v_23199;
  wire [7:0] v_23200;
  function [7:0] mux_23200(input [0:0] sel);
    case (sel) 0: mux_23200 = 8'h0; 1: mux_23200 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23201;
  wire [7:0] v_23202;
  wire [7:0] v_23203;
  function [7:0] mux_23203(input [0:0] sel);
    case (sel) 0: mux_23203 = 8'h0; 1: mux_23203 = v_23204;
    endcase
  endfunction
  reg [7:0] v_23204 = 8'h0;
  wire [7:0] v_23205;
  wire [7:0] v_23206;
  function [7:0] mux_23206(input [0:0] sel);
    case (sel) 0: mux_23206 = 8'h0; 1: mux_23206 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23207;
  wire [7:0] v_23208;
  wire [7:0] v_23209;
  function [7:0] mux_23209(input [0:0] sel);
    case (sel) 0: mux_23209 = 8'h0; 1: mux_23209 = vout_peek_19099;
    endcase
  endfunction
  wire [7:0] v_23210;
  function [7:0] mux_23210(input [0:0] sel);
    case (sel) 0: mux_23210 = 8'h0; 1: mux_23210 = vout_peek_19090;
    endcase
  endfunction
  wire [7:0] v_23211;
  function [7:0] mux_23211(input [0:0] sel);
    case (sel) 0: mux_23211 = 8'h0; 1: mux_23211 = v_23212;
    endcase
  endfunction
  reg [7:0] v_23212 = 8'h0;
  wire [7:0] v_23213;
  wire [7:0] v_23214;
  function [7:0] mux_23214(input [0:0] sel);
    case (sel) 0: mux_23214 = 8'h0; 1: mux_23214 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23215;
  wire [7:0] v_23216;
  wire [7:0] v_23217;
  function [7:0] mux_23217(input [0:0] sel);
    case (sel) 0: mux_23217 = 8'h0; 1: mux_23217 = vout_peek_19062;
    endcase
  endfunction
  wire [7:0] v_23218;
  function [7:0] mux_23218(input [0:0] sel);
    case (sel) 0: mux_23218 = 8'h0; 1: mux_23218 = vout_peek_19053;
    endcase
  endfunction
  wire [7:0] v_23219;
  function [7:0] mux_23219(input [0:0] sel);
    case (sel) 0: mux_23219 = 8'h0; 1: mux_23219 = v_23220;
    endcase
  endfunction
  reg [7:0] v_23220 = 8'h0;
  wire [7:0] v_23221;
  wire [7:0] v_23222;
  function [7:0] mux_23222(input [0:0] sel);
    case (sel) 0: mux_23222 = 8'h0; 1: mux_23222 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23223;
  wire [7:0] v_23224;
  wire [7:0] v_23225;
  function [7:0] mux_23225(input [0:0] sel);
    case (sel) 0: mux_23225 = 8'h0; 1: mux_23225 = v_23226;
    endcase
  endfunction
  reg [7:0] v_23226 = 8'h0;
  wire [7:0] v_23227;
  wire [7:0] v_23228;
  function [7:0] mux_23228(input [0:0] sel);
    case (sel) 0: mux_23228 = 8'h0; 1: mux_23228 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23229;
  wire [7:0] v_23230;
  wire [7:0] v_23231;
  function [7:0] mux_23231(input [0:0] sel);
    case (sel) 0: mux_23231 = 8'h0; 1: mux_23231 = vout_peek_19006;
    endcase
  endfunction
  wire [7:0] v_23232;
  function [7:0] mux_23232(input [0:0] sel);
    case (sel) 0: mux_23232 = 8'h0; 1: mux_23232 = vout_peek_18997;
    endcase
  endfunction
  wire [7:0] v_23233;
  function [7:0] mux_23233(input [0:0] sel);
    case (sel) 0: mux_23233 = 8'h0; 1: mux_23233 = v_23234;
    endcase
  endfunction
  reg [7:0] v_23234 = 8'h0;
  wire [7:0] v_23235;
  wire [7:0] v_23236;
  function [7:0] mux_23236(input [0:0] sel);
    case (sel) 0: mux_23236 = 8'h0; 1: mux_23236 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23237;
  wire [7:0] v_23238;
  wire [7:0] v_23239;
  function [7:0] mux_23239(input [0:0] sel);
    case (sel) 0: mux_23239 = 8'h0; 1: mux_23239 = vout_peek_18969;
    endcase
  endfunction
  wire [7:0] v_23240;
  function [7:0] mux_23240(input [0:0] sel);
    case (sel) 0: mux_23240 = 8'h0; 1: mux_23240 = vout_peek_18960;
    endcase
  endfunction
  wire [7:0] v_23241;
  function [7:0] mux_23241(input [0:0] sel);
    case (sel) 0: mux_23241 = 8'h0; 1: mux_23241 = v_23242;
    endcase
  endfunction
  reg [7:0] v_23242 = 8'h0;
  wire [7:0] v_23243;
  wire [7:0] v_23244;
  function [7:0] mux_23244(input [0:0] sel);
    case (sel) 0: mux_23244 = 8'h0; 1: mux_23244 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23245;
  wire [7:0] v_23246;
  wire [7:0] v_23247;
  function [7:0] mux_23247(input [0:0] sel);
    case (sel) 0: mux_23247 = 8'h0; 1: mux_23247 = v_23248;
    endcase
  endfunction
  reg [7:0] v_23248 = 8'h0;
  wire [7:0] v_23249;
  wire [7:0] v_23250;
  function [7:0] mux_23250(input [0:0] sel);
    case (sel) 0: mux_23250 = 8'h0; 1: mux_23250 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23251;
  wire [7:0] v_23252;
  wire [7:0] v_23253;
  function [7:0] mux_23253(input [0:0] sel);
    case (sel) 0: mux_23253 = 8'h0; 1: mux_23253 = v_23254;
    endcase
  endfunction
  reg [7:0] v_23254 = 8'h0;
  wire [7:0] v_23255;
  wire [7:0] v_23256;
  function [7:0] mux_23256(input [0:0] sel);
    case (sel) 0: mux_23256 = 8'h0; 1: mux_23256 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23257;
  wire [7:0] v_23258;
  wire [7:0] v_23259;
  function [7:0] mux_23259(input [0:0] sel);
    case (sel) 0: mux_23259 = 8'h0; 1: mux_23259 = vout_peek_18894;
    endcase
  endfunction
  wire [7:0] v_23260;
  function [7:0] mux_23260(input [0:0] sel);
    case (sel) 0: mux_23260 = 8'h0; 1: mux_23260 = vout_peek_18885;
    endcase
  endfunction
  wire [7:0] v_23261;
  function [7:0] mux_23261(input [0:0] sel);
    case (sel) 0: mux_23261 = 8'h0; 1: mux_23261 = v_23262;
    endcase
  endfunction
  reg [7:0] v_23262 = 8'h0;
  wire [7:0] v_23263;
  wire [7:0] v_23264;
  function [7:0] mux_23264(input [0:0] sel);
    case (sel) 0: mux_23264 = 8'h0; 1: mux_23264 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23265;
  wire [7:0] v_23266;
  wire [7:0] v_23267;
  function [7:0] mux_23267(input [0:0] sel);
    case (sel) 0: mux_23267 = 8'h0; 1: mux_23267 = vout_peek_18857;
    endcase
  endfunction
  wire [7:0] v_23268;
  function [7:0] mux_23268(input [0:0] sel);
    case (sel) 0: mux_23268 = 8'h0; 1: mux_23268 = vout_peek_18848;
    endcase
  endfunction
  wire [7:0] v_23269;
  function [7:0] mux_23269(input [0:0] sel);
    case (sel) 0: mux_23269 = 8'h0; 1: mux_23269 = v_23270;
    endcase
  endfunction
  reg [7:0] v_23270 = 8'h0;
  wire [7:0] v_23271;
  wire [7:0] v_23272;
  function [7:0] mux_23272(input [0:0] sel);
    case (sel) 0: mux_23272 = 8'h0; 1: mux_23272 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23273;
  wire [7:0] v_23274;
  wire [7:0] v_23275;
  function [7:0] mux_23275(input [0:0] sel);
    case (sel) 0: mux_23275 = 8'h0; 1: mux_23275 = v_23276;
    endcase
  endfunction
  reg [7:0] v_23276 = 8'h0;
  wire [7:0] v_23277;
  wire [7:0] v_23278;
  function [7:0] mux_23278(input [0:0] sel);
    case (sel) 0: mux_23278 = 8'h0; 1: mux_23278 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23279;
  wire [7:0] v_23280;
  wire [7:0] v_23281;
  function [7:0] mux_23281(input [0:0] sel);
    case (sel) 0: mux_23281 = 8'h0; 1: mux_23281 = vout_peek_18801;
    endcase
  endfunction
  wire [7:0] v_23282;
  function [7:0] mux_23282(input [0:0] sel);
    case (sel) 0: mux_23282 = 8'h0; 1: mux_23282 = vout_peek_18792;
    endcase
  endfunction
  wire [7:0] v_23283;
  function [7:0] mux_23283(input [0:0] sel);
    case (sel) 0: mux_23283 = 8'h0; 1: mux_23283 = v_23284;
    endcase
  endfunction
  reg [7:0] v_23284 = 8'h0;
  wire [7:0] v_23285;
  wire [7:0] v_23286;
  function [7:0] mux_23286(input [0:0] sel);
    case (sel) 0: mux_23286 = 8'h0; 1: mux_23286 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23287;
  wire [7:0] v_23288;
  wire [7:0] v_23289;
  function [7:0] mux_23289(input [0:0] sel);
    case (sel) 0: mux_23289 = 8'h0; 1: mux_23289 = vout_peek_18764;
    endcase
  endfunction
  wire [7:0] v_23290;
  function [7:0] mux_23290(input [0:0] sel);
    case (sel) 0: mux_23290 = 8'h0; 1: mux_23290 = vout_peek_18755;
    endcase
  endfunction
  wire [7:0] v_23291;
  function [7:0] mux_23291(input [0:0] sel);
    case (sel) 0: mux_23291 = 8'h0; 1: mux_23291 = v_23292;
    endcase
  endfunction
  reg [7:0] v_23292 = 8'h0;
  wire [7:0] v_23293;
  wire [7:0] v_23294;
  function [7:0] mux_23294(input [0:0] sel);
    case (sel) 0: mux_23294 = 8'h0; 1: mux_23294 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23295;
  wire [7:0] v_23296;
  wire [7:0] v_23297;
  function [7:0] mux_23297(input [0:0] sel);
    case (sel) 0: mux_23297 = 8'h0; 1: mux_23297 = v_23298;
    endcase
  endfunction
  reg [7:0] v_23298 = 8'h0;
  wire [7:0] v_23299;
  wire [7:0] v_23300;
  function [7:0] mux_23300(input [0:0] sel);
    case (sel) 0: mux_23300 = 8'h0; 1: mux_23300 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23301;
  wire [7:0] v_23302;
  wire [7:0] v_23303;
  function [7:0] mux_23303(input [0:0] sel);
    case (sel) 0: mux_23303 = 8'h0; 1: mux_23303 = v_23304;
    endcase
  endfunction
  reg [7:0] v_23304 = 8'h0;
  wire [7:0] v_23305;
  wire [7:0] v_23306;
  function [7:0] mux_23306(input [0:0] sel);
    case (sel) 0: mux_23306 = 8'h0; 1: mux_23306 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23307;
  wire [7:0] v_23308;
  wire [7:0] v_23309;
  function [7:0] mux_23309(input [0:0] sel);
    case (sel) 0: mux_23309 = 8'h0; 1: mux_23309 = v_23310;
    endcase
  endfunction
  reg [7:0] v_23310 = 8'h0;
  wire [7:0] v_23311;
  wire [7:0] v_23312;
  function [7:0] mux_23312(input [0:0] sel);
    case (sel) 0: mux_23312 = 8'h0; 1: mux_23312 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23313;
  wire [7:0] v_23314;
  wire [7:0] v_23315;
  function [7:0] mux_23315(input [0:0] sel);
    case (sel) 0: mux_23315 = 8'h0; 1: mux_23315 = v_23316;
    endcase
  endfunction
  reg [7:0] v_23316 = 8'h0;
  wire [7:0] v_23317;
  wire [7:0] v_23318;
  function [7:0] mux_23318(input [0:0] sel);
    case (sel) 0: mux_23318 = 8'h0; 1: mux_23318 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23319;
  wire [7:0] v_23320;
  wire [7:0] v_23321;
  function [7:0] mux_23321(input [0:0] sel);
    case (sel) 0: mux_23321 = 8'h0; 1: mux_23321 = v_23322;
    endcase
  endfunction
  reg [7:0] v_23322 = 8'h0;
  wire [7:0] v_23323;
  wire [7:0] v_23324;
  function [7:0] mux_23324(input [0:0] sel);
    case (sel) 0: mux_23324 = 8'h0; 1: mux_23324 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23325;
  wire [7:0] v_23326;
  wire [7:0] v_23327;
  function [7:0] mux_23327(input [0:0] sel);
    case (sel) 0: mux_23327 = 8'h0; 1: mux_23327 = v_23328;
    endcase
  endfunction
  reg [7:0] v_23328 = 8'h0;
  wire [7:0] v_23329;
  wire [7:0] v_23330;
  function [7:0] mux_23330(input [0:0] sel);
    case (sel) 0: mux_23330 = 8'h0; 1: mux_23330 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23331;
  wire [7:0] v_23332;
  wire [7:0] v_23333;
  function [7:0] mux_23333(input [0:0] sel);
    case (sel) 0: mux_23333 = 8'h0; 1: mux_23333 = vout_peek_18613;
    endcase
  endfunction
  wire [7:0] v_23334;
  function [7:0] mux_23334(input [0:0] sel);
    case (sel) 0: mux_23334 = 8'h0; 1: mux_23334 = vout_peek_18604;
    endcase
  endfunction
  wire [7:0] v_23335;
  function [7:0] mux_23335(input [0:0] sel);
    case (sel) 0: mux_23335 = 8'h0; 1: mux_23335 = v_23336;
    endcase
  endfunction
  reg [7:0] v_23336 = 8'h0;
  wire [7:0] v_23337;
  wire [7:0] v_23338;
  function [7:0] mux_23338(input [0:0] sel);
    case (sel) 0: mux_23338 = 8'h0; 1: mux_23338 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23339;
  wire [7:0] v_23340;
  wire [7:0] v_23341;
  function [7:0] mux_23341(input [0:0] sel);
    case (sel) 0: mux_23341 = 8'h0; 1: mux_23341 = vout_peek_18576;
    endcase
  endfunction
  wire [7:0] v_23342;
  function [7:0] mux_23342(input [0:0] sel);
    case (sel) 0: mux_23342 = 8'h0; 1: mux_23342 = vout_peek_18567;
    endcase
  endfunction
  wire [7:0] v_23343;
  function [7:0] mux_23343(input [0:0] sel);
    case (sel) 0: mux_23343 = 8'h0; 1: mux_23343 = v_23344;
    endcase
  endfunction
  reg [7:0] v_23344 = 8'h0;
  wire [7:0] v_23345;
  wire [7:0] v_23346;
  function [7:0] mux_23346(input [0:0] sel);
    case (sel) 0: mux_23346 = 8'h0; 1: mux_23346 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23347;
  wire [7:0] v_23348;
  wire [7:0] v_23349;
  function [7:0] mux_23349(input [0:0] sel);
    case (sel) 0: mux_23349 = 8'h0; 1: mux_23349 = v_23350;
    endcase
  endfunction
  reg [7:0] v_23350 = 8'h0;
  wire [7:0] v_23351;
  wire [7:0] v_23352;
  function [7:0] mux_23352(input [0:0] sel);
    case (sel) 0: mux_23352 = 8'h0; 1: mux_23352 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23353;
  wire [7:0] v_23354;
  wire [7:0] v_23355;
  function [7:0] mux_23355(input [0:0] sel);
    case (sel) 0: mux_23355 = 8'h0; 1: mux_23355 = vout_peek_18520;
    endcase
  endfunction
  wire [7:0] v_23356;
  function [7:0] mux_23356(input [0:0] sel);
    case (sel) 0: mux_23356 = 8'h0; 1: mux_23356 = vout_peek_18511;
    endcase
  endfunction
  wire [7:0] v_23357;
  function [7:0] mux_23357(input [0:0] sel);
    case (sel) 0: mux_23357 = 8'h0; 1: mux_23357 = v_23358;
    endcase
  endfunction
  reg [7:0] v_23358 = 8'h0;
  wire [7:0] v_23359;
  wire [7:0] v_23360;
  function [7:0] mux_23360(input [0:0] sel);
    case (sel) 0: mux_23360 = 8'h0; 1: mux_23360 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23361;
  wire [7:0] v_23362;
  wire [7:0] v_23363;
  function [7:0] mux_23363(input [0:0] sel);
    case (sel) 0: mux_23363 = 8'h0; 1: mux_23363 = vout_peek_18483;
    endcase
  endfunction
  wire [7:0] v_23364;
  function [7:0] mux_23364(input [0:0] sel);
    case (sel) 0: mux_23364 = 8'h0; 1: mux_23364 = vout_peek_18474;
    endcase
  endfunction
  wire [7:0] v_23365;
  function [7:0] mux_23365(input [0:0] sel);
    case (sel) 0: mux_23365 = 8'h0; 1: mux_23365 = v_23366;
    endcase
  endfunction
  reg [7:0] v_23366 = 8'h0;
  wire [7:0] v_23367;
  wire [7:0] v_23368;
  function [7:0] mux_23368(input [0:0] sel);
    case (sel) 0: mux_23368 = 8'h0; 1: mux_23368 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23369;
  wire [7:0] v_23370;
  wire [7:0] v_23371;
  function [7:0] mux_23371(input [0:0] sel);
    case (sel) 0: mux_23371 = 8'h0; 1: mux_23371 = v_23372;
    endcase
  endfunction
  reg [7:0] v_23372 = 8'h0;
  wire [7:0] v_23373;
  wire [7:0] v_23374;
  function [7:0] mux_23374(input [0:0] sel);
    case (sel) 0: mux_23374 = 8'h0; 1: mux_23374 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23375;
  wire [7:0] v_23376;
  wire [7:0] v_23377;
  function [7:0] mux_23377(input [0:0] sel);
    case (sel) 0: mux_23377 = 8'h0; 1: mux_23377 = v_23378;
    endcase
  endfunction
  reg [7:0] v_23378 = 8'h0;
  wire [7:0] v_23379;
  wire [7:0] v_23380;
  function [7:0] mux_23380(input [0:0] sel);
    case (sel) 0: mux_23380 = 8'h0; 1: mux_23380 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23381;
  wire [7:0] v_23382;
  wire [7:0] v_23383;
  function [7:0] mux_23383(input [0:0] sel);
    case (sel) 0: mux_23383 = 8'h0; 1: mux_23383 = vout_peek_18408;
    endcase
  endfunction
  wire [7:0] v_23384;
  function [7:0] mux_23384(input [0:0] sel);
    case (sel) 0: mux_23384 = 8'h0; 1: mux_23384 = vout_peek_18399;
    endcase
  endfunction
  wire [7:0] v_23385;
  function [7:0] mux_23385(input [0:0] sel);
    case (sel) 0: mux_23385 = 8'h0; 1: mux_23385 = v_23386;
    endcase
  endfunction
  reg [7:0] v_23386 = 8'h0;
  wire [7:0] v_23387;
  wire [7:0] v_23388;
  function [7:0] mux_23388(input [0:0] sel);
    case (sel) 0: mux_23388 = 8'h0; 1: mux_23388 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23389;
  wire [7:0] v_23390;
  wire [7:0] v_23391;
  function [7:0] mux_23391(input [0:0] sel);
    case (sel) 0: mux_23391 = 8'h0; 1: mux_23391 = vout_peek_18371;
    endcase
  endfunction
  wire [7:0] v_23392;
  function [7:0] mux_23392(input [0:0] sel);
    case (sel) 0: mux_23392 = 8'h0; 1: mux_23392 = vout_peek_18362;
    endcase
  endfunction
  wire [7:0] v_23393;
  function [7:0] mux_23393(input [0:0] sel);
    case (sel) 0: mux_23393 = 8'h0; 1: mux_23393 = v_23394;
    endcase
  endfunction
  reg [7:0] v_23394 = 8'h0;
  wire [7:0] v_23395;
  wire [7:0] v_23396;
  function [7:0] mux_23396(input [0:0] sel);
    case (sel) 0: mux_23396 = 8'h0; 1: mux_23396 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23397;
  wire [7:0] v_23398;
  wire [7:0] v_23399;
  function [7:0] mux_23399(input [0:0] sel);
    case (sel) 0: mux_23399 = 8'h0; 1: mux_23399 = v_23400;
    endcase
  endfunction
  reg [7:0] v_23400 = 8'h0;
  wire [7:0] v_23401;
  wire [7:0] v_23402;
  function [7:0] mux_23402(input [0:0] sel);
    case (sel) 0: mux_23402 = 8'h0; 1: mux_23402 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23403;
  wire [7:0] v_23404;
  wire [7:0] v_23405;
  function [7:0] mux_23405(input [0:0] sel);
    case (sel) 0: mux_23405 = 8'h0; 1: mux_23405 = vout_peek_18315;
    endcase
  endfunction
  wire [7:0] v_23406;
  function [7:0] mux_23406(input [0:0] sel);
    case (sel) 0: mux_23406 = 8'h0; 1: mux_23406 = vout_peek_18306;
    endcase
  endfunction
  wire [7:0] v_23407;
  function [7:0] mux_23407(input [0:0] sel);
    case (sel) 0: mux_23407 = 8'h0; 1: mux_23407 = v_23408;
    endcase
  endfunction
  reg [7:0] v_23408 = 8'h0;
  wire [7:0] v_23409;
  wire [7:0] v_23410;
  function [7:0] mux_23410(input [0:0] sel);
    case (sel) 0: mux_23410 = 8'h0; 1: mux_23410 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23411;
  wire [7:0] v_23412;
  wire [7:0] v_23413;
  function [7:0] mux_23413(input [0:0] sel);
    case (sel) 0: mux_23413 = 8'h0; 1: mux_23413 = vout_peek_18278;
    endcase
  endfunction
  wire [7:0] v_23414;
  function [7:0] mux_23414(input [0:0] sel);
    case (sel) 0: mux_23414 = 8'h0; 1: mux_23414 = vout_peek_18269;
    endcase
  endfunction
  wire [7:0] v_23415;
  function [7:0] mux_23415(input [0:0] sel);
    case (sel) 0: mux_23415 = 8'h0; 1: mux_23415 = v_23416;
    endcase
  endfunction
  reg [7:0] v_23416 = 8'h0;
  wire [7:0] v_23417;
  wire [7:0] v_23418;
  function [7:0] mux_23418(input [0:0] sel);
    case (sel) 0: mux_23418 = 8'h0; 1: mux_23418 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23419;
  wire [7:0] v_23420;
  wire [7:0] v_23421;
  function [7:0] mux_23421(input [0:0] sel);
    case (sel) 0: mux_23421 = 8'h0; 1: mux_23421 = v_23422;
    endcase
  endfunction
  reg [7:0] v_23422 = 8'h0;
  wire [7:0] v_23423;
  wire [7:0] v_23424;
  function [7:0] mux_23424(input [0:0] sel);
    case (sel) 0: mux_23424 = 8'h0; 1: mux_23424 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23425;
  wire [7:0] v_23426;
  wire [7:0] v_23427;
  function [7:0] mux_23427(input [0:0] sel);
    case (sel) 0: mux_23427 = 8'h0; 1: mux_23427 = v_23428;
    endcase
  endfunction
  reg [7:0] v_23428 = 8'h0;
  wire [7:0] v_23429;
  wire [7:0] v_23430;
  function [7:0] mux_23430(input [0:0] sel);
    case (sel) 0: mux_23430 = 8'h0; 1: mux_23430 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23431;
  wire [7:0] v_23432;
  wire [7:0] v_23433;
  function [7:0] mux_23433(input [0:0] sel);
    case (sel) 0: mux_23433 = 8'h0; 1: mux_23433 = v_23434;
    endcase
  endfunction
  reg [7:0] v_23434 = 8'h0;
  wire [7:0] v_23435;
  wire [7:0] v_23436;
  function [7:0] mux_23436(input [0:0] sel);
    case (sel) 0: mux_23436 = 8'h0; 1: mux_23436 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23437;
  wire [7:0] v_23438;
  wire [7:0] v_23439;
  function [7:0] mux_23439(input [0:0] sel);
    case (sel) 0: mux_23439 = 8'h0; 1: mux_23439 = vout_peek_18184;
    endcase
  endfunction
  wire [7:0] v_23440;
  function [7:0] mux_23440(input [0:0] sel);
    case (sel) 0: mux_23440 = 8'h0; 1: mux_23440 = vout_peek_18175;
    endcase
  endfunction
  wire [7:0] v_23441;
  function [7:0] mux_23441(input [0:0] sel);
    case (sel) 0: mux_23441 = 8'h0; 1: mux_23441 = v_23442;
    endcase
  endfunction
  reg [7:0] v_23442 = 8'h0;
  wire [7:0] v_23443;
  wire [7:0] v_23444;
  function [7:0] mux_23444(input [0:0] sel);
    case (sel) 0: mux_23444 = 8'h0; 1: mux_23444 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23445;
  wire [7:0] v_23446;
  wire [7:0] v_23447;
  function [7:0] mux_23447(input [0:0] sel);
    case (sel) 0: mux_23447 = 8'h0; 1: mux_23447 = vout_peek_18147;
    endcase
  endfunction
  wire [7:0] v_23448;
  function [7:0] mux_23448(input [0:0] sel);
    case (sel) 0: mux_23448 = 8'h0; 1: mux_23448 = vout_peek_18138;
    endcase
  endfunction
  wire [7:0] v_23449;
  function [7:0] mux_23449(input [0:0] sel);
    case (sel) 0: mux_23449 = 8'h0; 1: mux_23449 = v_23450;
    endcase
  endfunction
  reg [7:0] v_23450 = 8'h0;
  wire [7:0] v_23451;
  wire [7:0] v_23452;
  function [7:0] mux_23452(input [0:0] sel);
    case (sel) 0: mux_23452 = 8'h0; 1: mux_23452 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23453;
  wire [7:0] v_23454;
  wire [7:0] v_23455;
  function [7:0] mux_23455(input [0:0] sel);
    case (sel) 0: mux_23455 = 8'h0; 1: mux_23455 = v_23456;
    endcase
  endfunction
  reg [7:0] v_23456 = 8'h0;
  wire [7:0] v_23457;
  wire [7:0] v_23458;
  function [7:0] mux_23458(input [0:0] sel);
    case (sel) 0: mux_23458 = 8'h0; 1: mux_23458 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23459;
  wire [7:0] v_23460;
  wire [7:0] v_23461;
  function [7:0] mux_23461(input [0:0] sel);
    case (sel) 0: mux_23461 = 8'h0; 1: mux_23461 = vout_peek_18091;
    endcase
  endfunction
  wire [7:0] v_23462;
  function [7:0] mux_23462(input [0:0] sel);
    case (sel) 0: mux_23462 = 8'h0; 1: mux_23462 = vout_peek_18082;
    endcase
  endfunction
  wire [7:0] v_23463;
  function [7:0] mux_23463(input [0:0] sel);
    case (sel) 0: mux_23463 = 8'h0; 1: mux_23463 = v_23464;
    endcase
  endfunction
  reg [7:0] v_23464 = 8'h0;
  wire [7:0] v_23465;
  wire [7:0] v_23466;
  function [7:0] mux_23466(input [0:0] sel);
    case (sel) 0: mux_23466 = 8'h0; 1: mux_23466 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23467;
  wire [7:0] v_23468;
  wire [7:0] v_23469;
  function [7:0] mux_23469(input [0:0] sel);
    case (sel) 0: mux_23469 = 8'h0; 1: mux_23469 = vout_peek_18054;
    endcase
  endfunction
  wire [7:0] v_23470;
  function [7:0] mux_23470(input [0:0] sel);
    case (sel) 0: mux_23470 = 8'h0; 1: mux_23470 = vout_peek_18045;
    endcase
  endfunction
  wire [7:0] v_23471;
  function [7:0] mux_23471(input [0:0] sel);
    case (sel) 0: mux_23471 = 8'h0; 1: mux_23471 = v_23472;
    endcase
  endfunction
  reg [7:0] v_23472 = 8'h0;
  wire [7:0] v_23473;
  wire [7:0] v_23474;
  function [7:0] mux_23474(input [0:0] sel);
    case (sel) 0: mux_23474 = 8'h0; 1: mux_23474 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23475;
  wire [7:0] v_23476;
  wire [7:0] v_23477;
  function [7:0] mux_23477(input [0:0] sel);
    case (sel) 0: mux_23477 = 8'h0; 1: mux_23477 = v_23478;
    endcase
  endfunction
  reg [7:0] v_23478 = 8'h0;
  wire [7:0] v_23479;
  wire [7:0] v_23480;
  function [7:0] mux_23480(input [0:0] sel);
    case (sel) 0: mux_23480 = 8'h0; 1: mux_23480 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23481;
  wire [7:0] v_23482;
  wire [7:0] v_23483;
  function [7:0] mux_23483(input [0:0] sel);
    case (sel) 0: mux_23483 = 8'h0; 1: mux_23483 = v_23484;
    endcase
  endfunction
  reg [7:0] v_23484 = 8'h0;
  wire [7:0] v_23485;
  wire [7:0] v_23486;
  function [7:0] mux_23486(input [0:0] sel);
    case (sel) 0: mux_23486 = 8'h0; 1: mux_23486 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23487;
  wire [7:0] v_23488;
  wire [7:0] v_23489;
  function [7:0] mux_23489(input [0:0] sel);
    case (sel) 0: mux_23489 = 8'h0; 1: mux_23489 = vout_peek_17979;
    endcase
  endfunction
  wire [7:0] v_23490;
  function [7:0] mux_23490(input [0:0] sel);
    case (sel) 0: mux_23490 = 8'h0; 1: mux_23490 = vout_peek_17970;
    endcase
  endfunction
  wire [7:0] v_23491;
  function [7:0] mux_23491(input [0:0] sel);
    case (sel) 0: mux_23491 = 8'h0; 1: mux_23491 = v_23492;
    endcase
  endfunction
  reg [7:0] v_23492 = 8'h0;
  wire [7:0] v_23493;
  wire [7:0] v_23494;
  function [7:0] mux_23494(input [0:0] sel);
    case (sel) 0: mux_23494 = 8'h0; 1: mux_23494 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23495;
  wire [7:0] v_23496;
  wire [7:0] v_23497;
  function [7:0] mux_23497(input [0:0] sel);
    case (sel) 0: mux_23497 = 8'h0; 1: mux_23497 = vout_peek_17942;
    endcase
  endfunction
  wire [7:0] v_23498;
  function [7:0] mux_23498(input [0:0] sel);
    case (sel) 0: mux_23498 = 8'h0; 1: mux_23498 = vout_peek_17933;
    endcase
  endfunction
  wire [7:0] v_23499;
  function [7:0] mux_23499(input [0:0] sel);
    case (sel) 0: mux_23499 = 8'h0; 1: mux_23499 = v_23500;
    endcase
  endfunction
  reg [7:0] v_23500 = 8'h0;
  wire [7:0] v_23501;
  wire [7:0] v_23502;
  function [7:0] mux_23502(input [0:0] sel);
    case (sel) 0: mux_23502 = 8'h0; 1: mux_23502 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23503;
  wire [7:0] v_23504;
  wire [7:0] v_23505;
  function [7:0] mux_23505(input [0:0] sel);
    case (sel) 0: mux_23505 = 8'h0; 1: mux_23505 = v_23506;
    endcase
  endfunction
  reg [7:0] v_23506 = 8'h0;
  wire [7:0] v_23507;
  wire [7:0] v_23508;
  function [7:0] mux_23508(input [0:0] sel);
    case (sel) 0: mux_23508 = 8'h0; 1: mux_23508 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23509;
  wire [7:0] v_23510;
  wire [7:0] v_23511;
  function [7:0] mux_23511(input [0:0] sel);
    case (sel) 0: mux_23511 = 8'h0; 1: mux_23511 = vout_peek_17886;
    endcase
  endfunction
  wire [7:0] v_23512;
  function [7:0] mux_23512(input [0:0] sel);
    case (sel) 0: mux_23512 = 8'h0; 1: mux_23512 = vout_peek_17877;
    endcase
  endfunction
  wire [7:0] v_23513;
  function [7:0] mux_23513(input [0:0] sel);
    case (sel) 0: mux_23513 = 8'h0; 1: mux_23513 = v_23514;
    endcase
  endfunction
  reg [7:0] v_23514 = 8'h0;
  wire [7:0] v_23515;
  wire [7:0] v_23516;
  function [7:0] mux_23516(input [0:0] sel);
    case (sel) 0: mux_23516 = 8'h0; 1: mux_23516 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23517;
  wire [7:0] v_23518;
  wire [7:0] v_23519;
  function [7:0] mux_23519(input [0:0] sel);
    case (sel) 0: mux_23519 = 8'h0; 1: mux_23519 = vout_peek_17849;
    endcase
  endfunction
  wire [7:0] v_23520;
  function [7:0] mux_23520(input [0:0] sel);
    case (sel) 0: mux_23520 = 8'h0; 1: mux_23520 = vout_peek_17840;
    endcase
  endfunction
  wire [7:0] v_23521;
  function [7:0] mux_23521(input [0:0] sel);
    case (sel) 0: mux_23521 = 8'h0; 1: mux_23521 = v_23522;
    endcase
  endfunction
  reg [7:0] v_23522 = 8'h0;
  wire [7:0] v_23523;
  wire [7:0] v_23524;
  function [7:0] mux_23524(input [0:0] sel);
    case (sel) 0: mux_23524 = 8'h0; 1: mux_23524 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23525;
  wire [7:0] v_23526;
  wire [7:0] v_23527;
  function [7:0] mux_23527(input [0:0] sel);
    case (sel) 0: mux_23527 = 8'h0; 1: mux_23527 = v_23528;
    endcase
  endfunction
  reg [7:0] v_23528 = 8'h0;
  wire [7:0] v_23529;
  wire [7:0] v_23530;
  function [7:0] mux_23530(input [0:0] sel);
    case (sel) 0: mux_23530 = 8'h0; 1: mux_23530 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23531;
  wire [7:0] v_23532;
  wire [7:0] v_23533;
  function [7:0] mux_23533(input [0:0] sel);
    case (sel) 0: mux_23533 = 8'h0; 1: mux_23533 = v_23534;
    endcase
  endfunction
  reg [7:0] v_23534 = 8'h0;
  wire [7:0] v_23535;
  wire [7:0] v_23536;
  function [7:0] mux_23536(input [0:0] sel);
    case (sel) 0: mux_23536 = 8'h0; 1: mux_23536 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23537;
  wire [7:0] v_23538;
  wire [7:0] v_23539;
  function [7:0] mux_23539(input [0:0] sel);
    case (sel) 0: mux_23539 = 8'h0; 1: mux_23539 = v_23540;
    endcase
  endfunction
  reg [7:0] v_23540 = 8'h0;
  wire [7:0] v_23541;
  wire [7:0] v_23542;
  function [7:0] mux_23542(input [0:0] sel);
    case (sel) 0: mux_23542 = 8'h0; 1: mux_23542 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23543;
  wire [7:0] v_23544;
  wire [7:0] v_23545;
  function [7:0] mux_23545(input [0:0] sel);
    case (sel) 0: mux_23545 = 8'h0; 1: mux_23545 = v_23546;
    endcase
  endfunction
  reg [7:0] v_23546 = 8'h0;
  wire [7:0] v_23547;
  wire [7:0] v_23548;
  function [7:0] mux_23548(input [0:0] sel);
    case (sel) 0: mux_23548 = 8'h0; 1: mux_23548 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23549;
  wire [7:0] v_23550;
  wire [7:0] v_23551;
  function [7:0] mux_23551(input [0:0] sel);
    case (sel) 0: mux_23551 = 8'h0; 1: mux_23551 = vout_peek_17736;
    endcase
  endfunction
  wire [7:0] v_23552;
  function [7:0] mux_23552(input [0:0] sel);
    case (sel) 0: mux_23552 = 8'h0; 1: mux_23552 = vout_peek_17727;
    endcase
  endfunction
  wire [7:0] v_23553;
  function [7:0] mux_23553(input [0:0] sel);
    case (sel) 0: mux_23553 = 8'h0; 1: mux_23553 = v_23554;
    endcase
  endfunction
  reg [7:0] v_23554 = 8'h0;
  wire [7:0] v_23555;
  wire [7:0] v_23556;
  function [7:0] mux_23556(input [0:0] sel);
    case (sel) 0: mux_23556 = 8'h0; 1: mux_23556 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23557;
  wire [7:0] v_23558;
  wire [7:0] v_23559;
  function [7:0] mux_23559(input [0:0] sel);
    case (sel) 0: mux_23559 = 8'h0; 1: mux_23559 = vout_peek_17699;
    endcase
  endfunction
  wire [7:0] v_23560;
  function [7:0] mux_23560(input [0:0] sel);
    case (sel) 0: mux_23560 = 8'h0; 1: mux_23560 = vout_peek_17690;
    endcase
  endfunction
  wire [7:0] v_23561;
  function [7:0] mux_23561(input [0:0] sel);
    case (sel) 0: mux_23561 = 8'h0; 1: mux_23561 = v_23562;
    endcase
  endfunction
  reg [7:0] v_23562 = 8'h0;
  wire [7:0] v_23563;
  wire [7:0] v_23564;
  function [7:0] mux_23564(input [0:0] sel);
    case (sel) 0: mux_23564 = 8'h0; 1: mux_23564 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23565;
  wire [7:0] v_23566;
  wire [7:0] v_23567;
  function [7:0] mux_23567(input [0:0] sel);
    case (sel) 0: mux_23567 = 8'h0; 1: mux_23567 = v_23568;
    endcase
  endfunction
  reg [7:0] v_23568 = 8'h0;
  wire [7:0] v_23569;
  wire [7:0] v_23570;
  function [7:0] mux_23570(input [0:0] sel);
    case (sel) 0: mux_23570 = 8'h0; 1: mux_23570 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23571;
  wire [7:0] v_23572;
  wire [7:0] v_23573;
  function [7:0] mux_23573(input [0:0] sel);
    case (sel) 0: mux_23573 = 8'h0; 1: mux_23573 = vout_peek_17643;
    endcase
  endfunction
  wire [7:0] v_23574;
  function [7:0] mux_23574(input [0:0] sel);
    case (sel) 0: mux_23574 = 8'h0; 1: mux_23574 = vout_peek_17634;
    endcase
  endfunction
  wire [7:0] v_23575;
  function [7:0] mux_23575(input [0:0] sel);
    case (sel) 0: mux_23575 = 8'h0; 1: mux_23575 = v_23576;
    endcase
  endfunction
  reg [7:0] v_23576 = 8'h0;
  wire [7:0] v_23577;
  wire [7:0] v_23578;
  function [7:0] mux_23578(input [0:0] sel);
    case (sel) 0: mux_23578 = 8'h0; 1: mux_23578 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23579;
  wire [7:0] v_23580;
  wire [7:0] v_23581;
  function [7:0] mux_23581(input [0:0] sel);
    case (sel) 0: mux_23581 = 8'h0; 1: mux_23581 = vout_peek_17606;
    endcase
  endfunction
  wire [7:0] v_23582;
  function [7:0] mux_23582(input [0:0] sel);
    case (sel) 0: mux_23582 = 8'h0; 1: mux_23582 = vout_peek_17597;
    endcase
  endfunction
  wire [7:0] v_23583;
  function [7:0] mux_23583(input [0:0] sel);
    case (sel) 0: mux_23583 = 8'h0; 1: mux_23583 = v_23584;
    endcase
  endfunction
  reg [7:0] v_23584 = 8'h0;
  wire [7:0] v_23585;
  wire [7:0] v_23586;
  function [7:0] mux_23586(input [0:0] sel);
    case (sel) 0: mux_23586 = 8'h0; 1: mux_23586 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23587;
  wire [7:0] v_23588;
  wire [7:0] v_23589;
  function [7:0] mux_23589(input [0:0] sel);
    case (sel) 0: mux_23589 = 8'h0; 1: mux_23589 = v_23590;
    endcase
  endfunction
  reg [7:0] v_23590 = 8'h0;
  wire [7:0] v_23591;
  wire [7:0] v_23592;
  function [7:0] mux_23592(input [0:0] sel);
    case (sel) 0: mux_23592 = 8'h0; 1: mux_23592 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23593;
  wire [7:0] v_23594;
  wire [7:0] v_23595;
  function [7:0] mux_23595(input [0:0] sel);
    case (sel) 0: mux_23595 = 8'h0; 1: mux_23595 = v_23596;
    endcase
  endfunction
  reg [7:0] v_23596 = 8'h0;
  wire [7:0] v_23597;
  wire [7:0] v_23598;
  function [7:0] mux_23598(input [0:0] sel);
    case (sel) 0: mux_23598 = 8'h0; 1: mux_23598 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23599;
  wire [7:0] v_23600;
  wire [7:0] v_23601;
  function [7:0] mux_23601(input [0:0] sel);
    case (sel) 0: mux_23601 = 8'h0; 1: mux_23601 = vout_peek_17531;
    endcase
  endfunction
  wire [7:0] v_23602;
  function [7:0] mux_23602(input [0:0] sel);
    case (sel) 0: mux_23602 = 8'h0; 1: mux_23602 = vout_peek_17522;
    endcase
  endfunction
  wire [7:0] v_23603;
  function [7:0] mux_23603(input [0:0] sel);
    case (sel) 0: mux_23603 = 8'h0; 1: mux_23603 = v_23604;
    endcase
  endfunction
  reg [7:0] v_23604 = 8'h0;
  wire [7:0] v_23605;
  wire [7:0] v_23606;
  function [7:0] mux_23606(input [0:0] sel);
    case (sel) 0: mux_23606 = 8'h0; 1: mux_23606 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23607;
  wire [7:0] v_23608;
  wire [7:0] v_23609;
  function [7:0] mux_23609(input [0:0] sel);
    case (sel) 0: mux_23609 = 8'h0; 1: mux_23609 = vout_peek_17494;
    endcase
  endfunction
  wire [7:0] v_23610;
  function [7:0] mux_23610(input [0:0] sel);
    case (sel) 0: mux_23610 = 8'h0; 1: mux_23610 = vout_peek_17485;
    endcase
  endfunction
  wire [7:0] v_23611;
  function [7:0] mux_23611(input [0:0] sel);
    case (sel) 0: mux_23611 = 8'h0; 1: mux_23611 = v_23612;
    endcase
  endfunction
  reg [7:0] v_23612 = 8'h0;
  wire [7:0] v_23613;
  wire [7:0] v_23614;
  function [7:0] mux_23614(input [0:0] sel);
    case (sel) 0: mux_23614 = 8'h0; 1: mux_23614 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23615;
  wire [7:0] v_23616;
  wire [7:0] v_23617;
  function [7:0] mux_23617(input [0:0] sel);
    case (sel) 0: mux_23617 = 8'h0; 1: mux_23617 = v_23618;
    endcase
  endfunction
  reg [7:0] v_23618 = 8'h0;
  wire [7:0] v_23619;
  wire [7:0] v_23620;
  function [7:0] mux_23620(input [0:0] sel);
    case (sel) 0: mux_23620 = 8'h0; 1: mux_23620 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23621;
  wire [7:0] v_23622;
  wire [7:0] v_23623;
  function [7:0] mux_23623(input [0:0] sel);
    case (sel) 0: mux_23623 = 8'h0; 1: mux_23623 = vout_peek_17438;
    endcase
  endfunction
  wire [7:0] v_23624;
  function [7:0] mux_23624(input [0:0] sel);
    case (sel) 0: mux_23624 = 8'h0; 1: mux_23624 = vout_peek_17429;
    endcase
  endfunction
  wire [7:0] v_23625;
  function [7:0] mux_23625(input [0:0] sel);
    case (sel) 0: mux_23625 = 8'h0; 1: mux_23625 = v_23626;
    endcase
  endfunction
  reg [7:0] v_23626 = 8'h0;
  wire [7:0] v_23627;
  wire [7:0] v_23628;
  function [7:0] mux_23628(input [0:0] sel);
    case (sel) 0: mux_23628 = 8'h0; 1: mux_23628 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23629;
  wire [7:0] v_23630;
  wire [7:0] v_23631;
  function [7:0] mux_23631(input [0:0] sel);
    case (sel) 0: mux_23631 = 8'h0; 1: mux_23631 = vout_peek_17401;
    endcase
  endfunction
  wire [7:0] v_23632;
  function [7:0] mux_23632(input [0:0] sel);
    case (sel) 0: mux_23632 = 8'h0; 1: mux_23632 = vout_peek_17392;
    endcase
  endfunction
  wire [7:0] v_23633;
  function [7:0] mux_23633(input [0:0] sel);
    case (sel) 0: mux_23633 = 8'h0; 1: mux_23633 = v_23634;
    endcase
  endfunction
  reg [7:0] v_23634 = 8'h0;
  wire [7:0] v_23635;
  wire [7:0] v_23636;
  function [7:0] mux_23636(input [0:0] sel);
    case (sel) 0: mux_23636 = 8'h0; 1: mux_23636 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23637;
  wire [7:0] v_23638;
  wire [7:0] v_23639;
  function [7:0] mux_23639(input [0:0] sel);
    case (sel) 0: mux_23639 = 8'h0; 1: mux_23639 = v_23640;
    endcase
  endfunction
  reg [7:0] v_23640 = 8'h0;
  wire [7:0] v_23641;
  wire [7:0] v_23642;
  function [7:0] mux_23642(input [0:0] sel);
    case (sel) 0: mux_23642 = 8'h0; 1: mux_23642 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23643;
  wire [7:0] v_23644;
  wire [7:0] v_23645;
  function [7:0] mux_23645(input [0:0] sel);
    case (sel) 0: mux_23645 = 8'h0; 1: mux_23645 = v_23646;
    endcase
  endfunction
  reg [7:0] v_23646 = 8'h0;
  wire [7:0] v_23647;
  wire [7:0] v_23648;
  function [7:0] mux_23648(input [0:0] sel);
    case (sel) 0: mux_23648 = 8'h0; 1: mux_23648 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23649;
  wire [7:0] v_23650;
  wire [7:0] v_23651;
  function [7:0] mux_23651(input [0:0] sel);
    case (sel) 0: mux_23651 = 8'h0; 1: mux_23651 = v_23652;
    endcase
  endfunction
  reg [7:0] v_23652 = 8'h0;
  wire [7:0] v_23653;
  wire [7:0] v_23654;
  function [7:0] mux_23654(input [0:0] sel);
    case (sel) 0: mux_23654 = 8'h0; 1: mux_23654 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23655;
  wire [7:0] v_23656;
  wire [7:0] v_23657;
  function [7:0] mux_23657(input [0:0] sel);
    case (sel) 0: mux_23657 = 8'h0; 1: mux_23657 = vout_peek_17307;
    endcase
  endfunction
  wire [7:0] v_23658;
  function [7:0] mux_23658(input [0:0] sel);
    case (sel) 0: mux_23658 = 8'h0; 1: mux_23658 = vout_peek_17298;
    endcase
  endfunction
  wire [7:0] v_23659;
  function [7:0] mux_23659(input [0:0] sel);
    case (sel) 0: mux_23659 = 8'h0; 1: mux_23659 = v_23660;
    endcase
  endfunction
  reg [7:0] v_23660 = 8'h0;
  wire [7:0] v_23661;
  wire [7:0] v_23662;
  function [7:0] mux_23662(input [0:0] sel);
    case (sel) 0: mux_23662 = 8'h0; 1: mux_23662 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23663;
  wire [7:0] v_23664;
  wire [7:0] v_23665;
  function [7:0] mux_23665(input [0:0] sel);
    case (sel) 0: mux_23665 = 8'h0; 1: mux_23665 = vout_peek_17270;
    endcase
  endfunction
  wire [7:0] v_23666;
  function [7:0] mux_23666(input [0:0] sel);
    case (sel) 0: mux_23666 = 8'h0; 1: mux_23666 = vout_peek_17261;
    endcase
  endfunction
  wire [7:0] v_23667;
  function [7:0] mux_23667(input [0:0] sel);
    case (sel) 0: mux_23667 = 8'h0; 1: mux_23667 = v_23668;
    endcase
  endfunction
  reg [7:0] v_23668 = 8'h0;
  wire [7:0] v_23669;
  wire [7:0] v_23670;
  function [7:0] mux_23670(input [0:0] sel);
    case (sel) 0: mux_23670 = 8'h0; 1: mux_23670 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23671;
  wire [7:0] v_23672;
  wire [7:0] v_23673;
  function [7:0] mux_23673(input [0:0] sel);
    case (sel) 0: mux_23673 = 8'h0; 1: mux_23673 = v_23674;
    endcase
  endfunction
  reg [7:0] v_23674 = 8'h0;
  wire [7:0] v_23675;
  wire [7:0] v_23676;
  function [7:0] mux_23676(input [0:0] sel);
    case (sel) 0: mux_23676 = 8'h0; 1: mux_23676 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23677;
  wire [7:0] v_23678;
  wire [7:0] v_23679;
  function [7:0] mux_23679(input [0:0] sel);
    case (sel) 0: mux_23679 = 8'h0; 1: mux_23679 = vout_peek_17214;
    endcase
  endfunction
  wire [7:0] v_23680;
  function [7:0] mux_23680(input [0:0] sel);
    case (sel) 0: mux_23680 = 8'h0; 1: mux_23680 = vout_peek_17205;
    endcase
  endfunction
  wire [7:0] v_23681;
  function [7:0] mux_23681(input [0:0] sel);
    case (sel) 0: mux_23681 = 8'h0; 1: mux_23681 = v_23682;
    endcase
  endfunction
  reg [7:0] v_23682 = 8'h0;
  wire [7:0] v_23683;
  wire [7:0] v_23684;
  function [7:0] mux_23684(input [0:0] sel);
    case (sel) 0: mux_23684 = 8'h0; 1: mux_23684 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23685;
  wire [7:0] v_23686;
  wire [7:0] v_23687;
  function [7:0] mux_23687(input [0:0] sel);
    case (sel) 0: mux_23687 = 8'h0; 1: mux_23687 = vout_peek_17177;
    endcase
  endfunction
  wire [7:0] v_23688;
  function [7:0] mux_23688(input [0:0] sel);
    case (sel) 0: mux_23688 = 8'h0; 1: mux_23688 = vout_peek_17168;
    endcase
  endfunction
  wire [7:0] v_23689;
  function [7:0] mux_23689(input [0:0] sel);
    case (sel) 0: mux_23689 = 8'h0; 1: mux_23689 = v_23690;
    endcase
  endfunction
  reg [7:0] v_23690 = 8'h0;
  wire [7:0] v_23691;
  wire [7:0] v_23692;
  function [7:0] mux_23692(input [0:0] sel);
    case (sel) 0: mux_23692 = 8'h0; 1: mux_23692 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23693;
  wire [7:0] v_23694;
  wire [7:0] v_23695;
  function [7:0] mux_23695(input [0:0] sel);
    case (sel) 0: mux_23695 = 8'h0; 1: mux_23695 = v_23696;
    endcase
  endfunction
  reg [7:0] v_23696 = 8'h0;
  wire [7:0] v_23697;
  wire [7:0] v_23698;
  function [7:0] mux_23698(input [0:0] sel);
    case (sel) 0: mux_23698 = 8'h0; 1: mux_23698 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23699;
  wire [7:0] v_23700;
  wire [7:0] v_23701;
  function [7:0] mux_23701(input [0:0] sel);
    case (sel) 0: mux_23701 = 8'h0; 1: mux_23701 = v_23702;
    endcase
  endfunction
  reg [7:0] v_23702 = 8'h0;
  wire [7:0] v_23703;
  wire [7:0] v_23704;
  function [7:0] mux_23704(input [0:0] sel);
    case (sel) 0: mux_23704 = 8'h0; 1: mux_23704 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23705;
  wire [7:0] v_23706;
  wire [7:0] v_23707;
  function [7:0] mux_23707(input [0:0] sel);
    case (sel) 0: mux_23707 = 8'h0; 1: mux_23707 = vout_peek_17102;
    endcase
  endfunction
  wire [7:0] v_23708;
  function [7:0] mux_23708(input [0:0] sel);
    case (sel) 0: mux_23708 = 8'h0; 1: mux_23708 = vout_peek_17093;
    endcase
  endfunction
  wire [7:0] v_23709;
  function [7:0] mux_23709(input [0:0] sel);
    case (sel) 0: mux_23709 = 8'h0; 1: mux_23709 = v_23710;
    endcase
  endfunction
  reg [7:0] v_23710 = 8'h0;
  wire [7:0] v_23711;
  wire [7:0] v_23712;
  function [7:0] mux_23712(input [0:0] sel);
    case (sel) 0: mux_23712 = 8'h0; 1: mux_23712 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23713;
  wire [7:0] v_23714;
  wire [7:0] v_23715;
  function [7:0] mux_23715(input [0:0] sel);
    case (sel) 0: mux_23715 = 8'h0; 1: mux_23715 = vout_peek_17065;
    endcase
  endfunction
  wire [7:0] v_23716;
  function [7:0] mux_23716(input [0:0] sel);
    case (sel) 0: mux_23716 = 8'h0; 1: mux_23716 = vout_peek_17056;
    endcase
  endfunction
  wire [7:0] v_23717;
  function [7:0] mux_23717(input [0:0] sel);
    case (sel) 0: mux_23717 = 8'h0; 1: mux_23717 = v_23718;
    endcase
  endfunction
  reg [7:0] v_23718 = 8'h0;
  wire [7:0] v_23719;
  wire [7:0] v_23720;
  function [7:0] mux_23720(input [0:0] sel);
    case (sel) 0: mux_23720 = 8'h0; 1: mux_23720 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23721;
  wire [7:0] v_23722;
  wire [7:0] v_23723;
  function [7:0] mux_23723(input [0:0] sel);
    case (sel) 0: mux_23723 = 8'h0; 1: mux_23723 = v_23724;
    endcase
  endfunction
  reg [7:0] v_23724 = 8'h0;
  wire [7:0] v_23725;
  wire [7:0] v_23726;
  function [7:0] mux_23726(input [0:0] sel);
    case (sel) 0: mux_23726 = 8'h0; 1: mux_23726 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23727;
  wire [7:0] v_23728;
  wire [7:0] v_23729;
  function [7:0] mux_23729(input [0:0] sel);
    case (sel) 0: mux_23729 = 8'h0; 1: mux_23729 = vout_peek_17009;
    endcase
  endfunction
  wire [7:0] v_23730;
  function [7:0] mux_23730(input [0:0] sel);
    case (sel) 0: mux_23730 = 8'h0; 1: mux_23730 = vout_peek_17000;
    endcase
  endfunction
  wire [7:0] v_23731;
  function [7:0] mux_23731(input [0:0] sel);
    case (sel) 0: mux_23731 = 8'h0; 1: mux_23731 = v_23732;
    endcase
  endfunction
  reg [7:0] v_23732 = 8'h0;
  wire [7:0] v_23733;
  wire [7:0] v_23734;
  function [7:0] mux_23734(input [0:0] sel);
    case (sel) 0: mux_23734 = 8'h0; 1: mux_23734 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23735;
  wire [7:0] v_23736;
  wire [7:0] v_23737;
  function [7:0] mux_23737(input [0:0] sel);
    case (sel) 0: mux_23737 = 8'h0; 1: mux_23737 = vout_peek_16972;
    endcase
  endfunction
  wire [7:0] v_23738;
  function [7:0] mux_23738(input [0:0] sel);
    case (sel) 0: mux_23738 = 8'h0; 1: mux_23738 = vout_peek_16963;
    endcase
  endfunction
  wire [7:0] v_23739;
  function [7:0] mux_23739(input [0:0] sel);
    case (sel) 0: mux_23739 = 8'h0; 1: mux_23739 = v_23740;
    endcase
  endfunction
  reg [7:0] v_23740 = 8'h0;
  wire [7:0] v_23741;
  wire [7:0] v_23742;
  function [7:0] mux_23742(input [0:0] sel);
    case (sel) 0: mux_23742 = 8'h0; 1: mux_23742 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23743;
  wire [7:0] v_23744;
  wire [7:0] v_23745;
  function [7:0] mux_23745(input [0:0] sel);
    case (sel) 0: mux_23745 = 8'h0; 1: mux_23745 = v_23746;
    endcase
  endfunction
  reg [7:0] v_23746 = 8'h0;
  wire [7:0] v_23747;
  wire [7:0] v_23748;
  function [7:0] mux_23748(input [0:0] sel);
    case (sel) 0: mux_23748 = 8'h0; 1: mux_23748 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23749;
  wire [7:0] v_23750;
  wire [7:0] v_23751;
  function [7:0] mux_23751(input [0:0] sel);
    case (sel) 0: mux_23751 = 8'h0; 1: mux_23751 = v_23752;
    endcase
  endfunction
  reg [7:0] v_23752 = 8'h0;
  wire [7:0] v_23753;
  wire [7:0] v_23754;
  function [7:0] mux_23754(input [0:0] sel);
    case (sel) 0: mux_23754 = 8'h0; 1: mux_23754 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23755;
  wire [7:0] v_23756;
  wire [7:0] v_23757;
  function [7:0] mux_23757(input [0:0] sel);
    case (sel) 0: mux_23757 = 8'h0; 1: mux_23757 = v_23758;
    endcase
  endfunction
  reg [7:0] v_23758 = 8'h0;
  wire [7:0] v_23759;
  wire [7:0] v_23760;
  function [7:0] mux_23760(input [0:0] sel);
    case (sel) 0: mux_23760 = 8'h0; 1: mux_23760 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23761;
  wire [7:0] v_23762;
  wire [7:0] v_23763;
  function [7:0] mux_23763(input [0:0] sel);
    case (sel) 0: mux_23763 = 8'h0; 1: mux_23763 = v_23764;
    endcase
  endfunction
  reg [7:0] v_23764 = 8'h0;
  wire [7:0] v_23765;
  wire [7:0] v_23766;
  function [7:0] mux_23766(input [0:0] sel);
    case (sel) 0: mux_23766 = 8'h0; 1: mux_23766 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23767;
  wire [7:0] v_23768;
  wire [7:0] v_23769;
  function [7:0] mux_23769(input [0:0] sel);
    case (sel) 0: mux_23769 = 8'h0; 1: mux_23769 = v_23770;
    endcase
  endfunction
  reg [7:0] v_23770 = 8'h0;
  wire [7:0] v_23771;
  wire [7:0] v_23772;
  function [7:0] mux_23772(input [0:0] sel);
    case (sel) 0: mux_23772 = 8'h0; 1: mux_23772 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23773;
  wire [7:0] v_23774;
  wire [7:0] v_23775;
  function [7:0] mux_23775(input [0:0] sel);
    case (sel) 0: mux_23775 = 8'h0; 1: mux_23775 = vout_peek_16840;
    endcase
  endfunction
  wire [7:0] v_23776;
  function [7:0] mux_23776(input [0:0] sel);
    case (sel) 0: mux_23776 = 8'h0; 1: mux_23776 = vout_peek_16831;
    endcase
  endfunction
  wire [7:0] v_23777;
  function [7:0] mux_23777(input [0:0] sel);
    case (sel) 0: mux_23777 = 8'h0; 1: mux_23777 = v_23778;
    endcase
  endfunction
  reg [7:0] v_23778 = 8'h0;
  wire [7:0] v_23779;
  wire [7:0] v_23780;
  function [7:0] mux_23780(input [0:0] sel);
    case (sel) 0: mux_23780 = 8'h0; 1: mux_23780 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23781;
  wire [7:0] v_23782;
  wire [7:0] v_23783;
  function [7:0] mux_23783(input [0:0] sel);
    case (sel) 0: mux_23783 = 8'h0; 1: mux_23783 = vout_peek_16803;
    endcase
  endfunction
  wire [7:0] v_23784;
  function [7:0] mux_23784(input [0:0] sel);
    case (sel) 0: mux_23784 = 8'h0; 1: mux_23784 = vout_peek_16794;
    endcase
  endfunction
  wire [7:0] v_23785;
  function [7:0] mux_23785(input [0:0] sel);
    case (sel) 0: mux_23785 = 8'h0; 1: mux_23785 = v_23786;
    endcase
  endfunction
  reg [7:0] v_23786 = 8'h0;
  wire [7:0] v_23787;
  wire [7:0] v_23788;
  function [7:0] mux_23788(input [0:0] sel);
    case (sel) 0: mux_23788 = 8'h0; 1: mux_23788 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23789;
  wire [7:0] v_23790;
  wire [7:0] v_23791;
  function [7:0] mux_23791(input [0:0] sel);
    case (sel) 0: mux_23791 = 8'h0; 1: mux_23791 = v_23792;
    endcase
  endfunction
  reg [7:0] v_23792 = 8'h0;
  wire [7:0] v_23793;
  wire [7:0] v_23794;
  function [7:0] mux_23794(input [0:0] sel);
    case (sel) 0: mux_23794 = 8'h0; 1: mux_23794 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23795;
  wire [7:0] v_23796;
  wire [7:0] v_23797;
  function [7:0] mux_23797(input [0:0] sel);
    case (sel) 0: mux_23797 = 8'h0; 1: mux_23797 = vout_peek_16747;
    endcase
  endfunction
  wire [7:0] v_23798;
  function [7:0] mux_23798(input [0:0] sel);
    case (sel) 0: mux_23798 = 8'h0; 1: mux_23798 = vout_peek_16738;
    endcase
  endfunction
  wire [7:0] v_23799;
  function [7:0] mux_23799(input [0:0] sel);
    case (sel) 0: mux_23799 = 8'h0; 1: mux_23799 = v_23800;
    endcase
  endfunction
  reg [7:0] v_23800 = 8'h0;
  wire [7:0] v_23801;
  wire [7:0] v_23802;
  function [7:0] mux_23802(input [0:0] sel);
    case (sel) 0: mux_23802 = 8'h0; 1: mux_23802 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23803;
  wire [7:0] v_23804;
  wire [7:0] v_23805;
  function [7:0] mux_23805(input [0:0] sel);
    case (sel) 0: mux_23805 = 8'h0; 1: mux_23805 = vout_peek_16710;
    endcase
  endfunction
  wire [7:0] v_23806;
  function [7:0] mux_23806(input [0:0] sel);
    case (sel) 0: mux_23806 = 8'h0; 1: mux_23806 = vout_peek_16701;
    endcase
  endfunction
  wire [7:0] v_23807;
  function [7:0] mux_23807(input [0:0] sel);
    case (sel) 0: mux_23807 = 8'h0; 1: mux_23807 = v_23808;
    endcase
  endfunction
  reg [7:0] v_23808 = 8'h0;
  wire [7:0] v_23809;
  wire [7:0] v_23810;
  function [7:0] mux_23810(input [0:0] sel);
    case (sel) 0: mux_23810 = 8'h0; 1: mux_23810 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23811;
  wire [7:0] v_23812;
  wire [7:0] v_23813;
  function [7:0] mux_23813(input [0:0] sel);
    case (sel) 0: mux_23813 = 8'h0; 1: mux_23813 = v_23814;
    endcase
  endfunction
  reg [7:0] v_23814 = 8'h0;
  wire [7:0] v_23815;
  wire [7:0] v_23816;
  function [7:0] mux_23816(input [0:0] sel);
    case (sel) 0: mux_23816 = 8'h0; 1: mux_23816 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23817;
  wire [7:0] v_23818;
  wire [7:0] v_23819;
  function [7:0] mux_23819(input [0:0] sel);
    case (sel) 0: mux_23819 = 8'h0; 1: mux_23819 = v_23820;
    endcase
  endfunction
  reg [7:0] v_23820 = 8'h0;
  wire [7:0] v_23821;
  wire [7:0] v_23822;
  function [7:0] mux_23822(input [0:0] sel);
    case (sel) 0: mux_23822 = 8'h0; 1: mux_23822 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23823;
  wire [7:0] v_23824;
  wire [7:0] v_23825;
  function [7:0] mux_23825(input [0:0] sel);
    case (sel) 0: mux_23825 = 8'h0; 1: mux_23825 = vout_peek_16635;
    endcase
  endfunction
  wire [7:0] v_23826;
  function [7:0] mux_23826(input [0:0] sel);
    case (sel) 0: mux_23826 = 8'h0; 1: mux_23826 = vout_peek_16626;
    endcase
  endfunction
  wire [7:0] v_23827;
  function [7:0] mux_23827(input [0:0] sel);
    case (sel) 0: mux_23827 = 8'h0; 1: mux_23827 = v_23828;
    endcase
  endfunction
  reg [7:0] v_23828 = 8'h0;
  wire [7:0] v_23829;
  wire [7:0] v_23830;
  function [7:0] mux_23830(input [0:0] sel);
    case (sel) 0: mux_23830 = 8'h0; 1: mux_23830 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23831;
  wire [7:0] v_23832;
  wire [7:0] v_23833;
  function [7:0] mux_23833(input [0:0] sel);
    case (sel) 0: mux_23833 = 8'h0; 1: mux_23833 = vout_peek_16598;
    endcase
  endfunction
  wire [7:0] v_23834;
  function [7:0] mux_23834(input [0:0] sel);
    case (sel) 0: mux_23834 = 8'h0; 1: mux_23834 = vout_peek_16589;
    endcase
  endfunction
  wire [7:0] v_23835;
  function [7:0] mux_23835(input [0:0] sel);
    case (sel) 0: mux_23835 = 8'h0; 1: mux_23835 = v_23836;
    endcase
  endfunction
  reg [7:0] v_23836 = 8'h0;
  wire [7:0] v_23837;
  wire [7:0] v_23838;
  function [7:0] mux_23838(input [0:0] sel);
    case (sel) 0: mux_23838 = 8'h0; 1: mux_23838 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23839;
  wire [7:0] v_23840;
  wire [7:0] v_23841;
  function [7:0] mux_23841(input [0:0] sel);
    case (sel) 0: mux_23841 = 8'h0; 1: mux_23841 = v_23842;
    endcase
  endfunction
  reg [7:0] v_23842 = 8'h0;
  wire [7:0] v_23843;
  wire [7:0] v_23844;
  function [7:0] mux_23844(input [0:0] sel);
    case (sel) 0: mux_23844 = 8'h0; 1: mux_23844 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23845;
  wire [7:0] v_23846;
  wire [7:0] v_23847;
  function [7:0] mux_23847(input [0:0] sel);
    case (sel) 0: mux_23847 = 8'h0; 1: mux_23847 = vout_peek_16542;
    endcase
  endfunction
  wire [7:0] v_23848;
  function [7:0] mux_23848(input [0:0] sel);
    case (sel) 0: mux_23848 = 8'h0; 1: mux_23848 = vout_peek_16533;
    endcase
  endfunction
  wire [7:0] v_23849;
  function [7:0] mux_23849(input [0:0] sel);
    case (sel) 0: mux_23849 = 8'h0; 1: mux_23849 = v_23850;
    endcase
  endfunction
  reg [7:0] v_23850 = 8'h0;
  wire [7:0] v_23851;
  wire [7:0] v_23852;
  function [7:0] mux_23852(input [0:0] sel);
    case (sel) 0: mux_23852 = 8'h0; 1: mux_23852 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23853;
  wire [7:0] v_23854;
  wire [7:0] v_23855;
  function [7:0] mux_23855(input [0:0] sel);
    case (sel) 0: mux_23855 = 8'h0; 1: mux_23855 = vout_peek_16505;
    endcase
  endfunction
  wire [7:0] v_23856;
  function [7:0] mux_23856(input [0:0] sel);
    case (sel) 0: mux_23856 = 8'h0; 1: mux_23856 = vout_peek_16496;
    endcase
  endfunction
  wire [7:0] v_23857;
  function [7:0] mux_23857(input [0:0] sel);
    case (sel) 0: mux_23857 = 8'h0; 1: mux_23857 = v_23858;
    endcase
  endfunction
  reg [7:0] v_23858 = 8'h0;
  wire [7:0] v_23859;
  wire [7:0] v_23860;
  function [7:0] mux_23860(input [0:0] sel);
    case (sel) 0: mux_23860 = 8'h0; 1: mux_23860 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23861;
  wire [7:0] v_23862;
  wire [7:0] v_23863;
  function [7:0] mux_23863(input [0:0] sel);
    case (sel) 0: mux_23863 = 8'h0; 1: mux_23863 = v_23864;
    endcase
  endfunction
  reg [7:0] v_23864 = 8'h0;
  wire [7:0] v_23865;
  wire [7:0] v_23866;
  function [7:0] mux_23866(input [0:0] sel);
    case (sel) 0: mux_23866 = 8'h0; 1: mux_23866 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23867;
  wire [7:0] v_23868;
  wire [7:0] v_23869;
  function [7:0] mux_23869(input [0:0] sel);
    case (sel) 0: mux_23869 = 8'h0; 1: mux_23869 = v_23870;
    endcase
  endfunction
  reg [7:0] v_23870 = 8'h0;
  wire [7:0] v_23871;
  wire [7:0] v_23872;
  function [7:0] mux_23872(input [0:0] sel);
    case (sel) 0: mux_23872 = 8'h0; 1: mux_23872 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23873;
  wire [7:0] v_23874;
  wire [7:0] v_23875;
  function [7:0] mux_23875(input [0:0] sel);
    case (sel) 0: mux_23875 = 8'h0; 1: mux_23875 = v_23876;
    endcase
  endfunction
  reg [7:0] v_23876 = 8'h0;
  wire [7:0] v_23877;
  wire [7:0] v_23878;
  function [7:0] mux_23878(input [0:0] sel);
    case (sel) 0: mux_23878 = 8'h0; 1: mux_23878 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23879;
  wire [7:0] v_23880;
  wire [7:0] v_23881;
  function [7:0] mux_23881(input [0:0] sel);
    case (sel) 0: mux_23881 = 8'h0; 1: mux_23881 = vout_peek_16411;
    endcase
  endfunction
  wire [7:0] v_23882;
  function [7:0] mux_23882(input [0:0] sel);
    case (sel) 0: mux_23882 = 8'h0; 1: mux_23882 = vout_peek_16402;
    endcase
  endfunction
  wire [7:0] v_23883;
  function [7:0] mux_23883(input [0:0] sel);
    case (sel) 0: mux_23883 = 8'h0; 1: mux_23883 = v_23884;
    endcase
  endfunction
  reg [7:0] v_23884 = 8'h0;
  wire [7:0] v_23885;
  wire [7:0] v_23886;
  function [7:0] mux_23886(input [0:0] sel);
    case (sel) 0: mux_23886 = 8'h0; 1: mux_23886 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23887;
  wire [7:0] v_23888;
  wire [7:0] v_23889;
  function [7:0] mux_23889(input [0:0] sel);
    case (sel) 0: mux_23889 = 8'h0; 1: mux_23889 = vout_peek_16374;
    endcase
  endfunction
  wire [7:0] v_23890;
  function [7:0] mux_23890(input [0:0] sel);
    case (sel) 0: mux_23890 = 8'h0; 1: mux_23890 = vout_peek_16365;
    endcase
  endfunction
  wire [7:0] v_23891;
  function [7:0] mux_23891(input [0:0] sel);
    case (sel) 0: mux_23891 = 8'h0; 1: mux_23891 = v_23892;
    endcase
  endfunction
  reg [7:0] v_23892 = 8'h0;
  wire [7:0] v_23893;
  wire [7:0] v_23894;
  function [7:0] mux_23894(input [0:0] sel);
    case (sel) 0: mux_23894 = 8'h0; 1: mux_23894 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23895;
  wire [7:0] v_23896;
  wire [7:0] v_23897;
  function [7:0] mux_23897(input [0:0] sel);
    case (sel) 0: mux_23897 = 8'h0; 1: mux_23897 = v_23898;
    endcase
  endfunction
  reg [7:0] v_23898 = 8'h0;
  wire [7:0] v_23899;
  wire [7:0] v_23900;
  function [7:0] mux_23900(input [0:0] sel);
    case (sel) 0: mux_23900 = 8'h0; 1: mux_23900 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23901;
  wire [7:0] v_23902;
  wire [7:0] v_23903;
  function [7:0] mux_23903(input [0:0] sel);
    case (sel) 0: mux_23903 = 8'h0; 1: mux_23903 = vout_peek_16318;
    endcase
  endfunction
  wire [7:0] v_23904;
  function [7:0] mux_23904(input [0:0] sel);
    case (sel) 0: mux_23904 = 8'h0; 1: mux_23904 = vout_peek_16309;
    endcase
  endfunction
  wire [7:0] v_23905;
  function [7:0] mux_23905(input [0:0] sel);
    case (sel) 0: mux_23905 = 8'h0; 1: mux_23905 = v_23906;
    endcase
  endfunction
  reg [7:0] v_23906 = 8'h0;
  wire [7:0] v_23907;
  wire [7:0] v_23908;
  function [7:0] mux_23908(input [0:0] sel);
    case (sel) 0: mux_23908 = 8'h0; 1: mux_23908 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23909;
  wire [7:0] v_23910;
  wire [7:0] v_23911;
  function [7:0] mux_23911(input [0:0] sel);
    case (sel) 0: mux_23911 = 8'h0; 1: mux_23911 = vout_peek_16281;
    endcase
  endfunction
  wire [7:0] v_23912;
  function [7:0] mux_23912(input [0:0] sel);
    case (sel) 0: mux_23912 = 8'h0; 1: mux_23912 = vout_peek_16272;
    endcase
  endfunction
  wire [7:0] v_23913;
  function [7:0] mux_23913(input [0:0] sel);
    case (sel) 0: mux_23913 = 8'h0; 1: mux_23913 = v_23914;
    endcase
  endfunction
  reg [7:0] v_23914 = 8'h0;
  wire [7:0] v_23915;
  wire [7:0] v_23916;
  function [7:0] mux_23916(input [0:0] sel);
    case (sel) 0: mux_23916 = 8'h0; 1: mux_23916 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23917;
  wire [7:0] v_23918;
  wire [7:0] v_23919;
  function [7:0] mux_23919(input [0:0] sel);
    case (sel) 0: mux_23919 = 8'h0; 1: mux_23919 = v_23920;
    endcase
  endfunction
  reg [7:0] v_23920 = 8'h0;
  wire [7:0] v_23921;
  wire [7:0] v_23922;
  function [7:0] mux_23922(input [0:0] sel);
    case (sel) 0: mux_23922 = 8'h0; 1: mux_23922 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23923;
  wire [7:0] v_23924;
  wire [7:0] v_23925;
  function [7:0] mux_23925(input [0:0] sel);
    case (sel) 0: mux_23925 = 8'h0; 1: mux_23925 = v_23926;
    endcase
  endfunction
  reg [7:0] v_23926 = 8'h0;
  wire [7:0] v_23927;
  wire [7:0] v_23928;
  function [7:0] mux_23928(input [0:0] sel);
    case (sel) 0: mux_23928 = 8'h0; 1: mux_23928 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23929;
  wire [7:0] v_23930;
  wire [7:0] v_23931;
  function [7:0] mux_23931(input [0:0] sel);
    case (sel) 0: mux_23931 = 8'h0; 1: mux_23931 = vout_peek_16206;
    endcase
  endfunction
  wire [7:0] v_23932;
  function [7:0] mux_23932(input [0:0] sel);
    case (sel) 0: mux_23932 = 8'h0; 1: mux_23932 = vout_peek_16197;
    endcase
  endfunction
  wire [7:0] v_23933;
  function [7:0] mux_23933(input [0:0] sel);
    case (sel) 0: mux_23933 = 8'h0; 1: mux_23933 = v_23934;
    endcase
  endfunction
  reg [7:0] v_23934 = 8'h0;
  wire [7:0] v_23935;
  wire [7:0] v_23936;
  function [7:0] mux_23936(input [0:0] sel);
    case (sel) 0: mux_23936 = 8'h0; 1: mux_23936 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23937;
  wire [7:0] v_23938;
  wire [7:0] v_23939;
  function [7:0] mux_23939(input [0:0] sel);
    case (sel) 0: mux_23939 = 8'h0; 1: mux_23939 = vout_peek_16169;
    endcase
  endfunction
  wire [7:0] v_23940;
  function [7:0] mux_23940(input [0:0] sel);
    case (sel) 0: mux_23940 = 8'h0; 1: mux_23940 = vout_peek_16160;
    endcase
  endfunction
  wire [7:0] v_23941;
  function [7:0] mux_23941(input [0:0] sel);
    case (sel) 0: mux_23941 = 8'h0; 1: mux_23941 = v_23942;
    endcase
  endfunction
  reg [7:0] v_23942 = 8'h0;
  wire [7:0] v_23943;
  wire [7:0] v_23944;
  function [7:0] mux_23944(input [0:0] sel);
    case (sel) 0: mux_23944 = 8'h0; 1: mux_23944 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23945;
  wire [7:0] v_23946;
  wire [7:0] v_23947;
  function [7:0] mux_23947(input [0:0] sel);
    case (sel) 0: mux_23947 = 8'h0; 1: mux_23947 = v_23948;
    endcase
  endfunction
  reg [7:0] v_23948 = 8'h0;
  wire [7:0] v_23949;
  wire [7:0] v_23950;
  function [7:0] mux_23950(input [0:0] sel);
    case (sel) 0: mux_23950 = 8'h0; 1: mux_23950 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23951;
  wire [7:0] v_23952;
  wire [7:0] v_23953;
  function [7:0] mux_23953(input [0:0] sel);
    case (sel) 0: mux_23953 = 8'h0; 1: mux_23953 = vout_peek_16113;
    endcase
  endfunction
  wire [7:0] v_23954;
  function [7:0] mux_23954(input [0:0] sel);
    case (sel) 0: mux_23954 = 8'h0; 1: mux_23954 = vout_peek_16104;
    endcase
  endfunction
  wire [7:0] v_23955;
  function [7:0] mux_23955(input [0:0] sel);
    case (sel) 0: mux_23955 = 8'h0; 1: mux_23955 = v_23956;
    endcase
  endfunction
  reg [7:0] v_23956 = 8'h0;
  wire [7:0] v_23957;
  wire [7:0] v_23958;
  function [7:0] mux_23958(input [0:0] sel);
    case (sel) 0: mux_23958 = 8'h0; 1: mux_23958 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23959;
  wire [7:0] v_23960;
  wire [7:0] v_23961;
  function [7:0] mux_23961(input [0:0] sel);
    case (sel) 0: mux_23961 = 8'h0; 1: mux_23961 = vout_peek_16076;
    endcase
  endfunction
  wire [7:0] v_23962;
  function [7:0] mux_23962(input [0:0] sel);
    case (sel) 0: mux_23962 = 8'h0; 1: mux_23962 = vout_peek_16067;
    endcase
  endfunction
  wire [7:0] v_23963;
  function [7:0] mux_23963(input [0:0] sel);
    case (sel) 0: mux_23963 = 8'h0; 1: mux_23963 = v_23964;
    endcase
  endfunction
  reg [7:0] v_23964 = 8'h0;
  wire [7:0] v_23965;
  wire [7:0] v_23966;
  function [7:0] mux_23966(input [0:0] sel);
    case (sel) 0: mux_23966 = 8'h0; 1: mux_23966 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23967;
  wire [7:0] v_23968;
  wire [7:0] v_23969;
  function [7:0] mux_23969(input [0:0] sel);
    case (sel) 0: mux_23969 = 8'h0; 1: mux_23969 = v_23970;
    endcase
  endfunction
  reg [7:0] v_23970 = 8'h0;
  wire [7:0] v_23971;
  wire [7:0] v_23972;
  function [7:0] mux_23972(input [0:0] sel);
    case (sel) 0: mux_23972 = 8'h0; 1: mux_23972 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23973;
  wire [7:0] v_23974;
  wire [7:0] v_23975;
  function [7:0] mux_23975(input [0:0] sel);
    case (sel) 0: mux_23975 = 8'h0; 1: mux_23975 = v_23976;
    endcase
  endfunction
  reg [7:0] v_23976 = 8'h0;
  wire [7:0] v_23977;
  wire [7:0] v_23978;
  function [7:0] mux_23978(input [0:0] sel);
    case (sel) 0: mux_23978 = 8'h0; 1: mux_23978 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23979;
  wire [7:0] v_23980;
  wire [7:0] v_23981;
  function [7:0] mux_23981(input [0:0] sel);
    case (sel) 0: mux_23981 = 8'h0; 1: mux_23981 = v_23982;
    endcase
  endfunction
  reg [7:0] v_23982 = 8'h0;
  wire [7:0] v_23983;
  wire [7:0] v_23984;
  function [7:0] mux_23984(input [0:0] sel);
    case (sel) 0: mux_23984 = 8'h0; 1: mux_23984 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23985;
  wire [7:0] v_23986;
  wire [7:0] v_23987;
  function [7:0] mux_23987(input [0:0] sel);
    case (sel) 0: mux_23987 = 8'h0; 1: mux_23987 = v_23988;
    endcase
  endfunction
  reg [7:0] v_23988 = 8'h0;
  wire [7:0] v_23989;
  wire [7:0] v_23990;
  function [7:0] mux_23990(input [0:0] sel);
    case (sel) 0: mux_23990 = 8'h0; 1: mux_23990 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23991;
  wire [7:0] v_23992;
  wire [7:0] v_23993;
  function [7:0] mux_23993(input [0:0] sel);
    case (sel) 0: mux_23993 = 8'h0; 1: mux_23993 = vout_peek_15963;
    endcase
  endfunction
  wire [7:0] v_23994;
  function [7:0] mux_23994(input [0:0] sel);
    case (sel) 0: mux_23994 = 8'h0; 1: mux_23994 = vout_peek_15954;
    endcase
  endfunction
  wire [7:0] v_23995;
  function [7:0] mux_23995(input [0:0] sel);
    case (sel) 0: mux_23995 = 8'h0; 1: mux_23995 = v_23996;
    endcase
  endfunction
  reg [7:0] v_23996 = 8'h0;
  wire [7:0] v_23997;
  wire [7:0] v_23998;
  function [7:0] mux_23998(input [0:0] sel);
    case (sel) 0: mux_23998 = 8'h0; 1: mux_23998 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_23999;
  wire [7:0] v_24000;
  wire [7:0] v_24001;
  function [7:0] mux_24001(input [0:0] sel);
    case (sel) 0: mux_24001 = 8'h0; 1: mux_24001 = vout_peek_15926;
    endcase
  endfunction
  wire [7:0] v_24002;
  function [7:0] mux_24002(input [0:0] sel);
    case (sel) 0: mux_24002 = 8'h0; 1: mux_24002 = vout_peek_15917;
    endcase
  endfunction
  wire [7:0] v_24003;
  function [7:0] mux_24003(input [0:0] sel);
    case (sel) 0: mux_24003 = 8'h0; 1: mux_24003 = v_24004;
    endcase
  endfunction
  reg [7:0] v_24004 = 8'h0;
  wire [7:0] v_24005;
  wire [7:0] v_24006;
  function [7:0] mux_24006(input [0:0] sel);
    case (sel) 0: mux_24006 = 8'h0; 1: mux_24006 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24007;
  wire [7:0] v_24008;
  wire [7:0] v_24009;
  function [7:0] mux_24009(input [0:0] sel);
    case (sel) 0: mux_24009 = 8'h0; 1: mux_24009 = v_24010;
    endcase
  endfunction
  reg [7:0] v_24010 = 8'h0;
  wire [7:0] v_24011;
  wire [7:0] v_24012;
  function [7:0] mux_24012(input [0:0] sel);
    case (sel) 0: mux_24012 = 8'h0; 1: mux_24012 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24013;
  wire [7:0] v_24014;
  wire [7:0] v_24015;
  function [7:0] mux_24015(input [0:0] sel);
    case (sel) 0: mux_24015 = 8'h0; 1: mux_24015 = vout_peek_15870;
    endcase
  endfunction
  wire [7:0] v_24016;
  function [7:0] mux_24016(input [0:0] sel);
    case (sel) 0: mux_24016 = 8'h0; 1: mux_24016 = vout_peek_15861;
    endcase
  endfunction
  wire [7:0] v_24017;
  function [7:0] mux_24017(input [0:0] sel);
    case (sel) 0: mux_24017 = 8'h0; 1: mux_24017 = v_24018;
    endcase
  endfunction
  reg [7:0] v_24018 = 8'h0;
  wire [7:0] v_24019;
  wire [7:0] v_24020;
  function [7:0] mux_24020(input [0:0] sel);
    case (sel) 0: mux_24020 = 8'h0; 1: mux_24020 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24021;
  wire [7:0] v_24022;
  wire [7:0] v_24023;
  function [7:0] mux_24023(input [0:0] sel);
    case (sel) 0: mux_24023 = 8'h0; 1: mux_24023 = vout_peek_15833;
    endcase
  endfunction
  wire [7:0] v_24024;
  function [7:0] mux_24024(input [0:0] sel);
    case (sel) 0: mux_24024 = 8'h0; 1: mux_24024 = vout_peek_15824;
    endcase
  endfunction
  wire [7:0] v_24025;
  function [7:0] mux_24025(input [0:0] sel);
    case (sel) 0: mux_24025 = 8'h0; 1: mux_24025 = v_24026;
    endcase
  endfunction
  reg [7:0] v_24026 = 8'h0;
  wire [7:0] v_24027;
  wire [7:0] v_24028;
  function [7:0] mux_24028(input [0:0] sel);
    case (sel) 0: mux_24028 = 8'h0; 1: mux_24028 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24029;
  wire [7:0] v_24030;
  wire [7:0] v_24031;
  function [7:0] mux_24031(input [0:0] sel);
    case (sel) 0: mux_24031 = 8'h0; 1: mux_24031 = v_24032;
    endcase
  endfunction
  reg [7:0] v_24032 = 8'h0;
  wire [7:0] v_24033;
  wire [7:0] v_24034;
  function [7:0] mux_24034(input [0:0] sel);
    case (sel) 0: mux_24034 = 8'h0; 1: mux_24034 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24035;
  wire [7:0] v_24036;
  wire [7:0] v_24037;
  function [7:0] mux_24037(input [0:0] sel);
    case (sel) 0: mux_24037 = 8'h0; 1: mux_24037 = v_24038;
    endcase
  endfunction
  reg [7:0] v_24038 = 8'h0;
  wire [7:0] v_24039;
  wire [7:0] v_24040;
  function [7:0] mux_24040(input [0:0] sel);
    case (sel) 0: mux_24040 = 8'h0; 1: mux_24040 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24041;
  wire [7:0] v_24042;
  wire [7:0] v_24043;
  function [7:0] mux_24043(input [0:0] sel);
    case (sel) 0: mux_24043 = 8'h0; 1: mux_24043 = vout_peek_15758;
    endcase
  endfunction
  wire [7:0] v_24044;
  function [7:0] mux_24044(input [0:0] sel);
    case (sel) 0: mux_24044 = 8'h0; 1: mux_24044 = vout_peek_15749;
    endcase
  endfunction
  wire [7:0] v_24045;
  function [7:0] mux_24045(input [0:0] sel);
    case (sel) 0: mux_24045 = 8'h0; 1: mux_24045 = v_24046;
    endcase
  endfunction
  reg [7:0] v_24046 = 8'h0;
  wire [7:0] v_24047;
  wire [7:0] v_24048;
  function [7:0] mux_24048(input [0:0] sel);
    case (sel) 0: mux_24048 = 8'h0; 1: mux_24048 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24049;
  wire [7:0] v_24050;
  wire [7:0] v_24051;
  function [7:0] mux_24051(input [0:0] sel);
    case (sel) 0: mux_24051 = 8'h0; 1: mux_24051 = vout_peek_15721;
    endcase
  endfunction
  wire [7:0] v_24052;
  function [7:0] mux_24052(input [0:0] sel);
    case (sel) 0: mux_24052 = 8'h0; 1: mux_24052 = vout_peek_15712;
    endcase
  endfunction
  wire [7:0] v_24053;
  function [7:0] mux_24053(input [0:0] sel);
    case (sel) 0: mux_24053 = 8'h0; 1: mux_24053 = v_24054;
    endcase
  endfunction
  reg [7:0] v_24054 = 8'h0;
  wire [7:0] v_24055;
  wire [7:0] v_24056;
  function [7:0] mux_24056(input [0:0] sel);
    case (sel) 0: mux_24056 = 8'h0; 1: mux_24056 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24057;
  wire [7:0] v_24058;
  wire [7:0] v_24059;
  function [7:0] mux_24059(input [0:0] sel);
    case (sel) 0: mux_24059 = 8'h0; 1: mux_24059 = v_24060;
    endcase
  endfunction
  reg [7:0] v_24060 = 8'h0;
  wire [7:0] v_24061;
  wire [7:0] v_24062;
  function [7:0] mux_24062(input [0:0] sel);
    case (sel) 0: mux_24062 = 8'h0; 1: mux_24062 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24063;
  wire [7:0] v_24064;
  wire [7:0] v_24065;
  function [7:0] mux_24065(input [0:0] sel);
    case (sel) 0: mux_24065 = 8'h0; 1: mux_24065 = vout_peek_15665;
    endcase
  endfunction
  wire [7:0] v_24066;
  function [7:0] mux_24066(input [0:0] sel);
    case (sel) 0: mux_24066 = 8'h0; 1: mux_24066 = vout_peek_15656;
    endcase
  endfunction
  wire [7:0] v_24067;
  function [7:0] mux_24067(input [0:0] sel);
    case (sel) 0: mux_24067 = 8'h0; 1: mux_24067 = v_24068;
    endcase
  endfunction
  reg [7:0] v_24068 = 8'h0;
  wire [7:0] v_24069;
  wire [7:0] v_24070;
  function [7:0] mux_24070(input [0:0] sel);
    case (sel) 0: mux_24070 = 8'h0; 1: mux_24070 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24071;
  wire [7:0] v_24072;
  wire [7:0] v_24073;
  function [7:0] mux_24073(input [0:0] sel);
    case (sel) 0: mux_24073 = 8'h0; 1: mux_24073 = vout_peek_15628;
    endcase
  endfunction
  wire [7:0] v_24074;
  function [7:0] mux_24074(input [0:0] sel);
    case (sel) 0: mux_24074 = 8'h0; 1: mux_24074 = vout_peek_15619;
    endcase
  endfunction
  wire [7:0] v_24075;
  function [7:0] mux_24075(input [0:0] sel);
    case (sel) 0: mux_24075 = 8'h0; 1: mux_24075 = v_24076;
    endcase
  endfunction
  reg [7:0] v_24076 = 8'h0;
  wire [7:0] v_24077;
  wire [7:0] v_24078;
  function [7:0] mux_24078(input [0:0] sel);
    case (sel) 0: mux_24078 = 8'h0; 1: mux_24078 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24079;
  wire [7:0] v_24080;
  wire [7:0] v_24081;
  function [7:0] mux_24081(input [0:0] sel);
    case (sel) 0: mux_24081 = 8'h0; 1: mux_24081 = v_24082;
    endcase
  endfunction
  reg [7:0] v_24082 = 8'h0;
  wire [7:0] v_24083;
  wire [7:0] v_24084;
  function [7:0] mux_24084(input [0:0] sel);
    case (sel) 0: mux_24084 = 8'h0; 1: mux_24084 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24085;
  wire [7:0] v_24086;
  wire [7:0] v_24087;
  function [7:0] mux_24087(input [0:0] sel);
    case (sel) 0: mux_24087 = 8'h0; 1: mux_24087 = v_24088;
    endcase
  endfunction
  reg [7:0] v_24088 = 8'h0;
  wire [7:0] v_24089;
  wire [7:0] v_24090;
  function [7:0] mux_24090(input [0:0] sel);
    case (sel) 0: mux_24090 = 8'h0; 1: mux_24090 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24091;
  wire [7:0] v_24092;
  wire [7:0] v_24093;
  function [7:0] mux_24093(input [0:0] sel);
    case (sel) 0: mux_24093 = 8'h0; 1: mux_24093 = v_24094;
    endcase
  endfunction
  reg [7:0] v_24094 = 8'h0;
  wire [7:0] v_24095;
  wire [7:0] v_24096;
  function [7:0] mux_24096(input [0:0] sel);
    case (sel) 0: mux_24096 = 8'h0; 1: mux_24096 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24097;
  wire [7:0] v_24098;
  wire [7:0] v_24099;
  function [7:0] mux_24099(input [0:0] sel);
    case (sel) 0: mux_24099 = 8'h0; 1: mux_24099 = vout_peek_15534;
    endcase
  endfunction
  wire [7:0] v_24100;
  function [7:0] mux_24100(input [0:0] sel);
    case (sel) 0: mux_24100 = 8'h0; 1: mux_24100 = vout_peek_15525;
    endcase
  endfunction
  wire [7:0] v_24101;
  function [7:0] mux_24101(input [0:0] sel);
    case (sel) 0: mux_24101 = 8'h0; 1: mux_24101 = v_24102;
    endcase
  endfunction
  reg [7:0] v_24102 = 8'h0;
  wire [7:0] v_24103;
  wire [7:0] v_24104;
  function [7:0] mux_24104(input [0:0] sel);
    case (sel) 0: mux_24104 = 8'h0; 1: mux_24104 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24105;
  wire [7:0] v_24106;
  wire [7:0] v_24107;
  function [7:0] mux_24107(input [0:0] sel);
    case (sel) 0: mux_24107 = 8'h0; 1: mux_24107 = vout_peek_15497;
    endcase
  endfunction
  wire [7:0] v_24108;
  function [7:0] mux_24108(input [0:0] sel);
    case (sel) 0: mux_24108 = 8'h0; 1: mux_24108 = vout_peek_15488;
    endcase
  endfunction
  wire [7:0] v_24109;
  function [7:0] mux_24109(input [0:0] sel);
    case (sel) 0: mux_24109 = 8'h0; 1: mux_24109 = v_24110;
    endcase
  endfunction
  reg [7:0] v_24110 = 8'h0;
  wire [7:0] v_24111;
  wire [7:0] v_24112;
  function [7:0] mux_24112(input [0:0] sel);
    case (sel) 0: mux_24112 = 8'h0; 1: mux_24112 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24113;
  wire [7:0] v_24114;
  wire [7:0] v_24115;
  function [7:0] mux_24115(input [0:0] sel);
    case (sel) 0: mux_24115 = 8'h0; 1: mux_24115 = v_24116;
    endcase
  endfunction
  reg [7:0] v_24116 = 8'h0;
  wire [7:0] v_24117;
  wire [7:0] v_24118;
  function [7:0] mux_24118(input [0:0] sel);
    case (sel) 0: mux_24118 = 8'h0; 1: mux_24118 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24119;
  wire [7:0] v_24120;
  wire [7:0] v_24121;
  function [7:0] mux_24121(input [0:0] sel);
    case (sel) 0: mux_24121 = 8'h0; 1: mux_24121 = vout_peek_15441;
    endcase
  endfunction
  wire [7:0] v_24122;
  function [7:0] mux_24122(input [0:0] sel);
    case (sel) 0: mux_24122 = 8'h0; 1: mux_24122 = vout_peek_15432;
    endcase
  endfunction
  wire [7:0] v_24123;
  function [7:0] mux_24123(input [0:0] sel);
    case (sel) 0: mux_24123 = 8'h0; 1: mux_24123 = v_24124;
    endcase
  endfunction
  reg [7:0] v_24124 = 8'h0;
  wire [7:0] v_24125;
  wire [7:0] v_24126;
  function [7:0] mux_24126(input [0:0] sel);
    case (sel) 0: mux_24126 = 8'h0; 1: mux_24126 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24127;
  wire [7:0] v_24128;
  wire [7:0] v_24129;
  function [7:0] mux_24129(input [0:0] sel);
    case (sel) 0: mux_24129 = 8'h0; 1: mux_24129 = vout_peek_15404;
    endcase
  endfunction
  wire [7:0] v_24130;
  function [7:0] mux_24130(input [0:0] sel);
    case (sel) 0: mux_24130 = 8'h0; 1: mux_24130 = vout_peek_15395;
    endcase
  endfunction
  wire [7:0] v_24131;
  function [7:0] mux_24131(input [0:0] sel);
    case (sel) 0: mux_24131 = 8'h0; 1: mux_24131 = v_24132;
    endcase
  endfunction
  reg [7:0] v_24132 = 8'h0;
  wire [7:0] v_24133;
  wire [7:0] v_24134;
  function [7:0] mux_24134(input [0:0] sel);
    case (sel) 0: mux_24134 = 8'h0; 1: mux_24134 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24135;
  wire [7:0] v_24136;
  wire [7:0] v_24137;
  function [7:0] mux_24137(input [0:0] sel);
    case (sel) 0: mux_24137 = 8'h0; 1: mux_24137 = v_24138;
    endcase
  endfunction
  reg [7:0] v_24138 = 8'h0;
  wire [7:0] v_24139;
  wire [7:0] v_24140;
  function [7:0] mux_24140(input [0:0] sel);
    case (sel) 0: mux_24140 = 8'h0; 1: mux_24140 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24141;
  wire [7:0] v_24142;
  wire [7:0] v_24143;
  function [7:0] mux_24143(input [0:0] sel);
    case (sel) 0: mux_24143 = 8'h0; 1: mux_24143 = v_24144;
    endcase
  endfunction
  reg [7:0] v_24144 = 8'h0;
  wire [7:0] v_24145;
  wire [7:0] v_24146;
  function [7:0] mux_24146(input [0:0] sel);
    case (sel) 0: mux_24146 = 8'h0; 1: mux_24146 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24147;
  wire [7:0] v_24148;
  wire [7:0] v_24149;
  function [7:0] mux_24149(input [0:0] sel);
    case (sel) 0: mux_24149 = 8'h0; 1: mux_24149 = vout_peek_15329;
    endcase
  endfunction
  wire [7:0] v_24150;
  function [7:0] mux_24150(input [0:0] sel);
    case (sel) 0: mux_24150 = 8'h0; 1: mux_24150 = vout_peek_15320;
    endcase
  endfunction
  wire [7:0] v_24151;
  function [7:0] mux_24151(input [0:0] sel);
    case (sel) 0: mux_24151 = 8'h0; 1: mux_24151 = v_24152;
    endcase
  endfunction
  reg [7:0] v_24152 = 8'h0;
  wire [7:0] v_24153;
  wire [7:0] v_24154;
  function [7:0] mux_24154(input [0:0] sel);
    case (sel) 0: mux_24154 = 8'h0; 1: mux_24154 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24155;
  wire [7:0] v_24156;
  wire [7:0] v_24157;
  function [7:0] mux_24157(input [0:0] sel);
    case (sel) 0: mux_24157 = 8'h0; 1: mux_24157 = vout_peek_15292;
    endcase
  endfunction
  wire [7:0] v_24158;
  function [7:0] mux_24158(input [0:0] sel);
    case (sel) 0: mux_24158 = 8'h0; 1: mux_24158 = vout_peek_15283;
    endcase
  endfunction
  wire [7:0] v_24159;
  function [7:0] mux_24159(input [0:0] sel);
    case (sel) 0: mux_24159 = 8'h0; 1: mux_24159 = v_24160;
    endcase
  endfunction
  reg [7:0] v_24160 = 8'h0;
  wire [7:0] v_24161;
  wire [7:0] v_24162;
  function [7:0] mux_24162(input [0:0] sel);
    case (sel) 0: mux_24162 = 8'h0; 1: mux_24162 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24163;
  wire [7:0] v_24164;
  wire [7:0] v_24165;
  function [7:0] mux_24165(input [0:0] sel);
    case (sel) 0: mux_24165 = 8'h0; 1: mux_24165 = v_24166;
    endcase
  endfunction
  reg [7:0] v_24166 = 8'h0;
  wire [7:0] v_24167;
  wire [7:0] v_24168;
  function [7:0] mux_24168(input [0:0] sel);
    case (sel) 0: mux_24168 = 8'h0; 1: mux_24168 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24169;
  wire [7:0] v_24170;
  wire [7:0] v_24171;
  function [7:0] mux_24171(input [0:0] sel);
    case (sel) 0: mux_24171 = 8'h0; 1: mux_24171 = vout_peek_15236;
    endcase
  endfunction
  wire [7:0] v_24172;
  function [7:0] mux_24172(input [0:0] sel);
    case (sel) 0: mux_24172 = 8'h0; 1: mux_24172 = vout_peek_15227;
    endcase
  endfunction
  wire [7:0] v_24173;
  function [7:0] mux_24173(input [0:0] sel);
    case (sel) 0: mux_24173 = 8'h0; 1: mux_24173 = v_24174;
    endcase
  endfunction
  reg [7:0] v_24174 = 8'h0;
  wire [7:0] v_24175;
  wire [7:0] v_24176;
  function [7:0] mux_24176(input [0:0] sel);
    case (sel) 0: mux_24176 = 8'h0; 1: mux_24176 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24177;
  wire [7:0] v_24178;
  wire [7:0] v_24179;
  function [7:0] mux_24179(input [0:0] sel);
    case (sel) 0: mux_24179 = 8'h0; 1: mux_24179 = vout_peek_15199;
    endcase
  endfunction
  wire [7:0] v_24180;
  function [7:0] mux_24180(input [0:0] sel);
    case (sel) 0: mux_24180 = 8'h0; 1: mux_24180 = vout_peek_15190;
    endcase
  endfunction
  wire [7:0] v_24181;
  function [7:0] mux_24181(input [0:0] sel);
    case (sel) 0: mux_24181 = 8'h0; 1: mux_24181 = v_24182;
    endcase
  endfunction
  reg [7:0] v_24182 = 8'h0;
  wire [7:0] v_24183;
  wire [7:0] v_24184;
  function [7:0] mux_24184(input [0:0] sel);
    case (sel) 0: mux_24184 = 8'h0; 1: mux_24184 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24185;
  wire [7:0] v_24186;
  wire [7:0] v_24187;
  function [7:0] mux_24187(input [0:0] sel);
    case (sel) 0: mux_24187 = 8'h0; 1: mux_24187 = v_24188;
    endcase
  endfunction
  reg [7:0] v_24188 = 8'h0;
  wire [7:0] v_24189;
  wire [7:0] v_24190;
  function [7:0] mux_24190(input [0:0] sel);
    case (sel) 0: mux_24190 = 8'h0; 1: mux_24190 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24191;
  wire [7:0] v_24192;
  wire [7:0] v_24193;
  function [7:0] mux_24193(input [0:0] sel);
    case (sel) 0: mux_24193 = 8'h0; 1: mux_24193 = v_24194;
    endcase
  endfunction
  reg [7:0] v_24194 = 8'h0;
  wire [7:0] v_24195;
  wire [7:0] v_24196;
  function [7:0] mux_24196(input [0:0] sel);
    case (sel) 0: mux_24196 = 8'h0; 1: mux_24196 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24197;
  wire [7:0] v_24198;
  wire [7:0] v_24199;
  function [7:0] mux_24199(input [0:0] sel);
    case (sel) 0: mux_24199 = 8'h0; 1: mux_24199 = v_24200;
    endcase
  endfunction
  reg [7:0] v_24200 = 8'h0;
  wire [7:0] v_24201;
  wire [7:0] v_24202;
  function [7:0] mux_24202(input [0:0] sel);
    case (sel) 0: mux_24202 = 8'h0; 1: mux_24202 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24203;
  wire [7:0] v_24204;
  wire [7:0] v_24205;
  function [7:0] mux_24205(input [0:0] sel);
    case (sel) 0: mux_24205 = 8'h0; 1: mux_24205 = v_24206;
    endcase
  endfunction
  reg [7:0] v_24206 = 8'h0;
  wire [7:0] v_24207;
  wire [7:0] v_24208;
  function [7:0] mux_24208(input [0:0] sel);
    case (sel) 0: mux_24208 = 8'h0; 1: mux_24208 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24209;
  wire [7:0] v_24210;
  wire [7:0] v_24211;
  function [7:0] mux_24211(input [0:0] sel);
    case (sel) 0: mux_24211 = 8'h0; 1: mux_24211 = v_24212;
    endcase
  endfunction
  reg [7:0] v_24212 = 8'h0;
  wire [7:0] v_24213;
  wire [7:0] v_24214;
  function [7:0] mux_24214(input [0:0] sel);
    case (sel) 0: mux_24214 = 8'h0; 1: mux_24214 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24215;
  wire [7:0] v_24216;
  wire [7:0] v_24217;
  function [7:0] mux_24217(input [0:0] sel);
    case (sel) 0: mux_24217 = 8'h0; 1: mux_24217 = v_24218;
    endcase
  endfunction
  reg [7:0] v_24218 = 8'h0;
  wire [7:0] v_24219;
  wire [7:0] v_24220;
  function [7:0] mux_24220(input [0:0] sel);
    case (sel) 0: mux_24220 = 8'h0; 1: mux_24220 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24221;
  wire [7:0] v_24222;
  wire [7:0] v_24223;
  function [7:0] mux_24223(input [0:0] sel);
    case (sel) 0: mux_24223 = 8'h0; 1: mux_24223 = v_24224;
    endcase
  endfunction
  reg [7:0] v_24224 = 8'h0;
  wire [7:0] v_24225;
  wire [7:0] v_24226;
  function [7:0] mux_24226(input [0:0] sel);
    case (sel) 0: mux_24226 = 8'h0; 1: mux_24226 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24227;
  wire [7:0] v_24228;
  wire [7:0] v_24229;
  function [7:0] mux_24229(input [0:0] sel);
    case (sel) 0: mux_24229 = 8'h0; 1: mux_24229 = vout_peek_15029;
    endcase
  endfunction
  wire [7:0] v_24230;
  function [7:0] mux_24230(input [0:0] sel);
    case (sel) 0: mux_24230 = 8'h0; 1: mux_24230 = vout_peek_15020;
    endcase
  endfunction
  wire [7:0] v_24231;
  function [7:0] mux_24231(input [0:0] sel);
    case (sel) 0: mux_24231 = 8'h0; 1: mux_24231 = v_24232;
    endcase
  endfunction
  reg [7:0] v_24232 = 8'h0;
  wire [7:0] v_24233;
  wire [7:0] v_24234;
  function [7:0] mux_24234(input [0:0] sel);
    case (sel) 0: mux_24234 = 8'h0; 1: mux_24234 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24235;
  wire [7:0] v_24236;
  wire [7:0] v_24237;
  function [7:0] mux_24237(input [0:0] sel);
    case (sel) 0: mux_24237 = 8'h0; 1: mux_24237 = vout_peek_14992;
    endcase
  endfunction
  wire [7:0] v_24238;
  function [7:0] mux_24238(input [0:0] sel);
    case (sel) 0: mux_24238 = 8'h0; 1: mux_24238 = vout_peek_14983;
    endcase
  endfunction
  wire [7:0] v_24239;
  function [7:0] mux_24239(input [0:0] sel);
    case (sel) 0: mux_24239 = 8'h0; 1: mux_24239 = v_24240;
    endcase
  endfunction
  reg [7:0] v_24240 = 8'h0;
  wire [7:0] v_24241;
  wire [7:0] v_24242;
  function [7:0] mux_24242(input [0:0] sel);
    case (sel) 0: mux_24242 = 8'h0; 1: mux_24242 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24243;
  wire [7:0] v_24244;
  wire [7:0] v_24245;
  function [7:0] mux_24245(input [0:0] sel);
    case (sel) 0: mux_24245 = 8'h0; 1: mux_24245 = v_24246;
    endcase
  endfunction
  reg [7:0] v_24246 = 8'h0;
  wire [7:0] v_24247;
  wire [7:0] v_24248;
  function [7:0] mux_24248(input [0:0] sel);
    case (sel) 0: mux_24248 = 8'h0; 1: mux_24248 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24249;
  wire [7:0] v_24250;
  wire [7:0] v_24251;
  function [7:0] mux_24251(input [0:0] sel);
    case (sel) 0: mux_24251 = 8'h0; 1: mux_24251 = vout_peek_14936;
    endcase
  endfunction
  wire [7:0] v_24252;
  function [7:0] mux_24252(input [0:0] sel);
    case (sel) 0: mux_24252 = 8'h0; 1: mux_24252 = vout_peek_14927;
    endcase
  endfunction
  wire [7:0] v_24253;
  function [7:0] mux_24253(input [0:0] sel);
    case (sel) 0: mux_24253 = 8'h0; 1: mux_24253 = v_24254;
    endcase
  endfunction
  reg [7:0] v_24254 = 8'h0;
  wire [7:0] v_24255;
  wire [7:0] v_24256;
  function [7:0] mux_24256(input [0:0] sel);
    case (sel) 0: mux_24256 = 8'h0; 1: mux_24256 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24257;
  wire [7:0] v_24258;
  wire [7:0] v_24259;
  function [7:0] mux_24259(input [0:0] sel);
    case (sel) 0: mux_24259 = 8'h0; 1: mux_24259 = vout_peek_14899;
    endcase
  endfunction
  wire [7:0] v_24260;
  function [7:0] mux_24260(input [0:0] sel);
    case (sel) 0: mux_24260 = 8'h0; 1: mux_24260 = vout_peek_14890;
    endcase
  endfunction
  wire [7:0] v_24261;
  function [7:0] mux_24261(input [0:0] sel);
    case (sel) 0: mux_24261 = 8'h0; 1: mux_24261 = v_24262;
    endcase
  endfunction
  reg [7:0] v_24262 = 8'h0;
  wire [7:0] v_24263;
  wire [7:0] v_24264;
  function [7:0] mux_24264(input [0:0] sel);
    case (sel) 0: mux_24264 = 8'h0; 1: mux_24264 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24265;
  wire [7:0] v_24266;
  wire [7:0] v_24267;
  function [7:0] mux_24267(input [0:0] sel);
    case (sel) 0: mux_24267 = 8'h0; 1: mux_24267 = v_24268;
    endcase
  endfunction
  reg [7:0] v_24268 = 8'h0;
  wire [7:0] v_24269;
  wire [7:0] v_24270;
  function [7:0] mux_24270(input [0:0] sel);
    case (sel) 0: mux_24270 = 8'h0; 1: mux_24270 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24271;
  wire [7:0] v_24272;
  wire [7:0] v_24273;
  function [7:0] mux_24273(input [0:0] sel);
    case (sel) 0: mux_24273 = 8'h0; 1: mux_24273 = v_24274;
    endcase
  endfunction
  reg [7:0] v_24274 = 8'h0;
  wire [7:0] v_24275;
  wire [7:0] v_24276;
  function [7:0] mux_24276(input [0:0] sel);
    case (sel) 0: mux_24276 = 8'h0; 1: mux_24276 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24277;
  wire [7:0] v_24278;
  wire [7:0] v_24279;
  function [7:0] mux_24279(input [0:0] sel);
    case (sel) 0: mux_24279 = 8'h0; 1: mux_24279 = vout_peek_14824;
    endcase
  endfunction
  wire [7:0] v_24280;
  function [7:0] mux_24280(input [0:0] sel);
    case (sel) 0: mux_24280 = 8'h0; 1: mux_24280 = vout_peek_14815;
    endcase
  endfunction
  wire [7:0] v_24281;
  function [7:0] mux_24281(input [0:0] sel);
    case (sel) 0: mux_24281 = 8'h0; 1: mux_24281 = v_24282;
    endcase
  endfunction
  reg [7:0] v_24282 = 8'h0;
  wire [7:0] v_24283;
  wire [7:0] v_24284;
  function [7:0] mux_24284(input [0:0] sel);
    case (sel) 0: mux_24284 = 8'h0; 1: mux_24284 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24285;
  wire [7:0] v_24286;
  wire [7:0] v_24287;
  function [7:0] mux_24287(input [0:0] sel);
    case (sel) 0: mux_24287 = 8'h0; 1: mux_24287 = vout_peek_14787;
    endcase
  endfunction
  wire [7:0] v_24288;
  function [7:0] mux_24288(input [0:0] sel);
    case (sel) 0: mux_24288 = 8'h0; 1: mux_24288 = vout_peek_14778;
    endcase
  endfunction
  wire [7:0] v_24289;
  function [7:0] mux_24289(input [0:0] sel);
    case (sel) 0: mux_24289 = 8'h0; 1: mux_24289 = v_24290;
    endcase
  endfunction
  reg [7:0] v_24290 = 8'h0;
  wire [7:0] v_24291;
  wire [7:0] v_24292;
  function [7:0] mux_24292(input [0:0] sel);
    case (sel) 0: mux_24292 = 8'h0; 1: mux_24292 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24293;
  wire [7:0] v_24294;
  wire [7:0] v_24295;
  function [7:0] mux_24295(input [0:0] sel);
    case (sel) 0: mux_24295 = 8'h0; 1: mux_24295 = v_24296;
    endcase
  endfunction
  reg [7:0] v_24296 = 8'h0;
  wire [7:0] v_24297;
  wire [7:0] v_24298;
  function [7:0] mux_24298(input [0:0] sel);
    case (sel) 0: mux_24298 = 8'h0; 1: mux_24298 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24299;
  wire [7:0] v_24300;
  wire [7:0] v_24301;
  function [7:0] mux_24301(input [0:0] sel);
    case (sel) 0: mux_24301 = 8'h0; 1: mux_24301 = vout_peek_14731;
    endcase
  endfunction
  wire [7:0] v_24302;
  function [7:0] mux_24302(input [0:0] sel);
    case (sel) 0: mux_24302 = 8'h0; 1: mux_24302 = vout_peek_14722;
    endcase
  endfunction
  wire [7:0] v_24303;
  function [7:0] mux_24303(input [0:0] sel);
    case (sel) 0: mux_24303 = 8'h0; 1: mux_24303 = v_24304;
    endcase
  endfunction
  reg [7:0] v_24304 = 8'h0;
  wire [7:0] v_24305;
  wire [7:0] v_24306;
  function [7:0] mux_24306(input [0:0] sel);
    case (sel) 0: mux_24306 = 8'h0; 1: mux_24306 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24307;
  wire [7:0] v_24308;
  wire [7:0] v_24309;
  function [7:0] mux_24309(input [0:0] sel);
    case (sel) 0: mux_24309 = 8'h0; 1: mux_24309 = vout_peek_14694;
    endcase
  endfunction
  wire [7:0] v_24310;
  function [7:0] mux_24310(input [0:0] sel);
    case (sel) 0: mux_24310 = 8'h0; 1: mux_24310 = vout_peek_14685;
    endcase
  endfunction
  wire [7:0] v_24311;
  function [7:0] mux_24311(input [0:0] sel);
    case (sel) 0: mux_24311 = 8'h0; 1: mux_24311 = v_24312;
    endcase
  endfunction
  reg [7:0] v_24312 = 8'h0;
  wire [7:0] v_24313;
  wire [7:0] v_24314;
  function [7:0] mux_24314(input [0:0] sel);
    case (sel) 0: mux_24314 = 8'h0; 1: mux_24314 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24315;
  wire [7:0] v_24316;
  wire [7:0] v_24317;
  function [7:0] mux_24317(input [0:0] sel);
    case (sel) 0: mux_24317 = 8'h0; 1: mux_24317 = v_24318;
    endcase
  endfunction
  reg [7:0] v_24318 = 8'h0;
  wire [7:0] v_24319;
  wire [7:0] v_24320;
  function [7:0] mux_24320(input [0:0] sel);
    case (sel) 0: mux_24320 = 8'h0; 1: mux_24320 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24321;
  wire [7:0] v_24322;
  wire [7:0] v_24323;
  function [7:0] mux_24323(input [0:0] sel);
    case (sel) 0: mux_24323 = 8'h0; 1: mux_24323 = v_24324;
    endcase
  endfunction
  reg [7:0] v_24324 = 8'h0;
  wire [7:0] v_24325;
  wire [7:0] v_24326;
  function [7:0] mux_24326(input [0:0] sel);
    case (sel) 0: mux_24326 = 8'h0; 1: mux_24326 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24327;
  wire [7:0] v_24328;
  wire [7:0] v_24329;
  function [7:0] mux_24329(input [0:0] sel);
    case (sel) 0: mux_24329 = 8'h0; 1: mux_24329 = v_24330;
    endcase
  endfunction
  reg [7:0] v_24330 = 8'h0;
  wire [7:0] v_24331;
  wire [7:0] v_24332;
  function [7:0] mux_24332(input [0:0] sel);
    case (sel) 0: mux_24332 = 8'h0; 1: mux_24332 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24333;
  wire [7:0] v_24334;
  wire [7:0] v_24335;
  function [7:0] mux_24335(input [0:0] sel);
    case (sel) 0: mux_24335 = 8'h0; 1: mux_24335 = vout_peek_14600;
    endcase
  endfunction
  wire [7:0] v_24336;
  function [7:0] mux_24336(input [0:0] sel);
    case (sel) 0: mux_24336 = 8'h0; 1: mux_24336 = vout_peek_14591;
    endcase
  endfunction
  wire [7:0] v_24337;
  function [7:0] mux_24337(input [0:0] sel);
    case (sel) 0: mux_24337 = 8'h0; 1: mux_24337 = v_24338;
    endcase
  endfunction
  reg [7:0] v_24338 = 8'h0;
  wire [7:0] v_24339;
  wire [7:0] v_24340;
  function [7:0] mux_24340(input [0:0] sel);
    case (sel) 0: mux_24340 = 8'h0; 1: mux_24340 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24341;
  wire [7:0] v_24342;
  wire [7:0] v_24343;
  function [7:0] mux_24343(input [0:0] sel);
    case (sel) 0: mux_24343 = 8'h0; 1: mux_24343 = vout_peek_14563;
    endcase
  endfunction
  wire [7:0] v_24344;
  function [7:0] mux_24344(input [0:0] sel);
    case (sel) 0: mux_24344 = 8'h0; 1: mux_24344 = vout_peek_14554;
    endcase
  endfunction
  wire [7:0] v_24345;
  function [7:0] mux_24345(input [0:0] sel);
    case (sel) 0: mux_24345 = 8'h0; 1: mux_24345 = v_24346;
    endcase
  endfunction
  reg [7:0] v_24346 = 8'h0;
  wire [7:0] v_24347;
  wire [7:0] v_24348;
  function [7:0] mux_24348(input [0:0] sel);
    case (sel) 0: mux_24348 = 8'h0; 1: mux_24348 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24349;
  wire [7:0] v_24350;
  wire [7:0] v_24351;
  function [7:0] mux_24351(input [0:0] sel);
    case (sel) 0: mux_24351 = 8'h0; 1: mux_24351 = v_24352;
    endcase
  endfunction
  reg [7:0] v_24352 = 8'h0;
  wire [7:0] v_24353;
  wire [7:0] v_24354;
  function [7:0] mux_24354(input [0:0] sel);
    case (sel) 0: mux_24354 = 8'h0; 1: mux_24354 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24355;
  wire [7:0] v_24356;
  wire [7:0] v_24357;
  function [7:0] mux_24357(input [0:0] sel);
    case (sel) 0: mux_24357 = 8'h0; 1: mux_24357 = vout_peek_14507;
    endcase
  endfunction
  wire [7:0] v_24358;
  function [7:0] mux_24358(input [0:0] sel);
    case (sel) 0: mux_24358 = 8'h0; 1: mux_24358 = vout_peek_14498;
    endcase
  endfunction
  wire [7:0] v_24359;
  function [7:0] mux_24359(input [0:0] sel);
    case (sel) 0: mux_24359 = 8'h0; 1: mux_24359 = v_24360;
    endcase
  endfunction
  reg [7:0] v_24360 = 8'h0;
  wire [7:0] v_24361;
  wire [7:0] v_24362;
  function [7:0] mux_24362(input [0:0] sel);
    case (sel) 0: mux_24362 = 8'h0; 1: mux_24362 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24363;
  wire [7:0] v_24364;
  wire [7:0] v_24365;
  function [7:0] mux_24365(input [0:0] sel);
    case (sel) 0: mux_24365 = 8'h0; 1: mux_24365 = vout_peek_14470;
    endcase
  endfunction
  wire [7:0] v_24366;
  function [7:0] mux_24366(input [0:0] sel);
    case (sel) 0: mux_24366 = 8'h0; 1: mux_24366 = vout_peek_14461;
    endcase
  endfunction
  wire [7:0] v_24367;
  function [7:0] mux_24367(input [0:0] sel);
    case (sel) 0: mux_24367 = 8'h0; 1: mux_24367 = v_24368;
    endcase
  endfunction
  reg [7:0] v_24368 = 8'h0;
  wire [7:0] v_24369;
  wire [7:0] v_24370;
  function [7:0] mux_24370(input [0:0] sel);
    case (sel) 0: mux_24370 = 8'h0; 1: mux_24370 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24371;
  wire [7:0] v_24372;
  wire [7:0] v_24373;
  function [7:0] mux_24373(input [0:0] sel);
    case (sel) 0: mux_24373 = 8'h0; 1: mux_24373 = v_24374;
    endcase
  endfunction
  reg [7:0] v_24374 = 8'h0;
  wire [7:0] v_24375;
  wire [7:0] v_24376;
  function [7:0] mux_24376(input [0:0] sel);
    case (sel) 0: mux_24376 = 8'h0; 1: mux_24376 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24377;
  wire [7:0] v_24378;
  wire [7:0] v_24379;
  function [7:0] mux_24379(input [0:0] sel);
    case (sel) 0: mux_24379 = 8'h0; 1: mux_24379 = v_24380;
    endcase
  endfunction
  reg [7:0] v_24380 = 8'h0;
  wire [7:0] v_24381;
  wire [7:0] v_24382;
  function [7:0] mux_24382(input [0:0] sel);
    case (sel) 0: mux_24382 = 8'h0; 1: mux_24382 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24383;
  wire [7:0] v_24384;
  wire [7:0] v_24385;
  function [7:0] mux_24385(input [0:0] sel);
    case (sel) 0: mux_24385 = 8'h0; 1: mux_24385 = vout_peek_14395;
    endcase
  endfunction
  wire [7:0] v_24386;
  function [7:0] mux_24386(input [0:0] sel);
    case (sel) 0: mux_24386 = 8'h0; 1: mux_24386 = vout_peek_14386;
    endcase
  endfunction
  wire [7:0] v_24387;
  function [7:0] mux_24387(input [0:0] sel);
    case (sel) 0: mux_24387 = 8'h0; 1: mux_24387 = v_24388;
    endcase
  endfunction
  reg [7:0] v_24388 = 8'h0;
  wire [7:0] v_24389;
  wire [7:0] v_24390;
  function [7:0] mux_24390(input [0:0] sel);
    case (sel) 0: mux_24390 = 8'h0; 1: mux_24390 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24391;
  wire [7:0] v_24392;
  wire [7:0] v_24393;
  function [7:0] mux_24393(input [0:0] sel);
    case (sel) 0: mux_24393 = 8'h0; 1: mux_24393 = vout_peek_14358;
    endcase
  endfunction
  wire [7:0] v_24394;
  function [7:0] mux_24394(input [0:0] sel);
    case (sel) 0: mux_24394 = 8'h0; 1: mux_24394 = vout_peek_14349;
    endcase
  endfunction
  wire [7:0] v_24395;
  function [7:0] mux_24395(input [0:0] sel);
    case (sel) 0: mux_24395 = 8'h0; 1: mux_24395 = v_24396;
    endcase
  endfunction
  reg [7:0] v_24396 = 8'h0;
  wire [7:0] v_24397;
  wire [7:0] v_24398;
  function [7:0] mux_24398(input [0:0] sel);
    case (sel) 0: mux_24398 = 8'h0; 1: mux_24398 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24399;
  wire [7:0] v_24400;
  wire [7:0] v_24401;
  function [7:0] mux_24401(input [0:0] sel);
    case (sel) 0: mux_24401 = 8'h0; 1: mux_24401 = v_24402;
    endcase
  endfunction
  reg [7:0] v_24402 = 8'h0;
  wire [7:0] v_24403;
  wire [7:0] v_24404;
  function [7:0] mux_24404(input [0:0] sel);
    case (sel) 0: mux_24404 = 8'h0; 1: mux_24404 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24405;
  wire [7:0] v_24406;
  wire [7:0] v_24407;
  function [7:0] mux_24407(input [0:0] sel);
    case (sel) 0: mux_24407 = 8'h0; 1: mux_24407 = vout_peek_14302;
    endcase
  endfunction
  wire [7:0] v_24408;
  function [7:0] mux_24408(input [0:0] sel);
    case (sel) 0: mux_24408 = 8'h0; 1: mux_24408 = vout_peek_14293;
    endcase
  endfunction
  wire [7:0] v_24409;
  function [7:0] mux_24409(input [0:0] sel);
    case (sel) 0: mux_24409 = 8'h0; 1: mux_24409 = v_24410;
    endcase
  endfunction
  reg [7:0] v_24410 = 8'h0;
  wire [7:0] v_24411;
  wire [7:0] v_24412;
  function [7:0] mux_24412(input [0:0] sel);
    case (sel) 0: mux_24412 = 8'h0; 1: mux_24412 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24413;
  wire [7:0] v_24414;
  wire [7:0] v_24415;
  function [7:0] mux_24415(input [0:0] sel);
    case (sel) 0: mux_24415 = 8'h0; 1: mux_24415 = vout_peek_14265;
    endcase
  endfunction
  wire [7:0] v_24416;
  function [7:0] mux_24416(input [0:0] sel);
    case (sel) 0: mux_24416 = 8'h0; 1: mux_24416 = vout_peek_14256;
    endcase
  endfunction
  wire [7:0] v_24417;
  function [7:0] mux_24417(input [0:0] sel);
    case (sel) 0: mux_24417 = 8'h0; 1: mux_24417 = v_24418;
    endcase
  endfunction
  reg [7:0] v_24418 = 8'h0;
  wire [7:0] v_24419;
  wire [7:0] v_24420;
  function [7:0] mux_24420(input [0:0] sel);
    case (sel) 0: mux_24420 = 8'h0; 1: mux_24420 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24421;
  wire [7:0] v_24422;
  wire [7:0] v_24423;
  function [7:0] mux_24423(input [0:0] sel);
    case (sel) 0: mux_24423 = 8'h0; 1: mux_24423 = v_24424;
    endcase
  endfunction
  reg [7:0] v_24424 = 8'h0;
  wire [7:0] v_24425;
  wire [7:0] v_24426;
  function [7:0] mux_24426(input [0:0] sel);
    case (sel) 0: mux_24426 = 8'h0; 1: mux_24426 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24427;
  wire [7:0] v_24428;
  wire [7:0] v_24429;
  function [7:0] mux_24429(input [0:0] sel);
    case (sel) 0: mux_24429 = 8'h0; 1: mux_24429 = v_24430;
    endcase
  endfunction
  reg [7:0] v_24430 = 8'h0;
  wire [7:0] v_24431;
  wire [7:0] v_24432;
  function [7:0] mux_24432(input [0:0] sel);
    case (sel) 0: mux_24432 = 8'h0; 1: mux_24432 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24433;
  wire [7:0] v_24434;
  wire [7:0] v_24435;
  function [7:0] mux_24435(input [0:0] sel);
    case (sel) 0: mux_24435 = 8'h0; 1: mux_24435 = v_24436;
    endcase
  endfunction
  reg [7:0] v_24436 = 8'h0;
  wire [7:0] v_24437;
  wire [7:0] v_24438;
  function [7:0] mux_24438(input [0:0] sel);
    case (sel) 0: mux_24438 = 8'h0; 1: mux_24438 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24439;
  wire [7:0] v_24440;
  wire [7:0] v_24441;
  function [7:0] mux_24441(input [0:0] sel);
    case (sel) 0: mux_24441 = 8'h0; 1: mux_24441 = v_24442;
    endcase
  endfunction
  reg [7:0] v_24442 = 8'h0;
  wire [7:0] v_24443;
  wire [7:0] v_24444;
  function [7:0] mux_24444(input [0:0] sel);
    case (sel) 0: mux_24444 = 8'h0; 1: mux_24444 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24445;
  wire [7:0] v_24446;
  wire [7:0] v_24447;
  function [7:0] mux_24447(input [0:0] sel);
    case (sel) 0: mux_24447 = 8'h0; 1: mux_24447 = vout_peek_14152;
    endcase
  endfunction
  wire [7:0] v_24448;
  function [7:0] mux_24448(input [0:0] sel);
    case (sel) 0: mux_24448 = 8'h0; 1: mux_24448 = vout_peek_14143;
    endcase
  endfunction
  wire [7:0] v_24449;
  function [7:0] mux_24449(input [0:0] sel);
    case (sel) 0: mux_24449 = 8'h0; 1: mux_24449 = v_24450;
    endcase
  endfunction
  reg [7:0] v_24450 = 8'h0;
  wire [7:0] v_24451;
  wire [7:0] v_24452;
  function [7:0] mux_24452(input [0:0] sel);
    case (sel) 0: mux_24452 = 8'h0; 1: mux_24452 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24453;
  wire [7:0] v_24454;
  wire [7:0] v_24455;
  function [7:0] mux_24455(input [0:0] sel);
    case (sel) 0: mux_24455 = 8'h0; 1: mux_24455 = vout_peek_14115;
    endcase
  endfunction
  wire [7:0] v_24456;
  function [7:0] mux_24456(input [0:0] sel);
    case (sel) 0: mux_24456 = 8'h0; 1: mux_24456 = vout_peek_14106;
    endcase
  endfunction
  wire [7:0] v_24457;
  function [7:0] mux_24457(input [0:0] sel);
    case (sel) 0: mux_24457 = 8'h0; 1: mux_24457 = v_24458;
    endcase
  endfunction
  reg [7:0] v_24458 = 8'h0;
  wire [7:0] v_24459;
  wire [7:0] v_24460;
  function [7:0] mux_24460(input [0:0] sel);
    case (sel) 0: mux_24460 = 8'h0; 1: mux_24460 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24461;
  wire [7:0] v_24462;
  wire [7:0] v_24463;
  function [7:0] mux_24463(input [0:0] sel);
    case (sel) 0: mux_24463 = 8'h0; 1: mux_24463 = v_24464;
    endcase
  endfunction
  reg [7:0] v_24464 = 8'h0;
  wire [7:0] v_24465;
  wire [7:0] v_24466;
  function [7:0] mux_24466(input [0:0] sel);
    case (sel) 0: mux_24466 = 8'h0; 1: mux_24466 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24467;
  wire [7:0] v_24468;
  wire [7:0] v_24469;
  function [7:0] mux_24469(input [0:0] sel);
    case (sel) 0: mux_24469 = 8'h0; 1: mux_24469 = vout_peek_14059;
    endcase
  endfunction
  wire [7:0] v_24470;
  function [7:0] mux_24470(input [0:0] sel);
    case (sel) 0: mux_24470 = 8'h0; 1: mux_24470 = vout_peek_14050;
    endcase
  endfunction
  wire [7:0] v_24471;
  function [7:0] mux_24471(input [0:0] sel);
    case (sel) 0: mux_24471 = 8'h0; 1: mux_24471 = v_24472;
    endcase
  endfunction
  reg [7:0] v_24472 = 8'h0;
  wire [7:0] v_24473;
  wire [7:0] v_24474;
  function [7:0] mux_24474(input [0:0] sel);
    case (sel) 0: mux_24474 = 8'h0; 1: mux_24474 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24475;
  wire [7:0] v_24476;
  wire [7:0] v_24477;
  function [7:0] mux_24477(input [0:0] sel);
    case (sel) 0: mux_24477 = 8'h0; 1: mux_24477 = vout_peek_14022;
    endcase
  endfunction
  wire [7:0] v_24478;
  function [7:0] mux_24478(input [0:0] sel);
    case (sel) 0: mux_24478 = 8'h0; 1: mux_24478 = vout_peek_14013;
    endcase
  endfunction
  wire [7:0] v_24479;
  function [7:0] mux_24479(input [0:0] sel);
    case (sel) 0: mux_24479 = 8'h0; 1: mux_24479 = v_24480;
    endcase
  endfunction
  reg [7:0] v_24480 = 8'h0;
  wire [7:0] v_24481;
  wire [7:0] v_24482;
  function [7:0] mux_24482(input [0:0] sel);
    case (sel) 0: mux_24482 = 8'h0; 1: mux_24482 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24483;
  wire [7:0] v_24484;
  wire [7:0] v_24485;
  function [7:0] mux_24485(input [0:0] sel);
    case (sel) 0: mux_24485 = 8'h0; 1: mux_24485 = v_24486;
    endcase
  endfunction
  reg [7:0] v_24486 = 8'h0;
  wire [7:0] v_24487;
  wire [7:0] v_24488;
  function [7:0] mux_24488(input [0:0] sel);
    case (sel) 0: mux_24488 = 8'h0; 1: mux_24488 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24489;
  wire [7:0] v_24490;
  wire [7:0] v_24491;
  function [7:0] mux_24491(input [0:0] sel);
    case (sel) 0: mux_24491 = 8'h0; 1: mux_24491 = v_24492;
    endcase
  endfunction
  reg [7:0] v_24492 = 8'h0;
  wire [7:0] v_24493;
  wire [7:0] v_24494;
  function [7:0] mux_24494(input [0:0] sel);
    case (sel) 0: mux_24494 = 8'h0; 1: mux_24494 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24495;
  wire [7:0] v_24496;
  wire [7:0] v_24497;
  function [7:0] mux_24497(input [0:0] sel);
    case (sel) 0: mux_24497 = 8'h0; 1: mux_24497 = vout_peek_13947;
    endcase
  endfunction
  wire [7:0] v_24498;
  function [7:0] mux_24498(input [0:0] sel);
    case (sel) 0: mux_24498 = 8'h0; 1: mux_24498 = vout_peek_13938;
    endcase
  endfunction
  wire [7:0] v_24499;
  function [7:0] mux_24499(input [0:0] sel);
    case (sel) 0: mux_24499 = 8'h0; 1: mux_24499 = v_24500;
    endcase
  endfunction
  reg [7:0] v_24500 = 8'h0;
  wire [7:0] v_24501;
  wire [7:0] v_24502;
  function [7:0] mux_24502(input [0:0] sel);
    case (sel) 0: mux_24502 = 8'h0; 1: mux_24502 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24503;
  wire [7:0] v_24504;
  wire [7:0] v_24505;
  function [7:0] mux_24505(input [0:0] sel);
    case (sel) 0: mux_24505 = 8'h0; 1: mux_24505 = vout_peek_13910;
    endcase
  endfunction
  wire [7:0] v_24506;
  function [7:0] mux_24506(input [0:0] sel);
    case (sel) 0: mux_24506 = 8'h0; 1: mux_24506 = vout_peek_13901;
    endcase
  endfunction
  wire [7:0] v_24507;
  function [7:0] mux_24507(input [0:0] sel);
    case (sel) 0: mux_24507 = 8'h0; 1: mux_24507 = v_24508;
    endcase
  endfunction
  reg [7:0] v_24508 = 8'h0;
  wire [7:0] v_24509;
  wire [7:0] v_24510;
  function [7:0] mux_24510(input [0:0] sel);
    case (sel) 0: mux_24510 = 8'h0; 1: mux_24510 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24511;
  wire [7:0] v_24512;
  wire [7:0] v_24513;
  function [7:0] mux_24513(input [0:0] sel);
    case (sel) 0: mux_24513 = 8'h0; 1: mux_24513 = v_24514;
    endcase
  endfunction
  reg [7:0] v_24514 = 8'h0;
  wire [7:0] v_24515;
  wire [7:0] v_24516;
  function [7:0] mux_24516(input [0:0] sel);
    case (sel) 0: mux_24516 = 8'h0; 1: mux_24516 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24517;
  wire [7:0] v_24518;
  wire [7:0] v_24519;
  function [7:0] mux_24519(input [0:0] sel);
    case (sel) 0: mux_24519 = 8'h0; 1: mux_24519 = vout_peek_13854;
    endcase
  endfunction
  wire [7:0] v_24520;
  function [7:0] mux_24520(input [0:0] sel);
    case (sel) 0: mux_24520 = 8'h0; 1: mux_24520 = vout_peek_13845;
    endcase
  endfunction
  wire [7:0] v_24521;
  function [7:0] mux_24521(input [0:0] sel);
    case (sel) 0: mux_24521 = 8'h0; 1: mux_24521 = v_24522;
    endcase
  endfunction
  reg [7:0] v_24522 = 8'h0;
  wire [7:0] v_24523;
  wire [7:0] v_24524;
  function [7:0] mux_24524(input [0:0] sel);
    case (sel) 0: mux_24524 = 8'h0; 1: mux_24524 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24525;
  wire [7:0] v_24526;
  wire [7:0] v_24527;
  function [7:0] mux_24527(input [0:0] sel);
    case (sel) 0: mux_24527 = 8'h0; 1: mux_24527 = vout_peek_13817;
    endcase
  endfunction
  wire [7:0] v_24528;
  function [7:0] mux_24528(input [0:0] sel);
    case (sel) 0: mux_24528 = 8'h0; 1: mux_24528 = vout_peek_13808;
    endcase
  endfunction
  wire [7:0] v_24529;
  function [7:0] mux_24529(input [0:0] sel);
    case (sel) 0: mux_24529 = 8'h0; 1: mux_24529 = v_24530;
    endcase
  endfunction
  reg [7:0] v_24530 = 8'h0;
  wire [7:0] v_24531;
  wire [7:0] v_24532;
  function [7:0] mux_24532(input [0:0] sel);
    case (sel) 0: mux_24532 = 8'h0; 1: mux_24532 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24533;
  wire [7:0] v_24534;
  wire [7:0] v_24535;
  function [7:0] mux_24535(input [0:0] sel);
    case (sel) 0: mux_24535 = 8'h0; 1: mux_24535 = v_24536;
    endcase
  endfunction
  reg [7:0] v_24536 = 8'h0;
  wire [7:0] v_24537;
  wire [7:0] v_24538;
  function [7:0] mux_24538(input [0:0] sel);
    case (sel) 0: mux_24538 = 8'h0; 1: mux_24538 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24539;
  wire [7:0] v_24540;
  wire [7:0] v_24541;
  function [7:0] mux_24541(input [0:0] sel);
    case (sel) 0: mux_24541 = 8'h0; 1: mux_24541 = v_24542;
    endcase
  endfunction
  reg [7:0] v_24542 = 8'h0;
  wire [7:0] v_24543;
  wire [7:0] v_24544;
  function [7:0] mux_24544(input [0:0] sel);
    case (sel) 0: mux_24544 = 8'h0; 1: mux_24544 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24545;
  wire [7:0] v_24546;
  wire [7:0] v_24547;
  function [7:0] mux_24547(input [0:0] sel);
    case (sel) 0: mux_24547 = 8'h0; 1: mux_24547 = v_24548;
    endcase
  endfunction
  reg [7:0] v_24548 = 8'h0;
  wire [7:0] v_24549;
  wire [7:0] v_24550;
  function [7:0] mux_24550(input [0:0] sel);
    case (sel) 0: mux_24550 = 8'h0; 1: mux_24550 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24551;
  wire [7:0] v_24552;
  wire [7:0] v_24553;
  function [7:0] mux_24553(input [0:0] sel);
    case (sel) 0: mux_24553 = 8'h0; 1: mux_24553 = vout_peek_13723;
    endcase
  endfunction
  wire [7:0] v_24554;
  function [7:0] mux_24554(input [0:0] sel);
    case (sel) 0: mux_24554 = 8'h0; 1: mux_24554 = vout_peek_13714;
    endcase
  endfunction
  wire [7:0] v_24555;
  function [7:0] mux_24555(input [0:0] sel);
    case (sel) 0: mux_24555 = 8'h0; 1: mux_24555 = v_24556;
    endcase
  endfunction
  reg [7:0] v_24556 = 8'h0;
  wire [7:0] v_24557;
  wire [7:0] v_24558;
  function [7:0] mux_24558(input [0:0] sel);
    case (sel) 0: mux_24558 = 8'h0; 1: mux_24558 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24559;
  wire [7:0] v_24560;
  wire [7:0] v_24561;
  function [7:0] mux_24561(input [0:0] sel);
    case (sel) 0: mux_24561 = 8'h0; 1: mux_24561 = vout_peek_13686;
    endcase
  endfunction
  wire [7:0] v_24562;
  function [7:0] mux_24562(input [0:0] sel);
    case (sel) 0: mux_24562 = 8'h0; 1: mux_24562 = vout_peek_13677;
    endcase
  endfunction
  wire [7:0] v_24563;
  function [7:0] mux_24563(input [0:0] sel);
    case (sel) 0: mux_24563 = 8'h0; 1: mux_24563 = v_24564;
    endcase
  endfunction
  reg [7:0] v_24564 = 8'h0;
  wire [7:0] v_24565;
  wire [7:0] v_24566;
  function [7:0] mux_24566(input [0:0] sel);
    case (sel) 0: mux_24566 = 8'h0; 1: mux_24566 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24567;
  wire [7:0] v_24568;
  wire [7:0] v_24569;
  function [7:0] mux_24569(input [0:0] sel);
    case (sel) 0: mux_24569 = 8'h0; 1: mux_24569 = v_24570;
    endcase
  endfunction
  reg [7:0] v_24570 = 8'h0;
  wire [7:0] v_24571;
  wire [7:0] v_24572;
  function [7:0] mux_24572(input [0:0] sel);
    case (sel) 0: mux_24572 = 8'h0; 1: mux_24572 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24573;
  wire [7:0] v_24574;
  wire [7:0] v_24575;
  function [7:0] mux_24575(input [0:0] sel);
    case (sel) 0: mux_24575 = 8'h0; 1: mux_24575 = vout_peek_13630;
    endcase
  endfunction
  wire [7:0] v_24576;
  function [7:0] mux_24576(input [0:0] sel);
    case (sel) 0: mux_24576 = 8'h0; 1: mux_24576 = vout_peek_13621;
    endcase
  endfunction
  wire [7:0] v_24577;
  function [7:0] mux_24577(input [0:0] sel);
    case (sel) 0: mux_24577 = 8'h0; 1: mux_24577 = v_24578;
    endcase
  endfunction
  reg [7:0] v_24578 = 8'h0;
  wire [7:0] v_24579;
  wire [7:0] v_24580;
  function [7:0] mux_24580(input [0:0] sel);
    case (sel) 0: mux_24580 = 8'h0; 1: mux_24580 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24581;
  wire [7:0] v_24582;
  wire [7:0] v_24583;
  function [7:0] mux_24583(input [0:0] sel);
    case (sel) 0: mux_24583 = 8'h0; 1: mux_24583 = vout_peek_13593;
    endcase
  endfunction
  wire [7:0] v_24584;
  function [7:0] mux_24584(input [0:0] sel);
    case (sel) 0: mux_24584 = 8'h0; 1: mux_24584 = vout_peek_13584;
    endcase
  endfunction
  wire [7:0] v_24585;
  function [7:0] mux_24585(input [0:0] sel);
    case (sel) 0: mux_24585 = 8'h0; 1: mux_24585 = v_24586;
    endcase
  endfunction
  reg [7:0] v_24586 = 8'h0;
  wire [7:0] v_24587;
  wire [7:0] v_24588;
  function [7:0] mux_24588(input [0:0] sel);
    case (sel) 0: mux_24588 = 8'h0; 1: mux_24588 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24589;
  wire [7:0] v_24590;
  wire [7:0] v_24591;
  function [7:0] mux_24591(input [0:0] sel);
    case (sel) 0: mux_24591 = 8'h0; 1: mux_24591 = v_24592;
    endcase
  endfunction
  reg [7:0] v_24592 = 8'h0;
  wire [7:0] v_24593;
  wire [7:0] v_24594;
  function [7:0] mux_24594(input [0:0] sel);
    case (sel) 0: mux_24594 = 8'h0; 1: mux_24594 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24595;
  wire [7:0] v_24596;
  wire [7:0] v_24597;
  function [7:0] mux_24597(input [0:0] sel);
    case (sel) 0: mux_24597 = 8'h0; 1: mux_24597 = v_24598;
    endcase
  endfunction
  reg [7:0] v_24598 = 8'h0;
  wire [7:0] v_24599;
  wire [7:0] v_24600;
  function [7:0] mux_24600(input [0:0] sel);
    case (sel) 0: mux_24600 = 8'h0; 1: mux_24600 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24601;
  wire [7:0] v_24602;
  wire [7:0] v_24603;
  function [7:0] mux_24603(input [0:0] sel);
    case (sel) 0: mux_24603 = 8'h0; 1: mux_24603 = vout_peek_13518;
    endcase
  endfunction
  wire [7:0] v_24604;
  function [7:0] mux_24604(input [0:0] sel);
    case (sel) 0: mux_24604 = 8'h0; 1: mux_24604 = vout_peek_13509;
    endcase
  endfunction
  wire [7:0] v_24605;
  function [7:0] mux_24605(input [0:0] sel);
    case (sel) 0: mux_24605 = 8'h0; 1: mux_24605 = v_24606;
    endcase
  endfunction
  reg [7:0] v_24606 = 8'h0;
  wire [7:0] v_24607;
  wire [7:0] v_24608;
  function [7:0] mux_24608(input [0:0] sel);
    case (sel) 0: mux_24608 = 8'h0; 1: mux_24608 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24609;
  wire [7:0] v_24610;
  wire [7:0] v_24611;
  function [7:0] mux_24611(input [0:0] sel);
    case (sel) 0: mux_24611 = 8'h0; 1: mux_24611 = vout_peek_13481;
    endcase
  endfunction
  wire [7:0] v_24612;
  function [7:0] mux_24612(input [0:0] sel);
    case (sel) 0: mux_24612 = 8'h0; 1: mux_24612 = vout_peek_13472;
    endcase
  endfunction
  wire [7:0] v_24613;
  function [7:0] mux_24613(input [0:0] sel);
    case (sel) 0: mux_24613 = 8'h0; 1: mux_24613 = v_24614;
    endcase
  endfunction
  reg [7:0] v_24614 = 8'h0;
  wire [7:0] v_24615;
  wire [7:0] v_24616;
  function [7:0] mux_24616(input [0:0] sel);
    case (sel) 0: mux_24616 = 8'h0; 1: mux_24616 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24617;
  wire [7:0] v_24618;
  wire [7:0] v_24619;
  function [7:0] mux_24619(input [0:0] sel);
    case (sel) 0: mux_24619 = 8'h0; 1: mux_24619 = v_24620;
    endcase
  endfunction
  reg [7:0] v_24620 = 8'h0;
  wire [7:0] v_24621;
  wire [7:0] v_24622;
  function [7:0] mux_24622(input [0:0] sel);
    case (sel) 0: mux_24622 = 8'h0; 1: mux_24622 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24623;
  wire [7:0] v_24624;
  wire [7:0] v_24625;
  function [7:0] mux_24625(input [0:0] sel);
    case (sel) 0: mux_24625 = 8'h0; 1: mux_24625 = vout_peek_13425;
    endcase
  endfunction
  wire [7:0] v_24626;
  function [7:0] mux_24626(input [0:0] sel);
    case (sel) 0: mux_24626 = 8'h0; 1: mux_24626 = vout_peek_13416;
    endcase
  endfunction
  wire [7:0] v_24627;
  function [7:0] mux_24627(input [0:0] sel);
    case (sel) 0: mux_24627 = 8'h0; 1: mux_24627 = v_24628;
    endcase
  endfunction
  reg [7:0] v_24628 = 8'h0;
  wire [7:0] v_24629;
  wire [7:0] v_24630;
  function [7:0] mux_24630(input [0:0] sel);
    case (sel) 0: mux_24630 = 8'h0; 1: mux_24630 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24631;
  wire [7:0] v_24632;
  wire [7:0] v_24633;
  function [7:0] mux_24633(input [0:0] sel);
    case (sel) 0: mux_24633 = 8'h0; 1: mux_24633 = vout_peek_13388;
    endcase
  endfunction
  wire [7:0] v_24634;
  function [7:0] mux_24634(input [0:0] sel);
    case (sel) 0: mux_24634 = 8'h0; 1: mux_24634 = vout_peek_13379;
    endcase
  endfunction
  wire [7:0] v_24635;
  function [7:0] mux_24635(input [0:0] sel);
    case (sel) 0: mux_24635 = 8'h0; 1: mux_24635 = v_24636;
    endcase
  endfunction
  reg [7:0] v_24636 = 8'h0;
  wire [7:0] v_24637;
  wire [7:0] v_24638;
  function [7:0] mux_24638(input [0:0] sel);
    case (sel) 0: mux_24638 = 8'h0; 1: mux_24638 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24639;
  wire [7:0] v_24640;
  wire [7:0] v_24641;
  function [7:0] mux_24641(input [0:0] sel);
    case (sel) 0: mux_24641 = 8'h0; 1: mux_24641 = v_24642;
    endcase
  endfunction
  reg [7:0] v_24642 = 8'h0;
  wire [7:0] v_24643;
  wire [7:0] v_24644;
  function [7:0] mux_24644(input [0:0] sel);
    case (sel) 0: mux_24644 = 8'h0; 1: mux_24644 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24645;
  wire [7:0] v_24646;
  wire [7:0] v_24647;
  function [7:0] mux_24647(input [0:0] sel);
    case (sel) 0: mux_24647 = 8'h0; 1: mux_24647 = v_24648;
    endcase
  endfunction
  reg [7:0] v_24648 = 8'h0;
  wire [7:0] v_24649;
  wire [7:0] v_24650;
  function [7:0] mux_24650(input [0:0] sel);
    case (sel) 0: mux_24650 = 8'h0; 1: mux_24650 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24651;
  wire [7:0] v_24652;
  wire [7:0] v_24653;
  function [7:0] mux_24653(input [0:0] sel);
    case (sel) 0: mux_24653 = 8'h0; 1: mux_24653 = v_24654;
    endcase
  endfunction
  reg [7:0] v_24654 = 8'h0;
  wire [7:0] v_24655;
  wire [7:0] v_24656;
  function [7:0] mux_24656(input [0:0] sel);
    case (sel) 0: mux_24656 = 8'h0; 1: mux_24656 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24657;
  wire [7:0] v_24658;
  wire [7:0] v_24659;
  function [7:0] mux_24659(input [0:0] sel);
    case (sel) 0: mux_24659 = 8'h0; 1: mux_24659 = v_24660;
    endcase
  endfunction
  reg [7:0] v_24660 = 8'h0;
  wire [7:0] v_24661;
  wire [7:0] v_24662;
  function [7:0] mux_24662(input [0:0] sel);
    case (sel) 0: mux_24662 = 8'h0; 1: mux_24662 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24663;
  wire [7:0] v_24664;
  wire [7:0] v_24665;
  function [7:0] mux_24665(input [0:0] sel);
    case (sel) 0: mux_24665 = 8'h0; 1: mux_24665 = v_24666;
    endcase
  endfunction
  reg [7:0] v_24666 = 8'h0;
  wire [7:0] v_24667;
  wire [7:0] v_24668;
  function [7:0] mux_24668(input [0:0] sel);
    case (sel) 0: mux_24668 = 8'h0; 1: mux_24668 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24669;
  wire [7:0] v_24670;
  wire [7:0] v_24671;
  function [7:0] mux_24671(input [0:0] sel);
    case (sel) 0: mux_24671 = 8'h0; 1: mux_24671 = vout_peek_13256;
    endcase
  endfunction
  wire [7:0] v_24672;
  function [7:0] mux_24672(input [0:0] sel);
    case (sel) 0: mux_24672 = 8'h0; 1: mux_24672 = vout_peek_13247;
    endcase
  endfunction
  wire [7:0] v_24673;
  function [7:0] mux_24673(input [0:0] sel);
    case (sel) 0: mux_24673 = 8'h0; 1: mux_24673 = v_24674;
    endcase
  endfunction
  reg [7:0] v_24674 = 8'h0;
  wire [7:0] v_24675;
  wire [7:0] v_24676;
  function [7:0] mux_24676(input [0:0] sel);
    case (sel) 0: mux_24676 = 8'h0; 1: mux_24676 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24677;
  wire [7:0] v_24678;
  wire [7:0] v_24679;
  function [7:0] mux_24679(input [0:0] sel);
    case (sel) 0: mux_24679 = 8'h0; 1: mux_24679 = vout_peek_13219;
    endcase
  endfunction
  wire [7:0] v_24680;
  function [7:0] mux_24680(input [0:0] sel);
    case (sel) 0: mux_24680 = 8'h0; 1: mux_24680 = vout_peek_13210;
    endcase
  endfunction
  wire [7:0] v_24681;
  function [7:0] mux_24681(input [0:0] sel);
    case (sel) 0: mux_24681 = 8'h0; 1: mux_24681 = v_24682;
    endcase
  endfunction
  reg [7:0] v_24682 = 8'h0;
  wire [7:0] v_24683;
  wire [7:0] v_24684;
  function [7:0] mux_24684(input [0:0] sel);
    case (sel) 0: mux_24684 = 8'h0; 1: mux_24684 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24685;
  wire [7:0] v_24686;
  wire [7:0] v_24687;
  function [7:0] mux_24687(input [0:0] sel);
    case (sel) 0: mux_24687 = 8'h0; 1: mux_24687 = v_24688;
    endcase
  endfunction
  reg [7:0] v_24688 = 8'h0;
  wire [7:0] v_24689;
  wire [7:0] v_24690;
  function [7:0] mux_24690(input [0:0] sel);
    case (sel) 0: mux_24690 = 8'h0; 1: mux_24690 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24691;
  wire [7:0] v_24692;
  wire [7:0] v_24693;
  function [7:0] mux_24693(input [0:0] sel);
    case (sel) 0: mux_24693 = 8'h0; 1: mux_24693 = vout_peek_13163;
    endcase
  endfunction
  wire [7:0] v_24694;
  function [7:0] mux_24694(input [0:0] sel);
    case (sel) 0: mux_24694 = 8'h0; 1: mux_24694 = vout_peek_13154;
    endcase
  endfunction
  wire [7:0] v_24695;
  function [7:0] mux_24695(input [0:0] sel);
    case (sel) 0: mux_24695 = 8'h0; 1: mux_24695 = v_24696;
    endcase
  endfunction
  reg [7:0] v_24696 = 8'h0;
  wire [7:0] v_24697;
  wire [7:0] v_24698;
  function [7:0] mux_24698(input [0:0] sel);
    case (sel) 0: mux_24698 = 8'h0; 1: mux_24698 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24699;
  wire [7:0] v_24700;
  wire [7:0] v_24701;
  function [7:0] mux_24701(input [0:0] sel);
    case (sel) 0: mux_24701 = 8'h0; 1: mux_24701 = vout_peek_13126;
    endcase
  endfunction
  wire [7:0] v_24702;
  function [7:0] mux_24702(input [0:0] sel);
    case (sel) 0: mux_24702 = 8'h0; 1: mux_24702 = vout_peek_13117;
    endcase
  endfunction
  wire [7:0] v_24703;
  function [7:0] mux_24703(input [0:0] sel);
    case (sel) 0: mux_24703 = 8'h0; 1: mux_24703 = v_24704;
    endcase
  endfunction
  reg [7:0] v_24704 = 8'h0;
  wire [7:0] v_24705;
  wire [7:0] v_24706;
  function [7:0] mux_24706(input [0:0] sel);
    case (sel) 0: mux_24706 = 8'h0; 1: mux_24706 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24707;
  wire [7:0] v_24708;
  wire [7:0] v_24709;
  function [7:0] mux_24709(input [0:0] sel);
    case (sel) 0: mux_24709 = 8'h0; 1: mux_24709 = v_24710;
    endcase
  endfunction
  reg [7:0] v_24710 = 8'h0;
  wire [7:0] v_24711;
  wire [7:0] v_24712;
  function [7:0] mux_24712(input [0:0] sel);
    case (sel) 0: mux_24712 = 8'h0; 1: mux_24712 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24713;
  wire [7:0] v_24714;
  wire [7:0] v_24715;
  function [7:0] mux_24715(input [0:0] sel);
    case (sel) 0: mux_24715 = 8'h0; 1: mux_24715 = v_24716;
    endcase
  endfunction
  reg [7:0] v_24716 = 8'h0;
  wire [7:0] v_24717;
  wire [7:0] v_24718;
  function [7:0] mux_24718(input [0:0] sel);
    case (sel) 0: mux_24718 = 8'h0; 1: mux_24718 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24719;
  wire [7:0] v_24720;
  wire [7:0] v_24721;
  function [7:0] mux_24721(input [0:0] sel);
    case (sel) 0: mux_24721 = 8'h0; 1: mux_24721 = vout_peek_13051;
    endcase
  endfunction
  wire [7:0] v_24722;
  function [7:0] mux_24722(input [0:0] sel);
    case (sel) 0: mux_24722 = 8'h0; 1: mux_24722 = vout_peek_13042;
    endcase
  endfunction
  wire [7:0] v_24723;
  function [7:0] mux_24723(input [0:0] sel);
    case (sel) 0: mux_24723 = 8'h0; 1: mux_24723 = v_24724;
    endcase
  endfunction
  reg [7:0] v_24724 = 8'h0;
  wire [7:0] v_24725;
  wire [7:0] v_24726;
  function [7:0] mux_24726(input [0:0] sel);
    case (sel) 0: mux_24726 = 8'h0; 1: mux_24726 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24727;
  wire [7:0] v_24728;
  wire [7:0] v_24729;
  function [7:0] mux_24729(input [0:0] sel);
    case (sel) 0: mux_24729 = 8'h0; 1: mux_24729 = vout_peek_13014;
    endcase
  endfunction
  wire [7:0] v_24730;
  function [7:0] mux_24730(input [0:0] sel);
    case (sel) 0: mux_24730 = 8'h0; 1: mux_24730 = vout_peek_13005;
    endcase
  endfunction
  wire [7:0] v_24731;
  function [7:0] mux_24731(input [0:0] sel);
    case (sel) 0: mux_24731 = 8'h0; 1: mux_24731 = v_24732;
    endcase
  endfunction
  reg [7:0] v_24732 = 8'h0;
  wire [7:0] v_24733;
  wire [7:0] v_24734;
  function [7:0] mux_24734(input [0:0] sel);
    case (sel) 0: mux_24734 = 8'h0; 1: mux_24734 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24735;
  wire [7:0] v_24736;
  wire [7:0] v_24737;
  function [7:0] mux_24737(input [0:0] sel);
    case (sel) 0: mux_24737 = 8'h0; 1: mux_24737 = v_24738;
    endcase
  endfunction
  reg [7:0] v_24738 = 8'h0;
  wire [7:0] v_24739;
  wire [7:0] v_24740;
  function [7:0] mux_24740(input [0:0] sel);
    case (sel) 0: mux_24740 = 8'h0; 1: mux_24740 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24741;
  wire [7:0] v_24742;
  wire [7:0] v_24743;
  function [7:0] mux_24743(input [0:0] sel);
    case (sel) 0: mux_24743 = 8'h0; 1: mux_24743 = vout_peek_12958;
    endcase
  endfunction
  wire [7:0] v_24744;
  function [7:0] mux_24744(input [0:0] sel);
    case (sel) 0: mux_24744 = 8'h0; 1: mux_24744 = vout_peek_12949;
    endcase
  endfunction
  wire [7:0] v_24745;
  function [7:0] mux_24745(input [0:0] sel);
    case (sel) 0: mux_24745 = 8'h0; 1: mux_24745 = v_24746;
    endcase
  endfunction
  reg [7:0] v_24746 = 8'h0;
  wire [7:0] v_24747;
  wire [7:0] v_24748;
  function [7:0] mux_24748(input [0:0] sel);
    case (sel) 0: mux_24748 = 8'h0; 1: mux_24748 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24749;
  wire [7:0] v_24750;
  wire [7:0] v_24751;
  function [7:0] mux_24751(input [0:0] sel);
    case (sel) 0: mux_24751 = 8'h0; 1: mux_24751 = vout_peek_12921;
    endcase
  endfunction
  wire [7:0] v_24752;
  function [7:0] mux_24752(input [0:0] sel);
    case (sel) 0: mux_24752 = 8'h0; 1: mux_24752 = vout_peek_12912;
    endcase
  endfunction
  wire [7:0] v_24753;
  function [7:0] mux_24753(input [0:0] sel);
    case (sel) 0: mux_24753 = 8'h0; 1: mux_24753 = v_24754;
    endcase
  endfunction
  reg [7:0] v_24754 = 8'h0;
  wire [7:0] v_24755;
  wire [7:0] v_24756;
  function [7:0] mux_24756(input [0:0] sel);
    case (sel) 0: mux_24756 = 8'h0; 1: mux_24756 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24757;
  wire [7:0] v_24758;
  wire [7:0] v_24759;
  function [7:0] mux_24759(input [0:0] sel);
    case (sel) 0: mux_24759 = 8'h0; 1: mux_24759 = v_24760;
    endcase
  endfunction
  reg [7:0] v_24760 = 8'h0;
  wire [7:0] v_24761;
  wire [7:0] v_24762;
  function [7:0] mux_24762(input [0:0] sel);
    case (sel) 0: mux_24762 = 8'h0; 1: mux_24762 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24763;
  wire [7:0] v_24764;
  wire [7:0] v_24765;
  function [7:0] mux_24765(input [0:0] sel);
    case (sel) 0: mux_24765 = 8'h0; 1: mux_24765 = v_24766;
    endcase
  endfunction
  reg [7:0] v_24766 = 8'h0;
  wire [7:0] v_24767;
  wire [7:0] v_24768;
  function [7:0] mux_24768(input [0:0] sel);
    case (sel) 0: mux_24768 = 8'h0; 1: mux_24768 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24769;
  wire [7:0] v_24770;
  wire [7:0] v_24771;
  function [7:0] mux_24771(input [0:0] sel);
    case (sel) 0: mux_24771 = 8'h0; 1: mux_24771 = v_24772;
    endcase
  endfunction
  reg [7:0] v_24772 = 8'h0;
  wire [7:0] v_24773;
  wire [7:0] v_24774;
  function [7:0] mux_24774(input [0:0] sel);
    case (sel) 0: mux_24774 = 8'h0; 1: mux_24774 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24775;
  wire [7:0] v_24776;
  wire [7:0] v_24777;
  function [7:0] mux_24777(input [0:0] sel);
    case (sel) 0: mux_24777 = 8'h0; 1: mux_24777 = vout_peek_12827;
    endcase
  endfunction
  wire [7:0] v_24778;
  function [7:0] mux_24778(input [0:0] sel);
    case (sel) 0: mux_24778 = 8'h0; 1: mux_24778 = vout_peek_12818;
    endcase
  endfunction
  wire [7:0] v_24779;
  function [7:0] mux_24779(input [0:0] sel);
    case (sel) 0: mux_24779 = 8'h0; 1: mux_24779 = v_24780;
    endcase
  endfunction
  reg [7:0] v_24780 = 8'h0;
  wire [7:0] v_24781;
  wire [7:0] v_24782;
  function [7:0] mux_24782(input [0:0] sel);
    case (sel) 0: mux_24782 = 8'h0; 1: mux_24782 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24783;
  wire [7:0] v_24784;
  wire [7:0] v_24785;
  function [7:0] mux_24785(input [0:0] sel);
    case (sel) 0: mux_24785 = 8'h0; 1: mux_24785 = vout_peek_12790;
    endcase
  endfunction
  wire [7:0] v_24786;
  function [7:0] mux_24786(input [0:0] sel);
    case (sel) 0: mux_24786 = 8'h0; 1: mux_24786 = vout_peek_12781;
    endcase
  endfunction
  wire [7:0] v_24787;
  function [7:0] mux_24787(input [0:0] sel);
    case (sel) 0: mux_24787 = 8'h0; 1: mux_24787 = v_24788;
    endcase
  endfunction
  reg [7:0] v_24788 = 8'h0;
  wire [7:0] v_24789;
  wire [7:0] v_24790;
  function [7:0] mux_24790(input [0:0] sel);
    case (sel) 0: mux_24790 = 8'h0; 1: mux_24790 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24791;
  wire [7:0] v_24792;
  wire [7:0] v_24793;
  function [7:0] mux_24793(input [0:0] sel);
    case (sel) 0: mux_24793 = 8'h0; 1: mux_24793 = v_24794;
    endcase
  endfunction
  reg [7:0] v_24794 = 8'h0;
  wire [7:0] v_24795;
  wire [7:0] v_24796;
  function [7:0] mux_24796(input [0:0] sel);
    case (sel) 0: mux_24796 = 8'h0; 1: mux_24796 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24797;
  wire [7:0] v_24798;
  wire [7:0] v_24799;
  function [7:0] mux_24799(input [0:0] sel);
    case (sel) 0: mux_24799 = 8'h0; 1: mux_24799 = vout_peek_12734;
    endcase
  endfunction
  wire [7:0] v_24800;
  function [7:0] mux_24800(input [0:0] sel);
    case (sel) 0: mux_24800 = 8'h0; 1: mux_24800 = vout_peek_12725;
    endcase
  endfunction
  wire [7:0] v_24801;
  function [7:0] mux_24801(input [0:0] sel);
    case (sel) 0: mux_24801 = 8'h0; 1: mux_24801 = v_24802;
    endcase
  endfunction
  reg [7:0] v_24802 = 8'h0;
  wire [7:0] v_24803;
  wire [7:0] v_24804;
  function [7:0] mux_24804(input [0:0] sel);
    case (sel) 0: mux_24804 = 8'h0; 1: mux_24804 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24805;
  wire [7:0] v_24806;
  wire [7:0] v_24807;
  function [7:0] mux_24807(input [0:0] sel);
    case (sel) 0: mux_24807 = 8'h0; 1: mux_24807 = vout_peek_12697;
    endcase
  endfunction
  wire [7:0] v_24808;
  function [7:0] mux_24808(input [0:0] sel);
    case (sel) 0: mux_24808 = 8'h0; 1: mux_24808 = vout_peek_12688;
    endcase
  endfunction
  wire [7:0] v_24809;
  function [7:0] mux_24809(input [0:0] sel);
    case (sel) 0: mux_24809 = 8'h0; 1: mux_24809 = v_24810;
    endcase
  endfunction
  reg [7:0] v_24810 = 8'h0;
  wire [7:0] v_24811;
  wire [7:0] v_24812;
  function [7:0] mux_24812(input [0:0] sel);
    case (sel) 0: mux_24812 = 8'h0; 1: mux_24812 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24813;
  wire [7:0] v_24814;
  wire [7:0] v_24815;
  function [7:0] mux_24815(input [0:0] sel);
    case (sel) 0: mux_24815 = 8'h0; 1: mux_24815 = v_24816;
    endcase
  endfunction
  reg [7:0] v_24816 = 8'h0;
  wire [7:0] v_24817;
  wire [7:0] v_24818;
  function [7:0] mux_24818(input [0:0] sel);
    case (sel) 0: mux_24818 = 8'h0; 1: mux_24818 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24819;
  wire [7:0] v_24820;
  wire [7:0] v_24821;
  function [7:0] mux_24821(input [0:0] sel);
    case (sel) 0: mux_24821 = 8'h0; 1: mux_24821 = v_24822;
    endcase
  endfunction
  reg [7:0] v_24822 = 8'h0;
  wire [7:0] v_24823;
  wire [7:0] v_24824;
  function [7:0] mux_24824(input [0:0] sel);
    case (sel) 0: mux_24824 = 8'h0; 1: mux_24824 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24825;
  wire [7:0] v_24826;
  wire [7:0] v_24827;
  function [7:0] mux_24827(input [0:0] sel);
    case (sel) 0: mux_24827 = 8'h0; 1: mux_24827 = vout_peek_12622;
    endcase
  endfunction
  wire [7:0] v_24828;
  function [7:0] mux_24828(input [0:0] sel);
    case (sel) 0: mux_24828 = 8'h0; 1: mux_24828 = vout_peek_12613;
    endcase
  endfunction
  wire [7:0] v_24829;
  function [7:0] mux_24829(input [0:0] sel);
    case (sel) 0: mux_24829 = 8'h0; 1: mux_24829 = v_24830;
    endcase
  endfunction
  reg [7:0] v_24830 = 8'h0;
  wire [7:0] v_24831;
  wire [7:0] v_24832;
  function [7:0] mux_24832(input [0:0] sel);
    case (sel) 0: mux_24832 = 8'h0; 1: mux_24832 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24833;
  wire [7:0] v_24834;
  wire [7:0] v_24835;
  function [7:0] mux_24835(input [0:0] sel);
    case (sel) 0: mux_24835 = 8'h0; 1: mux_24835 = vout_peek_12585;
    endcase
  endfunction
  wire [7:0] v_24836;
  function [7:0] mux_24836(input [0:0] sel);
    case (sel) 0: mux_24836 = 8'h0; 1: mux_24836 = vout_peek_12576;
    endcase
  endfunction
  wire [7:0] v_24837;
  function [7:0] mux_24837(input [0:0] sel);
    case (sel) 0: mux_24837 = 8'h0; 1: mux_24837 = v_24838;
    endcase
  endfunction
  reg [7:0] v_24838 = 8'h0;
  wire [7:0] v_24839;
  wire [7:0] v_24840;
  function [7:0] mux_24840(input [0:0] sel);
    case (sel) 0: mux_24840 = 8'h0; 1: mux_24840 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24841;
  wire [7:0] v_24842;
  wire [7:0] v_24843;
  function [7:0] mux_24843(input [0:0] sel);
    case (sel) 0: mux_24843 = 8'h0; 1: mux_24843 = v_24844;
    endcase
  endfunction
  reg [7:0] v_24844 = 8'h0;
  wire [7:0] v_24845;
  wire [7:0] v_24846;
  function [7:0] mux_24846(input [0:0] sel);
    case (sel) 0: mux_24846 = 8'h0; 1: mux_24846 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24847;
  wire [7:0] v_24848;
  wire [7:0] v_24849;
  function [7:0] mux_24849(input [0:0] sel);
    case (sel) 0: mux_24849 = 8'h0; 1: mux_24849 = vout_peek_12529;
    endcase
  endfunction
  wire [7:0] v_24850;
  function [7:0] mux_24850(input [0:0] sel);
    case (sel) 0: mux_24850 = 8'h0; 1: mux_24850 = vout_peek_12520;
    endcase
  endfunction
  wire [7:0] v_24851;
  function [7:0] mux_24851(input [0:0] sel);
    case (sel) 0: mux_24851 = 8'h0; 1: mux_24851 = v_24852;
    endcase
  endfunction
  reg [7:0] v_24852 = 8'h0;
  wire [7:0] v_24853;
  wire [7:0] v_24854;
  function [7:0] mux_24854(input [0:0] sel);
    case (sel) 0: mux_24854 = 8'h0; 1: mux_24854 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24855;
  wire [7:0] v_24856;
  wire [7:0] v_24857;
  function [7:0] mux_24857(input [0:0] sel);
    case (sel) 0: mux_24857 = 8'h0; 1: mux_24857 = vout_peek_12492;
    endcase
  endfunction
  wire [7:0] v_24858;
  function [7:0] mux_24858(input [0:0] sel);
    case (sel) 0: mux_24858 = 8'h0; 1: mux_24858 = vout_peek_12483;
    endcase
  endfunction
  wire [7:0] v_24859;
  function [7:0] mux_24859(input [0:0] sel);
    case (sel) 0: mux_24859 = 8'h0; 1: mux_24859 = v_24860;
    endcase
  endfunction
  reg [7:0] v_24860 = 8'h0;
  wire [7:0] v_24861;
  wire [7:0] v_24862;
  function [7:0] mux_24862(input [0:0] sel);
    case (sel) 0: mux_24862 = 8'h0; 1: mux_24862 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24863;
  wire [7:0] v_24864;
  wire [7:0] v_24865;
  function [7:0] mux_24865(input [0:0] sel);
    case (sel) 0: mux_24865 = 8'h0; 1: mux_24865 = v_24866;
    endcase
  endfunction
  reg [7:0] v_24866 = 8'h0;
  wire [7:0] v_24867;
  wire [7:0] v_24868;
  function [7:0] mux_24868(input [0:0] sel);
    case (sel) 0: mux_24868 = 8'h0; 1: mux_24868 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24869;
  wire [7:0] v_24870;
  wire [7:0] v_24871;
  function [7:0] mux_24871(input [0:0] sel);
    case (sel) 0: mux_24871 = 8'h0; 1: mux_24871 = v_24872;
    endcase
  endfunction
  reg [7:0] v_24872 = 8'h0;
  wire [7:0] v_24873;
  wire [7:0] v_24874;
  function [7:0] mux_24874(input [0:0] sel);
    case (sel) 0: mux_24874 = 8'h0; 1: mux_24874 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24875;
  wire [7:0] v_24876;
  wire [7:0] v_24877;
  function [7:0] mux_24877(input [0:0] sel);
    case (sel) 0: mux_24877 = 8'h0; 1: mux_24877 = v_24878;
    endcase
  endfunction
  reg [7:0] v_24878 = 8'h0;
  wire [7:0] v_24879;
  wire [7:0] v_24880;
  function [7:0] mux_24880(input [0:0] sel);
    case (sel) 0: mux_24880 = 8'h0; 1: mux_24880 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24881;
  wire [7:0] v_24882;
  wire [7:0] v_24883;
  function [7:0] mux_24883(input [0:0] sel);
    case (sel) 0: mux_24883 = 8'h0; 1: mux_24883 = v_24884;
    endcase
  endfunction
  reg [7:0] v_24884 = 8'h0;
  wire [7:0] v_24885;
  wire [7:0] v_24886;
  function [7:0] mux_24886(input [0:0] sel);
    case (sel) 0: mux_24886 = 8'h0; 1: mux_24886 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24887;
  wire [7:0] v_24888;
  wire [7:0] v_24889;
  function [7:0] mux_24889(input [0:0] sel);
    case (sel) 0: mux_24889 = 8'h0; 1: mux_24889 = vout_peek_12379;
    endcase
  endfunction
  wire [7:0] v_24890;
  function [7:0] mux_24890(input [0:0] sel);
    case (sel) 0: mux_24890 = 8'h0; 1: mux_24890 = vout_peek_12370;
    endcase
  endfunction
  wire [7:0] v_24891;
  function [7:0] mux_24891(input [0:0] sel);
    case (sel) 0: mux_24891 = 8'h0; 1: mux_24891 = v_24892;
    endcase
  endfunction
  reg [7:0] v_24892 = 8'h0;
  wire [7:0] v_24893;
  wire [7:0] v_24894;
  function [7:0] mux_24894(input [0:0] sel);
    case (sel) 0: mux_24894 = 8'h0; 1: mux_24894 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24895;
  wire [7:0] v_24896;
  wire [7:0] v_24897;
  function [7:0] mux_24897(input [0:0] sel);
    case (sel) 0: mux_24897 = 8'h0; 1: mux_24897 = vout_peek_12342;
    endcase
  endfunction
  wire [7:0] v_24898;
  function [7:0] mux_24898(input [0:0] sel);
    case (sel) 0: mux_24898 = 8'h0; 1: mux_24898 = vout_peek_12333;
    endcase
  endfunction
  wire [7:0] v_24899;
  function [7:0] mux_24899(input [0:0] sel);
    case (sel) 0: mux_24899 = 8'h0; 1: mux_24899 = v_24900;
    endcase
  endfunction
  reg [7:0] v_24900 = 8'h0;
  wire [7:0] v_24901;
  wire [7:0] v_24902;
  function [7:0] mux_24902(input [0:0] sel);
    case (sel) 0: mux_24902 = 8'h0; 1: mux_24902 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24903;
  wire [7:0] v_24904;
  wire [7:0] v_24905;
  function [7:0] mux_24905(input [0:0] sel);
    case (sel) 0: mux_24905 = 8'h0; 1: mux_24905 = v_24906;
    endcase
  endfunction
  reg [7:0] v_24906 = 8'h0;
  wire [7:0] v_24907;
  wire [7:0] v_24908;
  function [7:0] mux_24908(input [0:0] sel);
    case (sel) 0: mux_24908 = 8'h0; 1: mux_24908 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24909;
  wire [7:0] v_24910;
  wire [7:0] v_24911;
  function [7:0] mux_24911(input [0:0] sel);
    case (sel) 0: mux_24911 = 8'h0; 1: mux_24911 = vout_peek_12286;
    endcase
  endfunction
  wire [7:0] v_24912;
  function [7:0] mux_24912(input [0:0] sel);
    case (sel) 0: mux_24912 = 8'h0; 1: mux_24912 = vout_peek_12277;
    endcase
  endfunction
  wire [7:0] v_24913;
  function [7:0] mux_24913(input [0:0] sel);
    case (sel) 0: mux_24913 = 8'h0; 1: mux_24913 = v_24914;
    endcase
  endfunction
  reg [7:0] v_24914 = 8'h0;
  wire [7:0] v_24915;
  wire [7:0] v_24916;
  function [7:0] mux_24916(input [0:0] sel);
    case (sel) 0: mux_24916 = 8'h0; 1: mux_24916 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24917;
  wire [7:0] v_24918;
  wire [7:0] v_24919;
  function [7:0] mux_24919(input [0:0] sel);
    case (sel) 0: mux_24919 = 8'h0; 1: mux_24919 = vout_peek_12249;
    endcase
  endfunction
  wire [7:0] v_24920;
  function [7:0] mux_24920(input [0:0] sel);
    case (sel) 0: mux_24920 = 8'h0; 1: mux_24920 = vout_peek_12240;
    endcase
  endfunction
  wire [7:0] v_24921;
  function [7:0] mux_24921(input [0:0] sel);
    case (sel) 0: mux_24921 = 8'h0; 1: mux_24921 = v_24922;
    endcase
  endfunction
  reg [7:0] v_24922 = 8'h0;
  wire [7:0] v_24923;
  wire [7:0] v_24924;
  function [7:0] mux_24924(input [0:0] sel);
    case (sel) 0: mux_24924 = 8'h0; 1: mux_24924 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24925;
  wire [7:0] v_24926;
  wire [7:0] v_24927;
  function [7:0] mux_24927(input [0:0] sel);
    case (sel) 0: mux_24927 = 8'h0; 1: mux_24927 = v_24928;
    endcase
  endfunction
  reg [7:0] v_24928 = 8'h0;
  wire [7:0] v_24929;
  wire [7:0] v_24930;
  function [7:0] mux_24930(input [0:0] sel);
    case (sel) 0: mux_24930 = 8'h0; 1: mux_24930 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24931;
  wire [7:0] v_24932;
  wire [7:0] v_24933;
  function [7:0] mux_24933(input [0:0] sel);
    case (sel) 0: mux_24933 = 8'h0; 1: mux_24933 = v_24934;
    endcase
  endfunction
  reg [7:0] v_24934 = 8'h0;
  wire [7:0] v_24935;
  wire [7:0] v_24936;
  function [7:0] mux_24936(input [0:0] sel);
    case (sel) 0: mux_24936 = 8'h0; 1: mux_24936 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24937;
  wire [7:0] v_24938;
  wire [7:0] v_24939;
  function [7:0] mux_24939(input [0:0] sel);
    case (sel) 0: mux_24939 = 8'h0; 1: mux_24939 = vout_peek_12174;
    endcase
  endfunction
  wire [7:0] v_24940;
  function [7:0] mux_24940(input [0:0] sel);
    case (sel) 0: mux_24940 = 8'h0; 1: mux_24940 = vout_peek_12165;
    endcase
  endfunction
  wire [7:0] v_24941;
  function [7:0] mux_24941(input [0:0] sel);
    case (sel) 0: mux_24941 = 8'h0; 1: mux_24941 = v_24942;
    endcase
  endfunction
  reg [7:0] v_24942 = 8'h0;
  wire [7:0] v_24943;
  wire [7:0] v_24944;
  function [7:0] mux_24944(input [0:0] sel);
    case (sel) 0: mux_24944 = 8'h0; 1: mux_24944 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24945;
  wire [7:0] v_24946;
  wire [7:0] v_24947;
  function [7:0] mux_24947(input [0:0] sel);
    case (sel) 0: mux_24947 = 8'h0; 1: mux_24947 = vout_peek_12137;
    endcase
  endfunction
  wire [7:0] v_24948;
  function [7:0] mux_24948(input [0:0] sel);
    case (sel) 0: mux_24948 = 8'h0; 1: mux_24948 = vout_peek_12128;
    endcase
  endfunction
  wire [7:0] v_24949;
  function [7:0] mux_24949(input [0:0] sel);
    case (sel) 0: mux_24949 = 8'h0; 1: mux_24949 = v_24950;
    endcase
  endfunction
  reg [7:0] v_24950 = 8'h0;
  wire [7:0] v_24951;
  wire [7:0] v_24952;
  function [7:0] mux_24952(input [0:0] sel);
    case (sel) 0: mux_24952 = 8'h0; 1: mux_24952 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24953;
  wire [7:0] v_24954;
  wire [7:0] v_24955;
  function [7:0] mux_24955(input [0:0] sel);
    case (sel) 0: mux_24955 = 8'h0; 1: mux_24955 = v_24956;
    endcase
  endfunction
  reg [7:0] v_24956 = 8'h0;
  wire [7:0] v_24957;
  wire [7:0] v_24958;
  function [7:0] mux_24958(input [0:0] sel);
    case (sel) 0: mux_24958 = 8'h0; 1: mux_24958 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24959;
  wire [7:0] v_24960;
  wire [7:0] v_24961;
  function [7:0] mux_24961(input [0:0] sel);
    case (sel) 0: mux_24961 = 8'h0; 1: mux_24961 = vout_peek_12081;
    endcase
  endfunction
  wire [7:0] v_24962;
  function [7:0] mux_24962(input [0:0] sel);
    case (sel) 0: mux_24962 = 8'h0; 1: mux_24962 = vout_peek_12072;
    endcase
  endfunction
  wire [7:0] v_24963;
  function [7:0] mux_24963(input [0:0] sel);
    case (sel) 0: mux_24963 = 8'h0; 1: mux_24963 = v_24964;
    endcase
  endfunction
  reg [7:0] v_24964 = 8'h0;
  wire [7:0] v_24965;
  wire [7:0] v_24966;
  function [7:0] mux_24966(input [0:0] sel);
    case (sel) 0: mux_24966 = 8'h0; 1: mux_24966 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24967;
  wire [7:0] v_24968;
  wire [7:0] v_24969;
  function [7:0] mux_24969(input [0:0] sel);
    case (sel) 0: mux_24969 = 8'h0; 1: mux_24969 = vout_peek_12044;
    endcase
  endfunction
  wire [7:0] v_24970;
  function [7:0] mux_24970(input [0:0] sel);
    case (sel) 0: mux_24970 = 8'h0; 1: mux_24970 = vout_peek_12035;
    endcase
  endfunction
  wire [7:0] v_24971;
  function [7:0] mux_24971(input [0:0] sel);
    case (sel) 0: mux_24971 = 8'h0; 1: mux_24971 = v_24972;
    endcase
  endfunction
  reg [7:0] v_24972 = 8'h0;
  wire [7:0] v_24973;
  wire [7:0] v_24974;
  function [7:0] mux_24974(input [0:0] sel);
    case (sel) 0: mux_24974 = 8'h0; 1: mux_24974 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24975;
  wire [7:0] v_24976;
  wire [7:0] v_24977;
  function [7:0] mux_24977(input [0:0] sel);
    case (sel) 0: mux_24977 = 8'h0; 1: mux_24977 = v_24978;
    endcase
  endfunction
  reg [7:0] v_24978 = 8'h0;
  wire [7:0] v_24979;
  wire [7:0] v_24980;
  function [7:0] mux_24980(input [0:0] sel);
    case (sel) 0: mux_24980 = 8'h0; 1: mux_24980 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24981;
  wire [7:0] v_24982;
  wire [7:0] v_24983;
  function [7:0] mux_24983(input [0:0] sel);
    case (sel) 0: mux_24983 = 8'h0; 1: mux_24983 = v_24984;
    endcase
  endfunction
  reg [7:0] v_24984 = 8'h0;
  wire [7:0] v_24985;
  wire [7:0] v_24986;
  function [7:0] mux_24986(input [0:0] sel);
    case (sel) 0: mux_24986 = 8'h0; 1: mux_24986 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24987;
  wire [7:0] v_24988;
  wire [7:0] v_24989;
  function [7:0] mux_24989(input [0:0] sel);
    case (sel) 0: mux_24989 = 8'h0; 1: mux_24989 = v_24990;
    endcase
  endfunction
  reg [7:0] v_24990 = 8'h0;
  wire [7:0] v_24991;
  wire [7:0] v_24992;
  function [7:0] mux_24992(input [0:0] sel);
    case (sel) 0: mux_24992 = 8'h0; 1: mux_24992 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_24993;
  wire [7:0] v_24994;
  wire [7:0] v_24995;
  function [7:0] mux_24995(input [0:0] sel);
    case (sel) 0: mux_24995 = 8'h0; 1: mux_24995 = vout_peek_11950;
    endcase
  endfunction
  wire [7:0] v_24996;
  function [7:0] mux_24996(input [0:0] sel);
    case (sel) 0: mux_24996 = 8'h0; 1: mux_24996 = vout_peek_11941;
    endcase
  endfunction
  wire [7:0] v_24997;
  function [7:0] mux_24997(input [0:0] sel);
    case (sel) 0: mux_24997 = 8'h0; 1: mux_24997 = v_24998;
    endcase
  endfunction
  reg [7:0] v_24998 = 8'h0;
  wire [7:0] v_24999;
  wire [7:0] v_25000;
  function [7:0] mux_25000(input [0:0] sel);
    case (sel) 0: mux_25000 = 8'h0; 1: mux_25000 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25001;
  wire [7:0] v_25002;
  wire [7:0] v_25003;
  function [7:0] mux_25003(input [0:0] sel);
    case (sel) 0: mux_25003 = 8'h0; 1: mux_25003 = vout_peek_11913;
    endcase
  endfunction
  wire [7:0] v_25004;
  function [7:0] mux_25004(input [0:0] sel);
    case (sel) 0: mux_25004 = 8'h0; 1: mux_25004 = vout_peek_11904;
    endcase
  endfunction
  wire [7:0] v_25005;
  function [7:0] mux_25005(input [0:0] sel);
    case (sel) 0: mux_25005 = 8'h0; 1: mux_25005 = v_25006;
    endcase
  endfunction
  reg [7:0] v_25006 = 8'h0;
  wire [7:0] v_25007;
  wire [7:0] v_25008;
  function [7:0] mux_25008(input [0:0] sel);
    case (sel) 0: mux_25008 = 8'h0; 1: mux_25008 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25009;
  wire [7:0] v_25010;
  wire [7:0] v_25011;
  function [7:0] mux_25011(input [0:0] sel);
    case (sel) 0: mux_25011 = 8'h0; 1: mux_25011 = v_25012;
    endcase
  endfunction
  reg [7:0] v_25012 = 8'h0;
  wire [7:0] v_25013;
  wire [7:0] v_25014;
  function [7:0] mux_25014(input [0:0] sel);
    case (sel) 0: mux_25014 = 8'h0; 1: mux_25014 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25015;
  wire [7:0] v_25016;
  wire [7:0] v_25017;
  function [7:0] mux_25017(input [0:0] sel);
    case (sel) 0: mux_25017 = 8'h0; 1: mux_25017 = vout_peek_11857;
    endcase
  endfunction
  wire [7:0] v_25018;
  function [7:0] mux_25018(input [0:0] sel);
    case (sel) 0: mux_25018 = 8'h0; 1: mux_25018 = vout_peek_11848;
    endcase
  endfunction
  wire [7:0] v_25019;
  function [7:0] mux_25019(input [0:0] sel);
    case (sel) 0: mux_25019 = 8'h0; 1: mux_25019 = v_25020;
    endcase
  endfunction
  reg [7:0] v_25020 = 8'h0;
  wire [7:0] v_25021;
  wire [7:0] v_25022;
  function [7:0] mux_25022(input [0:0] sel);
    case (sel) 0: mux_25022 = 8'h0; 1: mux_25022 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25023;
  wire [7:0] v_25024;
  wire [7:0] v_25025;
  function [7:0] mux_25025(input [0:0] sel);
    case (sel) 0: mux_25025 = 8'h0; 1: mux_25025 = vout_peek_11820;
    endcase
  endfunction
  wire [7:0] v_25026;
  function [7:0] mux_25026(input [0:0] sel);
    case (sel) 0: mux_25026 = 8'h0; 1: mux_25026 = vout_peek_11811;
    endcase
  endfunction
  wire [7:0] v_25027;
  function [7:0] mux_25027(input [0:0] sel);
    case (sel) 0: mux_25027 = 8'h0; 1: mux_25027 = v_25028;
    endcase
  endfunction
  reg [7:0] v_25028 = 8'h0;
  wire [7:0] v_25029;
  wire [7:0] v_25030;
  function [7:0] mux_25030(input [0:0] sel);
    case (sel) 0: mux_25030 = 8'h0; 1: mux_25030 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25031;
  wire [7:0] v_25032;
  wire [7:0] v_25033;
  function [7:0] mux_25033(input [0:0] sel);
    case (sel) 0: mux_25033 = 8'h0; 1: mux_25033 = v_25034;
    endcase
  endfunction
  reg [7:0] v_25034 = 8'h0;
  wire [7:0] v_25035;
  wire [7:0] v_25036;
  function [7:0] mux_25036(input [0:0] sel);
    case (sel) 0: mux_25036 = 8'h0; 1: mux_25036 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25037;
  wire [7:0] v_25038;
  wire [7:0] v_25039;
  function [7:0] mux_25039(input [0:0] sel);
    case (sel) 0: mux_25039 = 8'h0; 1: mux_25039 = v_25040;
    endcase
  endfunction
  reg [7:0] v_25040 = 8'h0;
  wire [7:0] v_25041;
  wire [7:0] v_25042;
  function [7:0] mux_25042(input [0:0] sel);
    case (sel) 0: mux_25042 = 8'h0; 1: mux_25042 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25043;
  wire [7:0] v_25044;
  wire [7:0] v_25045;
  function [7:0] mux_25045(input [0:0] sel);
    case (sel) 0: mux_25045 = 8'h0; 1: mux_25045 = vout_peek_11745;
    endcase
  endfunction
  wire [7:0] v_25046;
  function [7:0] mux_25046(input [0:0] sel);
    case (sel) 0: mux_25046 = 8'h0; 1: mux_25046 = vout_peek_11736;
    endcase
  endfunction
  wire [7:0] v_25047;
  function [7:0] mux_25047(input [0:0] sel);
    case (sel) 0: mux_25047 = 8'h0; 1: mux_25047 = v_25048;
    endcase
  endfunction
  reg [7:0] v_25048 = 8'h0;
  wire [7:0] v_25049;
  wire [7:0] v_25050;
  function [7:0] mux_25050(input [0:0] sel);
    case (sel) 0: mux_25050 = 8'h0; 1: mux_25050 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25051;
  wire [7:0] v_25052;
  wire [7:0] v_25053;
  function [7:0] mux_25053(input [0:0] sel);
    case (sel) 0: mux_25053 = 8'h0; 1: mux_25053 = vout_peek_11708;
    endcase
  endfunction
  wire [7:0] v_25054;
  function [7:0] mux_25054(input [0:0] sel);
    case (sel) 0: mux_25054 = 8'h0; 1: mux_25054 = vout_peek_11699;
    endcase
  endfunction
  wire [7:0] v_25055;
  function [7:0] mux_25055(input [0:0] sel);
    case (sel) 0: mux_25055 = 8'h0; 1: mux_25055 = v_25056;
    endcase
  endfunction
  reg [7:0] v_25056 = 8'h0;
  wire [7:0] v_25057;
  wire [7:0] v_25058;
  function [7:0] mux_25058(input [0:0] sel);
    case (sel) 0: mux_25058 = 8'h0; 1: mux_25058 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25059;
  wire [7:0] v_25060;
  wire [7:0] v_25061;
  function [7:0] mux_25061(input [0:0] sel);
    case (sel) 0: mux_25061 = 8'h0; 1: mux_25061 = v_25062;
    endcase
  endfunction
  reg [7:0] v_25062 = 8'h0;
  wire [7:0] v_25063;
  wire [7:0] v_25064;
  function [7:0] mux_25064(input [0:0] sel);
    case (sel) 0: mux_25064 = 8'h0; 1: mux_25064 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25065;
  wire [7:0] v_25066;
  wire [7:0] v_25067;
  function [7:0] mux_25067(input [0:0] sel);
    case (sel) 0: mux_25067 = 8'h0; 1: mux_25067 = vout_peek_11652;
    endcase
  endfunction
  wire [7:0] v_25068;
  function [7:0] mux_25068(input [0:0] sel);
    case (sel) 0: mux_25068 = 8'h0; 1: mux_25068 = vout_peek_11643;
    endcase
  endfunction
  wire [7:0] v_25069;
  function [7:0] mux_25069(input [0:0] sel);
    case (sel) 0: mux_25069 = 8'h0; 1: mux_25069 = v_25070;
    endcase
  endfunction
  reg [7:0] v_25070 = 8'h0;
  wire [7:0] v_25071;
  wire [7:0] v_25072;
  function [7:0] mux_25072(input [0:0] sel);
    case (sel) 0: mux_25072 = 8'h0; 1: mux_25072 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25073;
  wire [7:0] v_25074;
  wire [7:0] v_25075;
  function [7:0] mux_25075(input [0:0] sel);
    case (sel) 0: mux_25075 = 8'h0; 1: mux_25075 = vout_peek_11615;
    endcase
  endfunction
  wire [7:0] v_25076;
  function [7:0] mux_25076(input [0:0] sel);
    case (sel) 0: mux_25076 = 8'h0; 1: mux_25076 = vout_peek_11606;
    endcase
  endfunction
  wire [7:0] v_25077;
  function [7:0] mux_25077(input [0:0] sel);
    case (sel) 0: mux_25077 = 8'h0; 1: mux_25077 = v_25078;
    endcase
  endfunction
  reg [7:0] v_25078 = 8'h0;
  wire [7:0] v_25079;
  wire [7:0] v_25080;
  function [7:0] mux_25080(input [0:0] sel);
    case (sel) 0: mux_25080 = 8'h0; 1: mux_25080 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25081;
  wire [7:0] v_25082;
  wire [7:0] v_25083;
  function [7:0] mux_25083(input [0:0] sel);
    case (sel) 0: mux_25083 = 8'h0; 1: mux_25083 = v_25084;
    endcase
  endfunction
  reg [7:0] v_25084 = 8'h0;
  wire [7:0] v_25085;
  wire [7:0] v_25086;
  function [7:0] mux_25086(input [0:0] sel);
    case (sel) 0: mux_25086 = 8'h0; 1: mux_25086 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25087;
  wire [7:0] v_25088;
  wire [7:0] v_25089;
  function [7:0] mux_25089(input [0:0] sel);
    case (sel) 0: mux_25089 = 8'h0; 1: mux_25089 = v_25090;
    endcase
  endfunction
  reg [7:0] v_25090 = 8'h0;
  wire [7:0] v_25091;
  wire [7:0] v_25092;
  function [7:0] mux_25092(input [0:0] sel);
    case (sel) 0: mux_25092 = 8'h0; 1: mux_25092 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25093;
  wire [7:0] v_25094;
  wire [7:0] v_25095;
  function [7:0] mux_25095(input [0:0] sel);
    case (sel) 0: mux_25095 = 8'h0; 1: mux_25095 = v_25096;
    endcase
  endfunction
  reg [7:0] v_25096 = 8'h0;
  wire [7:0] v_25097;
  wire [7:0] v_25098;
  function [7:0] mux_25098(input [0:0] sel);
    case (sel) 0: mux_25098 = 8'h0; 1: mux_25098 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25099;
  wire [7:0] v_25100;
  wire [7:0] v_25101;
  function [7:0] mux_25101(input [0:0] sel);
    case (sel) 0: mux_25101 = 8'h0; 1: mux_25101 = v_25102;
    endcase
  endfunction
  reg [7:0] v_25102 = 8'h0;
  wire [7:0] v_25103;
  wire [7:0] v_25104;
  function [7:0] mux_25104(input [0:0] sel);
    case (sel) 0: mux_25104 = 8'h0; 1: mux_25104 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25105;
  wire [7:0] v_25106;
  wire [7:0] v_25107;
  function [7:0] mux_25107(input [0:0] sel);
    case (sel) 0: mux_25107 = 8'h0; 1: mux_25107 = v_25108;
    endcase
  endfunction
  reg [7:0] v_25108 = 8'h0;
  wire [7:0] v_25109;
  wire [7:0] v_25110;
  function [7:0] mux_25110(input [0:0] sel);
    case (sel) 0: mux_25110 = 8'h0; 1: mux_25110 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25111;
  wire [7:0] v_25112;
  wire [7:0] v_25113;
  function [7:0] mux_25113(input [0:0] sel);
    case (sel) 0: mux_25113 = 8'h0; 1: mux_25113 = v_25114;
    endcase
  endfunction
  reg [7:0] v_25114 = 8'h0;
  wire [7:0] v_25115;
  wire [7:0] v_25116;
  function [7:0] mux_25116(input [0:0] sel);
    case (sel) 0: mux_25116 = 8'h0; 1: mux_25116 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25117;
  wire [7:0] v_25118;
  wire [7:0] v_25119;
  function [7:0] mux_25119(input [0:0] sel);
    case (sel) 0: mux_25119 = 8'h0; 1: mux_25119 = vout_peek_11464;
    endcase
  endfunction
  wire [7:0] v_25120;
  function [7:0] mux_25120(input [0:0] sel);
    case (sel) 0: mux_25120 = 8'h0; 1: mux_25120 = vout_peek_11455;
    endcase
  endfunction
  wire [7:0] v_25121;
  function [7:0] mux_25121(input [0:0] sel);
    case (sel) 0: mux_25121 = 8'h0; 1: mux_25121 = v_25122;
    endcase
  endfunction
  reg [7:0] v_25122 = 8'h0;
  wire [7:0] v_25123;
  wire [7:0] v_25124;
  function [7:0] mux_25124(input [0:0] sel);
    case (sel) 0: mux_25124 = 8'h0; 1: mux_25124 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25125;
  wire [7:0] v_25126;
  wire [7:0] v_25127;
  function [7:0] mux_25127(input [0:0] sel);
    case (sel) 0: mux_25127 = 8'h0; 1: mux_25127 = vout_peek_11427;
    endcase
  endfunction
  wire [7:0] v_25128;
  function [7:0] mux_25128(input [0:0] sel);
    case (sel) 0: mux_25128 = 8'h0; 1: mux_25128 = vout_peek_11418;
    endcase
  endfunction
  wire [7:0] v_25129;
  function [7:0] mux_25129(input [0:0] sel);
    case (sel) 0: mux_25129 = 8'h0; 1: mux_25129 = v_25130;
    endcase
  endfunction
  reg [7:0] v_25130 = 8'h0;
  wire [7:0] v_25131;
  wire [7:0] v_25132;
  function [7:0] mux_25132(input [0:0] sel);
    case (sel) 0: mux_25132 = 8'h0; 1: mux_25132 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25133;
  wire [7:0] v_25134;
  wire [7:0] v_25135;
  function [7:0] mux_25135(input [0:0] sel);
    case (sel) 0: mux_25135 = 8'h0; 1: mux_25135 = v_25136;
    endcase
  endfunction
  reg [7:0] v_25136 = 8'h0;
  wire [7:0] v_25137;
  wire [7:0] v_25138;
  function [7:0] mux_25138(input [0:0] sel);
    case (sel) 0: mux_25138 = 8'h0; 1: mux_25138 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25139;
  wire [7:0] v_25140;
  wire [7:0] v_25141;
  function [7:0] mux_25141(input [0:0] sel);
    case (sel) 0: mux_25141 = 8'h0; 1: mux_25141 = vout_peek_11371;
    endcase
  endfunction
  wire [7:0] v_25142;
  function [7:0] mux_25142(input [0:0] sel);
    case (sel) 0: mux_25142 = 8'h0; 1: mux_25142 = vout_peek_11362;
    endcase
  endfunction
  wire [7:0] v_25143;
  function [7:0] mux_25143(input [0:0] sel);
    case (sel) 0: mux_25143 = 8'h0; 1: mux_25143 = v_25144;
    endcase
  endfunction
  reg [7:0] v_25144 = 8'h0;
  wire [7:0] v_25145;
  wire [7:0] v_25146;
  function [7:0] mux_25146(input [0:0] sel);
    case (sel) 0: mux_25146 = 8'h0; 1: mux_25146 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25147;
  wire [7:0] v_25148;
  wire [7:0] v_25149;
  function [7:0] mux_25149(input [0:0] sel);
    case (sel) 0: mux_25149 = 8'h0; 1: mux_25149 = vout_peek_11334;
    endcase
  endfunction
  wire [7:0] v_25150;
  function [7:0] mux_25150(input [0:0] sel);
    case (sel) 0: mux_25150 = 8'h0; 1: mux_25150 = vout_peek_11325;
    endcase
  endfunction
  wire [7:0] v_25151;
  function [7:0] mux_25151(input [0:0] sel);
    case (sel) 0: mux_25151 = 8'h0; 1: mux_25151 = v_25152;
    endcase
  endfunction
  reg [7:0] v_25152 = 8'h0;
  wire [7:0] v_25153;
  wire [7:0] v_25154;
  function [7:0] mux_25154(input [0:0] sel);
    case (sel) 0: mux_25154 = 8'h0; 1: mux_25154 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25155;
  wire [7:0] v_25156;
  wire [7:0] v_25157;
  function [7:0] mux_25157(input [0:0] sel);
    case (sel) 0: mux_25157 = 8'h0; 1: mux_25157 = v_25158;
    endcase
  endfunction
  reg [7:0] v_25158 = 8'h0;
  wire [7:0] v_25159;
  wire [7:0] v_25160;
  function [7:0] mux_25160(input [0:0] sel);
    case (sel) 0: mux_25160 = 8'h0; 1: mux_25160 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25161;
  wire [7:0] v_25162;
  wire [7:0] v_25163;
  function [7:0] mux_25163(input [0:0] sel);
    case (sel) 0: mux_25163 = 8'h0; 1: mux_25163 = v_25164;
    endcase
  endfunction
  reg [7:0] v_25164 = 8'h0;
  wire [7:0] v_25165;
  wire [7:0] v_25166;
  function [7:0] mux_25166(input [0:0] sel);
    case (sel) 0: mux_25166 = 8'h0; 1: mux_25166 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25167;
  wire [7:0] v_25168;
  wire [7:0] v_25169;
  function [7:0] mux_25169(input [0:0] sel);
    case (sel) 0: mux_25169 = 8'h0; 1: mux_25169 = vout_peek_11259;
    endcase
  endfunction
  wire [7:0] v_25170;
  function [7:0] mux_25170(input [0:0] sel);
    case (sel) 0: mux_25170 = 8'h0; 1: mux_25170 = vout_peek_11250;
    endcase
  endfunction
  wire [7:0] v_25171;
  function [7:0] mux_25171(input [0:0] sel);
    case (sel) 0: mux_25171 = 8'h0; 1: mux_25171 = v_25172;
    endcase
  endfunction
  reg [7:0] v_25172 = 8'h0;
  wire [7:0] v_25173;
  wire [7:0] v_25174;
  function [7:0] mux_25174(input [0:0] sel);
    case (sel) 0: mux_25174 = 8'h0; 1: mux_25174 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25175;
  wire [7:0] v_25176;
  wire [7:0] v_25177;
  function [7:0] mux_25177(input [0:0] sel);
    case (sel) 0: mux_25177 = 8'h0; 1: mux_25177 = vout_peek_11222;
    endcase
  endfunction
  wire [7:0] v_25178;
  function [7:0] mux_25178(input [0:0] sel);
    case (sel) 0: mux_25178 = 8'h0; 1: mux_25178 = vout_peek_11213;
    endcase
  endfunction
  wire [7:0] v_25179;
  function [7:0] mux_25179(input [0:0] sel);
    case (sel) 0: mux_25179 = 8'h0; 1: mux_25179 = v_25180;
    endcase
  endfunction
  reg [7:0] v_25180 = 8'h0;
  wire [7:0] v_25181;
  wire [7:0] v_25182;
  function [7:0] mux_25182(input [0:0] sel);
    case (sel) 0: mux_25182 = 8'h0; 1: mux_25182 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25183;
  wire [7:0] v_25184;
  wire [7:0] v_25185;
  function [7:0] mux_25185(input [0:0] sel);
    case (sel) 0: mux_25185 = 8'h0; 1: mux_25185 = v_25186;
    endcase
  endfunction
  reg [7:0] v_25186 = 8'h0;
  wire [7:0] v_25187;
  wire [7:0] v_25188;
  function [7:0] mux_25188(input [0:0] sel);
    case (sel) 0: mux_25188 = 8'h0; 1: mux_25188 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25189;
  wire [7:0] v_25190;
  wire [7:0] v_25191;
  function [7:0] mux_25191(input [0:0] sel);
    case (sel) 0: mux_25191 = 8'h0; 1: mux_25191 = vout_peek_11166;
    endcase
  endfunction
  wire [7:0] v_25192;
  function [7:0] mux_25192(input [0:0] sel);
    case (sel) 0: mux_25192 = 8'h0; 1: mux_25192 = vout_peek_11157;
    endcase
  endfunction
  wire [7:0] v_25193;
  function [7:0] mux_25193(input [0:0] sel);
    case (sel) 0: mux_25193 = 8'h0; 1: mux_25193 = v_25194;
    endcase
  endfunction
  reg [7:0] v_25194 = 8'h0;
  wire [7:0] v_25195;
  wire [7:0] v_25196;
  function [7:0] mux_25196(input [0:0] sel);
    case (sel) 0: mux_25196 = 8'h0; 1: mux_25196 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25197;
  wire [7:0] v_25198;
  wire [7:0] v_25199;
  function [7:0] mux_25199(input [0:0] sel);
    case (sel) 0: mux_25199 = 8'h0; 1: mux_25199 = vout_peek_11129;
    endcase
  endfunction
  wire [7:0] v_25200;
  function [7:0] mux_25200(input [0:0] sel);
    case (sel) 0: mux_25200 = 8'h0; 1: mux_25200 = vout_peek_11120;
    endcase
  endfunction
  wire [7:0] v_25201;
  function [7:0] mux_25201(input [0:0] sel);
    case (sel) 0: mux_25201 = 8'h0; 1: mux_25201 = v_25202;
    endcase
  endfunction
  reg [7:0] v_25202 = 8'h0;
  wire [7:0] v_25203;
  wire [7:0] v_25204;
  function [7:0] mux_25204(input [0:0] sel);
    case (sel) 0: mux_25204 = 8'h0; 1: mux_25204 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25205;
  wire [7:0] v_25206;
  wire [7:0] v_25207;
  function [7:0] mux_25207(input [0:0] sel);
    case (sel) 0: mux_25207 = 8'h0; 1: mux_25207 = v_25208;
    endcase
  endfunction
  reg [7:0] v_25208 = 8'h0;
  wire [7:0] v_25209;
  wire [7:0] v_25210;
  function [7:0] mux_25210(input [0:0] sel);
    case (sel) 0: mux_25210 = 8'h0; 1: mux_25210 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25211;
  wire [7:0] v_25212;
  wire [7:0] v_25213;
  function [7:0] mux_25213(input [0:0] sel);
    case (sel) 0: mux_25213 = 8'h0; 1: mux_25213 = v_25214;
    endcase
  endfunction
  reg [7:0] v_25214 = 8'h0;
  wire [7:0] v_25215;
  wire [7:0] v_25216;
  function [7:0] mux_25216(input [0:0] sel);
    case (sel) 0: mux_25216 = 8'h0; 1: mux_25216 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25217;
  wire [7:0] v_25218;
  wire [7:0] v_25219;
  function [7:0] mux_25219(input [0:0] sel);
    case (sel) 0: mux_25219 = 8'h0; 1: mux_25219 = v_25220;
    endcase
  endfunction
  reg [7:0] v_25220 = 8'h0;
  wire [7:0] v_25221;
  wire [7:0] v_25222;
  function [7:0] mux_25222(input [0:0] sel);
    case (sel) 0: mux_25222 = 8'h0; 1: mux_25222 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25223;
  wire [7:0] v_25224;
  wire [7:0] v_25225;
  function [7:0] mux_25225(input [0:0] sel);
    case (sel) 0: mux_25225 = 8'h0; 1: mux_25225 = vout_peek_11035;
    endcase
  endfunction
  wire [7:0] v_25226;
  function [7:0] mux_25226(input [0:0] sel);
    case (sel) 0: mux_25226 = 8'h0; 1: mux_25226 = vout_peek_11026;
    endcase
  endfunction
  wire [7:0] v_25227;
  function [7:0] mux_25227(input [0:0] sel);
    case (sel) 0: mux_25227 = 8'h0; 1: mux_25227 = v_25228;
    endcase
  endfunction
  reg [7:0] v_25228 = 8'h0;
  wire [7:0] v_25229;
  wire [7:0] v_25230;
  function [7:0] mux_25230(input [0:0] sel);
    case (sel) 0: mux_25230 = 8'h0; 1: mux_25230 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25231;
  wire [7:0] v_25232;
  wire [7:0] v_25233;
  function [7:0] mux_25233(input [0:0] sel);
    case (sel) 0: mux_25233 = 8'h0; 1: mux_25233 = vout_peek_10998;
    endcase
  endfunction
  wire [7:0] v_25234;
  function [7:0] mux_25234(input [0:0] sel);
    case (sel) 0: mux_25234 = 8'h0; 1: mux_25234 = vout_peek_10989;
    endcase
  endfunction
  wire [7:0] v_25235;
  function [7:0] mux_25235(input [0:0] sel);
    case (sel) 0: mux_25235 = 8'h0; 1: mux_25235 = v_25236;
    endcase
  endfunction
  reg [7:0] v_25236 = 8'h0;
  wire [7:0] v_25237;
  wire [7:0] v_25238;
  function [7:0] mux_25238(input [0:0] sel);
    case (sel) 0: mux_25238 = 8'h0; 1: mux_25238 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25239;
  wire [7:0] v_25240;
  wire [7:0] v_25241;
  function [7:0] mux_25241(input [0:0] sel);
    case (sel) 0: mux_25241 = 8'h0; 1: mux_25241 = v_25242;
    endcase
  endfunction
  reg [7:0] v_25242 = 8'h0;
  wire [7:0] v_25243;
  wire [7:0] v_25244;
  function [7:0] mux_25244(input [0:0] sel);
    case (sel) 0: mux_25244 = 8'h0; 1: mux_25244 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25245;
  wire [7:0] v_25246;
  wire [7:0] v_25247;
  function [7:0] mux_25247(input [0:0] sel);
    case (sel) 0: mux_25247 = 8'h0; 1: mux_25247 = vout_peek_10942;
    endcase
  endfunction
  wire [7:0] v_25248;
  function [7:0] mux_25248(input [0:0] sel);
    case (sel) 0: mux_25248 = 8'h0; 1: mux_25248 = vout_peek_10933;
    endcase
  endfunction
  wire [7:0] v_25249;
  function [7:0] mux_25249(input [0:0] sel);
    case (sel) 0: mux_25249 = 8'h0; 1: mux_25249 = v_25250;
    endcase
  endfunction
  reg [7:0] v_25250 = 8'h0;
  wire [7:0] v_25251;
  wire [7:0] v_25252;
  function [7:0] mux_25252(input [0:0] sel);
    case (sel) 0: mux_25252 = 8'h0; 1: mux_25252 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25253;
  wire [7:0] v_25254;
  wire [7:0] v_25255;
  function [7:0] mux_25255(input [0:0] sel);
    case (sel) 0: mux_25255 = 8'h0; 1: mux_25255 = vout_peek_10905;
    endcase
  endfunction
  wire [7:0] v_25256;
  function [7:0] mux_25256(input [0:0] sel);
    case (sel) 0: mux_25256 = 8'h0; 1: mux_25256 = vout_peek_10896;
    endcase
  endfunction
  wire [7:0] v_25257;
  function [7:0] mux_25257(input [0:0] sel);
    case (sel) 0: mux_25257 = 8'h0; 1: mux_25257 = v_25258;
    endcase
  endfunction
  reg [7:0] v_25258 = 8'h0;
  wire [7:0] v_25259;
  wire [7:0] v_25260;
  function [7:0] mux_25260(input [0:0] sel);
    case (sel) 0: mux_25260 = 8'h0; 1: mux_25260 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25261;
  wire [7:0] v_25262;
  wire [7:0] v_25263;
  function [7:0] mux_25263(input [0:0] sel);
    case (sel) 0: mux_25263 = 8'h0; 1: mux_25263 = v_25264;
    endcase
  endfunction
  reg [7:0] v_25264 = 8'h0;
  wire [7:0] v_25265;
  wire [7:0] v_25266;
  function [7:0] mux_25266(input [0:0] sel);
    case (sel) 0: mux_25266 = 8'h0; 1: mux_25266 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25267;
  wire [7:0] v_25268;
  wire [7:0] v_25269;
  function [7:0] mux_25269(input [0:0] sel);
    case (sel) 0: mux_25269 = 8'h0; 1: mux_25269 = v_25270;
    endcase
  endfunction
  reg [7:0] v_25270 = 8'h0;
  wire [7:0] v_25271;
  wire [7:0] v_25272;
  function [7:0] mux_25272(input [0:0] sel);
    case (sel) 0: mux_25272 = 8'h0; 1: mux_25272 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25273;
  wire [7:0] v_25274;
  wire [7:0] v_25275;
  function [7:0] mux_25275(input [0:0] sel);
    case (sel) 0: mux_25275 = 8'h0; 1: mux_25275 = vout_peek_10830;
    endcase
  endfunction
  wire [7:0] v_25276;
  function [7:0] mux_25276(input [0:0] sel);
    case (sel) 0: mux_25276 = 8'h0; 1: mux_25276 = vout_peek_10821;
    endcase
  endfunction
  wire [7:0] v_25277;
  function [7:0] mux_25277(input [0:0] sel);
    case (sel) 0: mux_25277 = 8'h0; 1: mux_25277 = v_25278;
    endcase
  endfunction
  reg [7:0] v_25278 = 8'h0;
  wire [7:0] v_25279;
  wire [7:0] v_25280;
  function [7:0] mux_25280(input [0:0] sel);
    case (sel) 0: mux_25280 = 8'h0; 1: mux_25280 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25281;
  wire [7:0] v_25282;
  wire [7:0] v_25283;
  function [7:0] mux_25283(input [0:0] sel);
    case (sel) 0: mux_25283 = 8'h0; 1: mux_25283 = vout_peek_10793;
    endcase
  endfunction
  wire [7:0] v_25284;
  function [7:0] mux_25284(input [0:0] sel);
    case (sel) 0: mux_25284 = 8'h0; 1: mux_25284 = vout_peek_10784;
    endcase
  endfunction
  wire [7:0] v_25285;
  function [7:0] mux_25285(input [0:0] sel);
    case (sel) 0: mux_25285 = 8'h0; 1: mux_25285 = v_25286;
    endcase
  endfunction
  reg [7:0] v_25286 = 8'h0;
  wire [7:0] v_25287;
  wire [7:0] v_25288;
  function [7:0] mux_25288(input [0:0] sel);
    case (sel) 0: mux_25288 = 8'h0; 1: mux_25288 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25289;
  wire [7:0] v_25290;
  wire [7:0] v_25291;
  function [7:0] mux_25291(input [0:0] sel);
    case (sel) 0: mux_25291 = 8'h0; 1: mux_25291 = v_25292;
    endcase
  endfunction
  reg [7:0] v_25292 = 8'h0;
  wire [7:0] v_25293;
  wire [7:0] v_25294;
  function [7:0] mux_25294(input [0:0] sel);
    case (sel) 0: mux_25294 = 8'h0; 1: mux_25294 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25295;
  wire [7:0] v_25296;
  wire [7:0] v_25297;
  function [7:0] mux_25297(input [0:0] sel);
    case (sel) 0: mux_25297 = 8'h0; 1: mux_25297 = vout_peek_10737;
    endcase
  endfunction
  wire [7:0] v_25298;
  function [7:0] mux_25298(input [0:0] sel);
    case (sel) 0: mux_25298 = 8'h0; 1: mux_25298 = vout_peek_10728;
    endcase
  endfunction
  wire [7:0] v_25299;
  function [7:0] mux_25299(input [0:0] sel);
    case (sel) 0: mux_25299 = 8'h0; 1: mux_25299 = v_25300;
    endcase
  endfunction
  reg [7:0] v_25300 = 8'h0;
  wire [7:0] v_25301;
  wire [7:0] v_25302;
  function [7:0] mux_25302(input [0:0] sel);
    case (sel) 0: mux_25302 = 8'h0; 1: mux_25302 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25303;
  wire [7:0] v_25304;
  wire [7:0] v_25305;
  function [7:0] mux_25305(input [0:0] sel);
    case (sel) 0: mux_25305 = 8'h0; 1: mux_25305 = vout_peek_10700;
    endcase
  endfunction
  wire [7:0] v_25306;
  function [7:0] mux_25306(input [0:0] sel);
    case (sel) 0: mux_25306 = 8'h0; 1: mux_25306 = vout_peek_10691;
    endcase
  endfunction
  wire [7:0] v_25307;
  function [7:0] mux_25307(input [0:0] sel);
    case (sel) 0: mux_25307 = 8'h0; 1: mux_25307 = v_25308;
    endcase
  endfunction
  reg [7:0] v_25308 = 8'h0;
  wire [7:0] v_25309;
  wire [7:0] v_25310;
  function [7:0] mux_25310(input [0:0] sel);
    case (sel) 0: mux_25310 = 8'h0; 1: mux_25310 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25311;
  wire [7:0] v_25312;
  wire [7:0] v_25313;
  function [7:0] mux_25313(input [0:0] sel);
    case (sel) 0: mux_25313 = 8'h0; 1: mux_25313 = v_25314;
    endcase
  endfunction
  reg [7:0] v_25314 = 8'h0;
  wire [7:0] v_25315;
  wire [7:0] v_25316;
  function [7:0] mux_25316(input [0:0] sel);
    case (sel) 0: mux_25316 = 8'h0; 1: mux_25316 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25317;
  wire [7:0] v_25318;
  wire [7:0] v_25319;
  function [7:0] mux_25319(input [0:0] sel);
    case (sel) 0: mux_25319 = 8'h0; 1: mux_25319 = v_25320;
    endcase
  endfunction
  reg [7:0] v_25320 = 8'h0;
  wire [7:0] v_25321;
  wire [7:0] v_25322;
  function [7:0] mux_25322(input [0:0] sel);
    case (sel) 0: mux_25322 = 8'h0; 1: mux_25322 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25323;
  wire [7:0] v_25324;
  wire [7:0] v_25325;
  function [7:0] mux_25325(input [0:0] sel);
    case (sel) 0: mux_25325 = 8'h0; 1: mux_25325 = v_25326;
    endcase
  endfunction
  reg [7:0] v_25326 = 8'h0;
  wire [7:0] v_25327;
  wire [7:0] v_25328;
  function [7:0] mux_25328(input [0:0] sel);
    case (sel) 0: mux_25328 = 8'h0; 1: mux_25328 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25329;
  wire [7:0] v_25330;
  wire [7:0] v_25331;
  function [7:0] mux_25331(input [0:0] sel);
    case (sel) 0: mux_25331 = 8'h0; 1: mux_25331 = v_25332;
    endcase
  endfunction
  reg [7:0] v_25332 = 8'h0;
  wire [7:0] v_25333;
  wire [7:0] v_25334;
  function [7:0] mux_25334(input [0:0] sel);
    case (sel) 0: mux_25334 = 8'h0; 1: mux_25334 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25335;
  wire [7:0] v_25336;
  wire [7:0] v_25337;
  function [7:0] mux_25337(input [0:0] sel);
    case (sel) 0: mux_25337 = 8'h0; 1: mux_25337 = vout_peek_10587;
    endcase
  endfunction
  wire [7:0] v_25338;
  function [7:0] mux_25338(input [0:0] sel);
    case (sel) 0: mux_25338 = 8'h0; 1: mux_25338 = vout_peek_10578;
    endcase
  endfunction
  wire [7:0] v_25339;
  function [7:0] mux_25339(input [0:0] sel);
    case (sel) 0: mux_25339 = 8'h0; 1: mux_25339 = v_25340;
    endcase
  endfunction
  reg [7:0] v_25340 = 8'h0;
  wire [7:0] v_25341;
  wire [7:0] v_25342;
  function [7:0] mux_25342(input [0:0] sel);
    case (sel) 0: mux_25342 = 8'h0; 1: mux_25342 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25343;
  wire [7:0] v_25344;
  wire [7:0] v_25345;
  function [7:0] mux_25345(input [0:0] sel);
    case (sel) 0: mux_25345 = 8'h0; 1: mux_25345 = vout_peek_10550;
    endcase
  endfunction
  wire [7:0] v_25346;
  function [7:0] mux_25346(input [0:0] sel);
    case (sel) 0: mux_25346 = 8'h0; 1: mux_25346 = vout_peek_10541;
    endcase
  endfunction
  wire [7:0] v_25347;
  function [7:0] mux_25347(input [0:0] sel);
    case (sel) 0: mux_25347 = 8'h0; 1: mux_25347 = v_25348;
    endcase
  endfunction
  reg [7:0] v_25348 = 8'h0;
  wire [7:0] v_25349;
  wire [7:0] v_25350;
  function [7:0] mux_25350(input [0:0] sel);
    case (sel) 0: mux_25350 = 8'h0; 1: mux_25350 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25351;
  wire [7:0] v_25352;
  wire [7:0] v_25353;
  function [7:0] mux_25353(input [0:0] sel);
    case (sel) 0: mux_25353 = 8'h0; 1: mux_25353 = v_25354;
    endcase
  endfunction
  reg [7:0] v_25354 = 8'h0;
  wire [7:0] v_25355;
  wire [7:0] v_25356;
  function [7:0] mux_25356(input [0:0] sel);
    case (sel) 0: mux_25356 = 8'h0; 1: mux_25356 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25357;
  wire [7:0] v_25358;
  wire [7:0] v_25359;
  function [7:0] mux_25359(input [0:0] sel);
    case (sel) 0: mux_25359 = 8'h0; 1: mux_25359 = vout_peek_10494;
    endcase
  endfunction
  wire [7:0] v_25360;
  function [7:0] mux_25360(input [0:0] sel);
    case (sel) 0: mux_25360 = 8'h0; 1: mux_25360 = vout_peek_10485;
    endcase
  endfunction
  wire [7:0] v_25361;
  function [7:0] mux_25361(input [0:0] sel);
    case (sel) 0: mux_25361 = 8'h0; 1: mux_25361 = v_25362;
    endcase
  endfunction
  reg [7:0] v_25362 = 8'h0;
  wire [7:0] v_25363;
  wire [7:0] v_25364;
  function [7:0] mux_25364(input [0:0] sel);
    case (sel) 0: mux_25364 = 8'h0; 1: mux_25364 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25365;
  wire [7:0] v_25366;
  wire [7:0] v_25367;
  function [7:0] mux_25367(input [0:0] sel);
    case (sel) 0: mux_25367 = 8'h0; 1: mux_25367 = vout_peek_10457;
    endcase
  endfunction
  wire [7:0] v_25368;
  function [7:0] mux_25368(input [0:0] sel);
    case (sel) 0: mux_25368 = 8'h0; 1: mux_25368 = vout_peek_10448;
    endcase
  endfunction
  wire [7:0] v_25369;
  function [7:0] mux_25369(input [0:0] sel);
    case (sel) 0: mux_25369 = 8'h0; 1: mux_25369 = v_25370;
    endcase
  endfunction
  reg [7:0] v_25370 = 8'h0;
  wire [7:0] v_25371;
  wire [7:0] v_25372;
  function [7:0] mux_25372(input [0:0] sel);
    case (sel) 0: mux_25372 = 8'h0; 1: mux_25372 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25373;
  wire [7:0] v_25374;
  wire [7:0] v_25375;
  function [7:0] mux_25375(input [0:0] sel);
    case (sel) 0: mux_25375 = 8'h0; 1: mux_25375 = v_25376;
    endcase
  endfunction
  reg [7:0] v_25376 = 8'h0;
  wire [7:0] v_25377;
  wire [7:0] v_25378;
  function [7:0] mux_25378(input [0:0] sel);
    case (sel) 0: mux_25378 = 8'h0; 1: mux_25378 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25379;
  wire [7:0] v_25380;
  wire [7:0] v_25381;
  function [7:0] mux_25381(input [0:0] sel);
    case (sel) 0: mux_25381 = 8'h0; 1: mux_25381 = v_25382;
    endcase
  endfunction
  reg [7:0] v_25382 = 8'h0;
  wire [7:0] v_25383;
  wire [7:0] v_25384;
  function [7:0] mux_25384(input [0:0] sel);
    case (sel) 0: mux_25384 = 8'h0; 1: mux_25384 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25385;
  wire [7:0] v_25386;
  wire [7:0] v_25387;
  function [7:0] mux_25387(input [0:0] sel);
    case (sel) 0: mux_25387 = 8'h0; 1: mux_25387 = vout_peek_10382;
    endcase
  endfunction
  wire [7:0] v_25388;
  function [7:0] mux_25388(input [0:0] sel);
    case (sel) 0: mux_25388 = 8'h0; 1: mux_25388 = vout_peek_10373;
    endcase
  endfunction
  wire [7:0] v_25389;
  function [7:0] mux_25389(input [0:0] sel);
    case (sel) 0: mux_25389 = 8'h0; 1: mux_25389 = v_25390;
    endcase
  endfunction
  reg [7:0] v_25390 = 8'h0;
  wire [7:0] v_25391;
  wire [7:0] v_25392;
  function [7:0] mux_25392(input [0:0] sel);
    case (sel) 0: mux_25392 = 8'h0; 1: mux_25392 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25393;
  wire [7:0] v_25394;
  wire [7:0] v_25395;
  function [7:0] mux_25395(input [0:0] sel);
    case (sel) 0: mux_25395 = 8'h0; 1: mux_25395 = vout_peek_10345;
    endcase
  endfunction
  wire [7:0] v_25396;
  function [7:0] mux_25396(input [0:0] sel);
    case (sel) 0: mux_25396 = 8'h0; 1: mux_25396 = vout_peek_10336;
    endcase
  endfunction
  wire [7:0] v_25397;
  function [7:0] mux_25397(input [0:0] sel);
    case (sel) 0: mux_25397 = 8'h0; 1: mux_25397 = v_25398;
    endcase
  endfunction
  reg [7:0] v_25398 = 8'h0;
  wire [7:0] v_25399;
  wire [7:0] v_25400;
  function [7:0] mux_25400(input [0:0] sel);
    case (sel) 0: mux_25400 = 8'h0; 1: mux_25400 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25401;
  wire [7:0] v_25402;
  wire [7:0] v_25403;
  function [7:0] mux_25403(input [0:0] sel);
    case (sel) 0: mux_25403 = 8'h0; 1: mux_25403 = v_25404;
    endcase
  endfunction
  reg [7:0] v_25404 = 8'h0;
  wire [7:0] v_25405;
  wire [7:0] v_25406;
  function [7:0] mux_25406(input [0:0] sel);
    case (sel) 0: mux_25406 = 8'h0; 1: mux_25406 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25407;
  wire [7:0] v_25408;
  wire [7:0] v_25409;
  function [7:0] mux_25409(input [0:0] sel);
    case (sel) 0: mux_25409 = 8'h0; 1: mux_25409 = vout_peek_10289;
    endcase
  endfunction
  wire [7:0] v_25410;
  function [7:0] mux_25410(input [0:0] sel);
    case (sel) 0: mux_25410 = 8'h0; 1: mux_25410 = vout_peek_10280;
    endcase
  endfunction
  wire [7:0] v_25411;
  function [7:0] mux_25411(input [0:0] sel);
    case (sel) 0: mux_25411 = 8'h0; 1: mux_25411 = v_25412;
    endcase
  endfunction
  reg [7:0] v_25412 = 8'h0;
  wire [7:0] v_25413;
  wire [7:0] v_25414;
  function [7:0] mux_25414(input [0:0] sel);
    case (sel) 0: mux_25414 = 8'h0; 1: mux_25414 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25415;
  wire [7:0] v_25416;
  wire [7:0] v_25417;
  function [7:0] mux_25417(input [0:0] sel);
    case (sel) 0: mux_25417 = 8'h0; 1: mux_25417 = vout_peek_10252;
    endcase
  endfunction
  wire [7:0] v_25418;
  function [7:0] mux_25418(input [0:0] sel);
    case (sel) 0: mux_25418 = 8'h0; 1: mux_25418 = vout_peek_10243;
    endcase
  endfunction
  wire [7:0] v_25419;
  function [7:0] mux_25419(input [0:0] sel);
    case (sel) 0: mux_25419 = 8'h0; 1: mux_25419 = v_25420;
    endcase
  endfunction
  reg [7:0] v_25420 = 8'h0;
  wire [7:0] v_25421;
  wire [7:0] v_25422;
  function [7:0] mux_25422(input [0:0] sel);
    case (sel) 0: mux_25422 = 8'h0; 1: mux_25422 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25423;
  wire [7:0] v_25424;
  wire [7:0] v_25425;
  function [7:0] mux_25425(input [0:0] sel);
    case (sel) 0: mux_25425 = 8'h0; 1: mux_25425 = v_25426;
    endcase
  endfunction
  reg [7:0] v_25426 = 8'h0;
  wire [7:0] v_25427;
  wire [7:0] v_25428;
  function [7:0] mux_25428(input [0:0] sel);
    case (sel) 0: mux_25428 = 8'h0; 1: mux_25428 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25429;
  wire [7:0] v_25430;
  wire [7:0] v_25431;
  function [7:0] mux_25431(input [0:0] sel);
    case (sel) 0: mux_25431 = 8'h0; 1: mux_25431 = v_25432;
    endcase
  endfunction
  reg [7:0] v_25432 = 8'h0;
  wire [7:0] v_25433;
  wire [7:0] v_25434;
  function [7:0] mux_25434(input [0:0] sel);
    case (sel) 0: mux_25434 = 8'h0; 1: mux_25434 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25435;
  wire [7:0] v_25436;
  wire [7:0] v_25437;
  function [7:0] mux_25437(input [0:0] sel);
    case (sel) 0: mux_25437 = 8'h0; 1: mux_25437 = v_25438;
    endcase
  endfunction
  reg [7:0] v_25438 = 8'h0;
  wire [7:0] v_25439;
  wire [7:0] v_25440;
  function [7:0] mux_25440(input [0:0] sel);
    case (sel) 0: mux_25440 = 8'h0; 1: mux_25440 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25441;
  wire [7:0] v_25442;
  wire [7:0] v_25443;
  function [7:0] mux_25443(input [0:0] sel);
    case (sel) 0: mux_25443 = 8'h0; 1: mux_25443 = vout_peek_10158;
    endcase
  endfunction
  wire [7:0] v_25444;
  function [7:0] mux_25444(input [0:0] sel);
    case (sel) 0: mux_25444 = 8'h0; 1: mux_25444 = vout_peek_10149;
    endcase
  endfunction
  wire [7:0] v_25445;
  function [7:0] mux_25445(input [0:0] sel);
    case (sel) 0: mux_25445 = 8'h0; 1: mux_25445 = v_25446;
    endcase
  endfunction
  reg [7:0] v_25446 = 8'h0;
  wire [7:0] v_25447;
  wire [7:0] v_25448;
  function [7:0] mux_25448(input [0:0] sel);
    case (sel) 0: mux_25448 = 8'h0; 1: mux_25448 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25449;
  wire [7:0] v_25450;
  wire [7:0] v_25451;
  function [7:0] mux_25451(input [0:0] sel);
    case (sel) 0: mux_25451 = 8'h0; 1: mux_25451 = vout_peek_10121;
    endcase
  endfunction
  wire [7:0] v_25452;
  function [7:0] mux_25452(input [0:0] sel);
    case (sel) 0: mux_25452 = 8'h0; 1: mux_25452 = vout_peek_10112;
    endcase
  endfunction
  wire [7:0] v_25453;
  function [7:0] mux_25453(input [0:0] sel);
    case (sel) 0: mux_25453 = 8'h0; 1: mux_25453 = v_25454;
    endcase
  endfunction
  reg [7:0] v_25454 = 8'h0;
  wire [7:0] v_25455;
  wire [7:0] v_25456;
  function [7:0] mux_25456(input [0:0] sel);
    case (sel) 0: mux_25456 = 8'h0; 1: mux_25456 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25457;
  wire [7:0] v_25458;
  wire [7:0] v_25459;
  function [7:0] mux_25459(input [0:0] sel);
    case (sel) 0: mux_25459 = 8'h0; 1: mux_25459 = v_25460;
    endcase
  endfunction
  reg [7:0] v_25460 = 8'h0;
  wire [7:0] v_25461;
  wire [7:0] v_25462;
  function [7:0] mux_25462(input [0:0] sel);
    case (sel) 0: mux_25462 = 8'h0; 1: mux_25462 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25463;
  wire [7:0] v_25464;
  wire [7:0] v_25465;
  function [7:0] mux_25465(input [0:0] sel);
    case (sel) 0: mux_25465 = 8'h0; 1: mux_25465 = vout_peek_10065;
    endcase
  endfunction
  wire [7:0] v_25466;
  function [7:0] mux_25466(input [0:0] sel);
    case (sel) 0: mux_25466 = 8'h0; 1: mux_25466 = vout_peek_10056;
    endcase
  endfunction
  wire [7:0] v_25467;
  function [7:0] mux_25467(input [0:0] sel);
    case (sel) 0: mux_25467 = 8'h0; 1: mux_25467 = v_25468;
    endcase
  endfunction
  reg [7:0] v_25468 = 8'h0;
  wire [7:0] v_25469;
  wire [7:0] v_25470;
  function [7:0] mux_25470(input [0:0] sel);
    case (sel) 0: mux_25470 = 8'h0; 1: mux_25470 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25471;
  wire [7:0] v_25472;
  wire [7:0] v_25473;
  function [7:0] mux_25473(input [0:0] sel);
    case (sel) 0: mux_25473 = 8'h0; 1: mux_25473 = vout_peek_10028;
    endcase
  endfunction
  wire [7:0] v_25474;
  function [7:0] mux_25474(input [0:0] sel);
    case (sel) 0: mux_25474 = 8'h0; 1: mux_25474 = vout_peek_10019;
    endcase
  endfunction
  wire [7:0] v_25475;
  function [7:0] mux_25475(input [0:0] sel);
    case (sel) 0: mux_25475 = 8'h0; 1: mux_25475 = v_25476;
    endcase
  endfunction
  reg [7:0] v_25476 = 8'h0;
  wire [7:0] v_25477;
  wire [7:0] v_25478;
  function [7:0] mux_25478(input [0:0] sel);
    case (sel) 0: mux_25478 = 8'h0; 1: mux_25478 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25479;
  wire [7:0] v_25480;
  wire [7:0] v_25481;
  function [7:0] mux_25481(input [0:0] sel);
    case (sel) 0: mux_25481 = 8'h0; 1: mux_25481 = v_25482;
    endcase
  endfunction
  reg [7:0] v_25482 = 8'h0;
  wire [7:0] v_25483;
  wire [7:0] v_25484;
  function [7:0] mux_25484(input [0:0] sel);
    case (sel) 0: mux_25484 = 8'h0; 1: mux_25484 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25485;
  wire [7:0] v_25486;
  wire [7:0] v_25487;
  function [7:0] mux_25487(input [0:0] sel);
    case (sel) 0: mux_25487 = 8'h0; 1: mux_25487 = v_25488;
    endcase
  endfunction
  reg [7:0] v_25488 = 8'h0;
  wire [7:0] v_25489;
  wire [7:0] v_25490;
  function [7:0] mux_25490(input [0:0] sel);
    case (sel) 0: mux_25490 = 8'h0; 1: mux_25490 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25491;
  wire [7:0] v_25492;
  wire [7:0] v_25493;
  function [7:0] mux_25493(input [0:0] sel);
    case (sel) 0: mux_25493 = 8'h0; 1: mux_25493 = vout_peek_9953;
    endcase
  endfunction
  wire [7:0] v_25494;
  function [7:0] mux_25494(input [0:0] sel);
    case (sel) 0: mux_25494 = 8'h0; 1: mux_25494 = vout_peek_9944;
    endcase
  endfunction
  wire [7:0] v_25495;
  function [7:0] mux_25495(input [0:0] sel);
    case (sel) 0: mux_25495 = 8'h0; 1: mux_25495 = v_25496;
    endcase
  endfunction
  reg [7:0] v_25496 = 8'h0;
  wire [7:0] v_25497;
  wire [7:0] v_25498;
  function [7:0] mux_25498(input [0:0] sel);
    case (sel) 0: mux_25498 = 8'h0; 1: mux_25498 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25499;
  wire [7:0] v_25500;
  wire [7:0] v_25501;
  function [7:0] mux_25501(input [0:0] sel);
    case (sel) 0: mux_25501 = 8'h0; 1: mux_25501 = vout_peek_9916;
    endcase
  endfunction
  wire [7:0] v_25502;
  function [7:0] mux_25502(input [0:0] sel);
    case (sel) 0: mux_25502 = 8'h0; 1: mux_25502 = vout_peek_9907;
    endcase
  endfunction
  wire [7:0] v_25503;
  function [7:0] mux_25503(input [0:0] sel);
    case (sel) 0: mux_25503 = 8'h0; 1: mux_25503 = v_25504;
    endcase
  endfunction
  reg [7:0] v_25504 = 8'h0;
  wire [7:0] v_25505;
  wire [7:0] v_25506;
  function [7:0] mux_25506(input [0:0] sel);
    case (sel) 0: mux_25506 = 8'h0; 1: mux_25506 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25507;
  wire [7:0] v_25508;
  wire [7:0] v_25509;
  function [7:0] mux_25509(input [0:0] sel);
    case (sel) 0: mux_25509 = 8'h0; 1: mux_25509 = v_25510;
    endcase
  endfunction
  reg [7:0] v_25510 = 8'h0;
  wire [7:0] v_25511;
  wire [7:0] v_25512;
  function [7:0] mux_25512(input [0:0] sel);
    case (sel) 0: mux_25512 = 8'h0; 1: mux_25512 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25513;
  wire [7:0] v_25514;
  wire [7:0] v_25515;
  function [7:0] mux_25515(input [0:0] sel);
    case (sel) 0: mux_25515 = 8'h0; 1: mux_25515 = vout_peek_9860;
    endcase
  endfunction
  wire [7:0] v_25516;
  function [7:0] mux_25516(input [0:0] sel);
    case (sel) 0: mux_25516 = 8'h0; 1: mux_25516 = vout_peek_9851;
    endcase
  endfunction
  wire [7:0] v_25517;
  function [7:0] mux_25517(input [0:0] sel);
    case (sel) 0: mux_25517 = 8'h0; 1: mux_25517 = v_25518;
    endcase
  endfunction
  reg [7:0] v_25518 = 8'h0;
  wire [7:0] v_25519;
  wire [7:0] v_25520;
  function [7:0] mux_25520(input [0:0] sel);
    case (sel) 0: mux_25520 = 8'h0; 1: mux_25520 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25521;
  wire [7:0] v_25522;
  wire [7:0] v_25523;
  function [7:0] mux_25523(input [0:0] sel);
    case (sel) 0: mux_25523 = 8'h0; 1: mux_25523 = vout_peek_9823;
    endcase
  endfunction
  wire [7:0] v_25524;
  function [7:0] mux_25524(input [0:0] sel);
    case (sel) 0: mux_25524 = 8'h0; 1: mux_25524 = vout_peek_9814;
    endcase
  endfunction
  wire [7:0] v_25525;
  function [7:0] mux_25525(input [0:0] sel);
    case (sel) 0: mux_25525 = 8'h0; 1: mux_25525 = v_25526;
    endcase
  endfunction
  reg [7:0] v_25526 = 8'h0;
  wire [7:0] v_25527;
  wire [7:0] v_25528;
  function [7:0] mux_25528(input [0:0] sel);
    case (sel) 0: mux_25528 = 8'h0; 1: mux_25528 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25529;
  wire [7:0] v_25530;
  wire [7:0] v_25531;
  function [7:0] mux_25531(input [0:0] sel);
    case (sel) 0: mux_25531 = 8'h0; 1: mux_25531 = v_25532;
    endcase
  endfunction
  reg [7:0] v_25532 = 8'h0;
  wire [7:0] v_25533;
  wire [7:0] v_25534;
  function [7:0] mux_25534(input [0:0] sel);
    case (sel) 0: mux_25534 = 8'h0; 1: mux_25534 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25535;
  wire [7:0] v_25536;
  wire [7:0] v_25537;
  function [7:0] mux_25537(input [0:0] sel);
    case (sel) 0: mux_25537 = 8'h0; 1: mux_25537 = v_25538;
    endcase
  endfunction
  reg [7:0] v_25538 = 8'h0;
  wire [7:0] v_25539;
  wire [7:0] v_25540;
  function [7:0] mux_25540(input [0:0] sel);
    case (sel) 0: mux_25540 = 8'h0; 1: mux_25540 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25541;
  wire [7:0] v_25542;
  wire [7:0] v_25543;
  function [7:0] mux_25543(input [0:0] sel);
    case (sel) 0: mux_25543 = 8'h0; 1: mux_25543 = v_25544;
    endcase
  endfunction
  reg [7:0] v_25544 = 8'h0;
  wire [7:0] v_25545;
  wire [7:0] v_25546;
  function [7:0] mux_25546(input [0:0] sel);
    case (sel) 0: mux_25546 = 8'h0; 1: mux_25546 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25547;
  wire [7:0] v_25548;
  wire [7:0] v_25549;
  function [7:0] mux_25549(input [0:0] sel);
    case (sel) 0: mux_25549 = 8'h0; 1: mux_25549 = v_25550;
    endcase
  endfunction
  reg [7:0] v_25550 = 8'h0;
  wire [7:0] v_25551;
  wire [7:0] v_25552;
  function [7:0] mux_25552(input [0:0] sel);
    case (sel) 0: mux_25552 = 8'h0; 1: mux_25552 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25553;
  wire [7:0] v_25554;
  wire [7:0] v_25555;
  function [7:0] mux_25555(input [0:0] sel);
    case (sel) 0: mux_25555 = 8'h0; 1: mux_25555 = v_25556;
    endcase
  endfunction
  reg [7:0] v_25556 = 8'h0;
  wire [7:0] v_25557;
  wire [7:0] v_25558;
  function [7:0] mux_25558(input [0:0] sel);
    case (sel) 0: mux_25558 = 8'h0; 1: mux_25558 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25559;
  wire [7:0] v_25560;
  wire [7:0] v_25561;
  function [7:0] mux_25561(input [0:0] sel);
    case (sel) 0: mux_25561 = 8'h0; 1: mux_25561 = vout_peek_9691;
    endcase
  endfunction
  wire [7:0] v_25562;
  function [7:0] mux_25562(input [0:0] sel);
    case (sel) 0: mux_25562 = 8'h0; 1: mux_25562 = vout_peek_9682;
    endcase
  endfunction
  wire [7:0] v_25563;
  function [7:0] mux_25563(input [0:0] sel);
    case (sel) 0: mux_25563 = 8'h0; 1: mux_25563 = v_25564;
    endcase
  endfunction
  reg [7:0] v_25564 = 8'h0;
  wire [7:0] v_25565;
  wire [7:0] v_25566;
  function [7:0] mux_25566(input [0:0] sel);
    case (sel) 0: mux_25566 = 8'h0; 1: mux_25566 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25567;
  wire [7:0] v_25568;
  wire [7:0] v_25569;
  function [7:0] mux_25569(input [0:0] sel);
    case (sel) 0: mux_25569 = 8'h0; 1: mux_25569 = vout_peek_9654;
    endcase
  endfunction
  wire [7:0] v_25570;
  function [7:0] mux_25570(input [0:0] sel);
    case (sel) 0: mux_25570 = 8'h0; 1: mux_25570 = vout_peek_9645;
    endcase
  endfunction
  wire [7:0] v_25571;
  function [7:0] mux_25571(input [0:0] sel);
    case (sel) 0: mux_25571 = 8'h0; 1: mux_25571 = v_25572;
    endcase
  endfunction
  reg [7:0] v_25572 = 8'h0;
  wire [7:0] v_25573;
  wire [7:0] v_25574;
  function [7:0] mux_25574(input [0:0] sel);
    case (sel) 0: mux_25574 = 8'h0; 1: mux_25574 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25575;
  wire [7:0] v_25576;
  wire [7:0] v_25577;
  function [7:0] mux_25577(input [0:0] sel);
    case (sel) 0: mux_25577 = 8'h0; 1: mux_25577 = v_25578;
    endcase
  endfunction
  reg [7:0] v_25578 = 8'h0;
  wire [7:0] v_25579;
  wire [7:0] v_25580;
  function [7:0] mux_25580(input [0:0] sel);
    case (sel) 0: mux_25580 = 8'h0; 1: mux_25580 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25581;
  wire [7:0] v_25582;
  wire [7:0] v_25583;
  function [7:0] mux_25583(input [0:0] sel);
    case (sel) 0: mux_25583 = 8'h0; 1: mux_25583 = vout_peek_9598;
    endcase
  endfunction
  wire [7:0] v_25584;
  function [7:0] mux_25584(input [0:0] sel);
    case (sel) 0: mux_25584 = 8'h0; 1: mux_25584 = vout_peek_9589;
    endcase
  endfunction
  wire [7:0] v_25585;
  function [7:0] mux_25585(input [0:0] sel);
    case (sel) 0: mux_25585 = 8'h0; 1: mux_25585 = v_25586;
    endcase
  endfunction
  reg [7:0] v_25586 = 8'h0;
  wire [7:0] v_25587;
  wire [7:0] v_25588;
  function [7:0] mux_25588(input [0:0] sel);
    case (sel) 0: mux_25588 = 8'h0; 1: mux_25588 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25589;
  wire [7:0] v_25590;
  wire [7:0] v_25591;
  function [7:0] mux_25591(input [0:0] sel);
    case (sel) 0: mux_25591 = 8'h0; 1: mux_25591 = vout_peek_9561;
    endcase
  endfunction
  wire [7:0] v_25592;
  function [7:0] mux_25592(input [0:0] sel);
    case (sel) 0: mux_25592 = 8'h0; 1: mux_25592 = vout_peek_9552;
    endcase
  endfunction
  wire [7:0] v_25593;
  function [7:0] mux_25593(input [0:0] sel);
    case (sel) 0: mux_25593 = 8'h0; 1: mux_25593 = v_25594;
    endcase
  endfunction
  reg [7:0] v_25594 = 8'h0;
  wire [7:0] v_25595;
  wire [7:0] v_25596;
  function [7:0] mux_25596(input [0:0] sel);
    case (sel) 0: mux_25596 = 8'h0; 1: mux_25596 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25597;
  wire [7:0] v_25598;
  wire [7:0] v_25599;
  function [7:0] mux_25599(input [0:0] sel);
    case (sel) 0: mux_25599 = 8'h0; 1: mux_25599 = v_25600;
    endcase
  endfunction
  reg [7:0] v_25600 = 8'h0;
  wire [7:0] v_25601;
  wire [7:0] v_25602;
  function [7:0] mux_25602(input [0:0] sel);
    case (sel) 0: mux_25602 = 8'h0; 1: mux_25602 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25603;
  wire [7:0] v_25604;
  wire [7:0] v_25605;
  function [7:0] mux_25605(input [0:0] sel);
    case (sel) 0: mux_25605 = 8'h0; 1: mux_25605 = v_25606;
    endcase
  endfunction
  reg [7:0] v_25606 = 8'h0;
  wire [7:0] v_25607;
  wire [7:0] v_25608;
  function [7:0] mux_25608(input [0:0] sel);
    case (sel) 0: mux_25608 = 8'h0; 1: mux_25608 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25609;
  wire [7:0] v_25610;
  wire [7:0] v_25611;
  function [7:0] mux_25611(input [0:0] sel);
    case (sel) 0: mux_25611 = 8'h0; 1: mux_25611 = vout_peek_9486;
    endcase
  endfunction
  wire [7:0] v_25612;
  function [7:0] mux_25612(input [0:0] sel);
    case (sel) 0: mux_25612 = 8'h0; 1: mux_25612 = vout_peek_9477;
    endcase
  endfunction
  wire [7:0] v_25613;
  function [7:0] mux_25613(input [0:0] sel);
    case (sel) 0: mux_25613 = 8'h0; 1: mux_25613 = v_25614;
    endcase
  endfunction
  reg [7:0] v_25614 = 8'h0;
  wire [7:0] v_25615;
  wire [7:0] v_25616;
  function [7:0] mux_25616(input [0:0] sel);
    case (sel) 0: mux_25616 = 8'h0; 1: mux_25616 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25617;
  wire [7:0] v_25618;
  wire [7:0] v_25619;
  function [7:0] mux_25619(input [0:0] sel);
    case (sel) 0: mux_25619 = 8'h0; 1: mux_25619 = vout_peek_9449;
    endcase
  endfunction
  wire [7:0] v_25620;
  function [7:0] mux_25620(input [0:0] sel);
    case (sel) 0: mux_25620 = 8'h0; 1: mux_25620 = vout_peek_9440;
    endcase
  endfunction
  wire [7:0] v_25621;
  function [7:0] mux_25621(input [0:0] sel);
    case (sel) 0: mux_25621 = 8'h0; 1: mux_25621 = v_25622;
    endcase
  endfunction
  reg [7:0] v_25622 = 8'h0;
  wire [7:0] v_25623;
  wire [7:0] v_25624;
  function [7:0] mux_25624(input [0:0] sel);
    case (sel) 0: mux_25624 = 8'h0; 1: mux_25624 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25625;
  wire [7:0] v_25626;
  wire [7:0] v_25627;
  function [7:0] mux_25627(input [0:0] sel);
    case (sel) 0: mux_25627 = 8'h0; 1: mux_25627 = v_25628;
    endcase
  endfunction
  reg [7:0] v_25628 = 8'h0;
  wire [7:0] v_25629;
  wire [7:0] v_25630;
  function [7:0] mux_25630(input [0:0] sel);
    case (sel) 0: mux_25630 = 8'h0; 1: mux_25630 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25631;
  wire [7:0] v_25632;
  wire [7:0] v_25633;
  function [7:0] mux_25633(input [0:0] sel);
    case (sel) 0: mux_25633 = 8'h0; 1: mux_25633 = vout_peek_9393;
    endcase
  endfunction
  wire [7:0] v_25634;
  function [7:0] mux_25634(input [0:0] sel);
    case (sel) 0: mux_25634 = 8'h0; 1: mux_25634 = vout_peek_9384;
    endcase
  endfunction
  wire [7:0] v_25635;
  function [7:0] mux_25635(input [0:0] sel);
    case (sel) 0: mux_25635 = 8'h0; 1: mux_25635 = v_25636;
    endcase
  endfunction
  reg [7:0] v_25636 = 8'h0;
  wire [7:0] v_25637;
  wire [7:0] v_25638;
  function [7:0] mux_25638(input [0:0] sel);
    case (sel) 0: mux_25638 = 8'h0; 1: mux_25638 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25639;
  wire [7:0] v_25640;
  wire [7:0] v_25641;
  function [7:0] mux_25641(input [0:0] sel);
    case (sel) 0: mux_25641 = 8'h0; 1: mux_25641 = vout_peek_9356;
    endcase
  endfunction
  wire [7:0] v_25642;
  function [7:0] mux_25642(input [0:0] sel);
    case (sel) 0: mux_25642 = 8'h0; 1: mux_25642 = vout_peek_9347;
    endcase
  endfunction
  wire [7:0] v_25643;
  function [7:0] mux_25643(input [0:0] sel);
    case (sel) 0: mux_25643 = 8'h0; 1: mux_25643 = v_25644;
    endcase
  endfunction
  reg [7:0] v_25644 = 8'h0;
  wire [7:0] v_25645;
  wire [7:0] v_25646;
  function [7:0] mux_25646(input [0:0] sel);
    case (sel) 0: mux_25646 = 8'h0; 1: mux_25646 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25647;
  wire [7:0] v_25648;
  wire [7:0] v_25649;
  function [7:0] mux_25649(input [0:0] sel);
    case (sel) 0: mux_25649 = 8'h0; 1: mux_25649 = v_25650;
    endcase
  endfunction
  reg [7:0] v_25650 = 8'h0;
  wire [7:0] v_25651;
  wire [7:0] v_25652;
  function [7:0] mux_25652(input [0:0] sel);
    case (sel) 0: mux_25652 = 8'h0; 1: mux_25652 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25653;
  wire [7:0] v_25654;
  wire [7:0] v_25655;
  function [7:0] mux_25655(input [0:0] sel);
    case (sel) 0: mux_25655 = 8'h0; 1: mux_25655 = v_25656;
    endcase
  endfunction
  reg [7:0] v_25656 = 8'h0;
  wire [7:0] v_25657;
  wire [7:0] v_25658;
  function [7:0] mux_25658(input [0:0] sel);
    case (sel) 0: mux_25658 = 8'h0; 1: mux_25658 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25659;
  wire [7:0] v_25660;
  wire [7:0] v_25661;
  function [7:0] mux_25661(input [0:0] sel);
    case (sel) 0: mux_25661 = 8'h0; 1: mux_25661 = v_25662;
    endcase
  endfunction
  reg [7:0] v_25662 = 8'h0;
  wire [7:0] v_25663;
  wire [7:0] v_25664;
  function [7:0] mux_25664(input [0:0] sel);
    case (sel) 0: mux_25664 = 8'h0; 1: mux_25664 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25665;
  wire [7:0] v_25666;
  wire [7:0] v_25667;
  function [7:0] mux_25667(input [0:0] sel);
    case (sel) 0: mux_25667 = 8'h0; 1: mux_25667 = vout_peek_9262;
    endcase
  endfunction
  wire [7:0] v_25668;
  function [7:0] mux_25668(input [0:0] sel);
    case (sel) 0: mux_25668 = 8'h0; 1: mux_25668 = vout_peek_9253;
    endcase
  endfunction
  wire [7:0] v_25669;
  function [7:0] mux_25669(input [0:0] sel);
    case (sel) 0: mux_25669 = 8'h0; 1: mux_25669 = v_25670;
    endcase
  endfunction
  reg [7:0] v_25670 = 8'h0;
  wire [7:0] v_25671;
  wire [7:0] v_25672;
  function [7:0] mux_25672(input [0:0] sel);
    case (sel) 0: mux_25672 = 8'h0; 1: mux_25672 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25673;
  wire [7:0] v_25674;
  wire [7:0] v_25675;
  function [7:0] mux_25675(input [0:0] sel);
    case (sel) 0: mux_25675 = 8'h0; 1: mux_25675 = vout_peek_9225;
    endcase
  endfunction
  wire [7:0] v_25676;
  function [7:0] mux_25676(input [0:0] sel);
    case (sel) 0: mux_25676 = 8'h0; 1: mux_25676 = vout_peek_9216;
    endcase
  endfunction
  wire [7:0] v_25677;
  function [7:0] mux_25677(input [0:0] sel);
    case (sel) 0: mux_25677 = 8'h0; 1: mux_25677 = v_25678;
    endcase
  endfunction
  reg [7:0] v_25678 = 8'h0;
  wire [7:0] v_25679;
  wire [7:0] v_25680;
  function [7:0] mux_25680(input [0:0] sel);
    case (sel) 0: mux_25680 = 8'h0; 1: mux_25680 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25681;
  wire [7:0] v_25682;
  wire [7:0] v_25683;
  function [7:0] mux_25683(input [0:0] sel);
    case (sel) 0: mux_25683 = 8'h0; 1: mux_25683 = v_25684;
    endcase
  endfunction
  reg [7:0] v_25684 = 8'h0;
  wire [7:0] v_25685;
  wire [7:0] v_25686;
  function [7:0] mux_25686(input [0:0] sel);
    case (sel) 0: mux_25686 = 8'h0; 1: mux_25686 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25687;
  wire [7:0] v_25688;
  wire [7:0] v_25689;
  function [7:0] mux_25689(input [0:0] sel);
    case (sel) 0: mux_25689 = 8'h0; 1: mux_25689 = vout_peek_9169;
    endcase
  endfunction
  wire [7:0] v_25690;
  function [7:0] mux_25690(input [0:0] sel);
    case (sel) 0: mux_25690 = 8'h0; 1: mux_25690 = vout_peek_9160;
    endcase
  endfunction
  wire [7:0] v_25691;
  function [7:0] mux_25691(input [0:0] sel);
    case (sel) 0: mux_25691 = 8'h0; 1: mux_25691 = v_25692;
    endcase
  endfunction
  reg [7:0] v_25692 = 8'h0;
  wire [7:0] v_25693;
  wire [7:0] v_25694;
  function [7:0] mux_25694(input [0:0] sel);
    case (sel) 0: mux_25694 = 8'h0; 1: mux_25694 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25695;
  wire [7:0] v_25696;
  wire [7:0] v_25697;
  function [7:0] mux_25697(input [0:0] sel);
    case (sel) 0: mux_25697 = 8'h0; 1: mux_25697 = vout_peek_9132;
    endcase
  endfunction
  wire [7:0] v_25698;
  function [7:0] mux_25698(input [0:0] sel);
    case (sel) 0: mux_25698 = 8'h0; 1: mux_25698 = vout_peek_9123;
    endcase
  endfunction
  wire [7:0] v_25699;
  function [7:0] mux_25699(input [0:0] sel);
    case (sel) 0: mux_25699 = 8'h0; 1: mux_25699 = v_25700;
    endcase
  endfunction
  reg [7:0] v_25700 = 8'h0;
  wire [7:0] v_25701;
  wire [7:0] v_25702;
  function [7:0] mux_25702(input [0:0] sel);
    case (sel) 0: mux_25702 = 8'h0; 1: mux_25702 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25703;
  wire [7:0] v_25704;
  wire [7:0] v_25705;
  function [7:0] mux_25705(input [0:0] sel);
    case (sel) 0: mux_25705 = 8'h0; 1: mux_25705 = v_25706;
    endcase
  endfunction
  reg [7:0] v_25706 = 8'h0;
  wire [7:0] v_25707;
  wire [7:0] v_25708;
  function [7:0] mux_25708(input [0:0] sel);
    case (sel) 0: mux_25708 = 8'h0; 1: mux_25708 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25709;
  wire [7:0] v_25710;
  wire [7:0] v_25711;
  function [7:0] mux_25711(input [0:0] sel);
    case (sel) 0: mux_25711 = 8'h0; 1: mux_25711 = v_25712;
    endcase
  endfunction
  reg [7:0] v_25712 = 8'h0;
  wire [7:0] v_25713;
  wire [7:0] v_25714;
  function [7:0] mux_25714(input [0:0] sel);
    case (sel) 0: mux_25714 = 8'h0; 1: mux_25714 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25715;
  wire [7:0] v_25716;
  wire [7:0] v_25717;
  function [7:0] mux_25717(input [0:0] sel);
    case (sel) 0: mux_25717 = 8'h0; 1: mux_25717 = vout_peek_9057;
    endcase
  endfunction
  wire [7:0] v_25718;
  function [7:0] mux_25718(input [0:0] sel);
    case (sel) 0: mux_25718 = 8'h0; 1: mux_25718 = vout_peek_9048;
    endcase
  endfunction
  wire [7:0] v_25719;
  function [7:0] mux_25719(input [0:0] sel);
    case (sel) 0: mux_25719 = 8'h0; 1: mux_25719 = v_25720;
    endcase
  endfunction
  reg [7:0] v_25720 = 8'h0;
  wire [7:0] v_25721;
  wire [7:0] v_25722;
  function [7:0] mux_25722(input [0:0] sel);
    case (sel) 0: mux_25722 = 8'h0; 1: mux_25722 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25723;
  wire [7:0] v_25724;
  wire [7:0] v_25725;
  function [7:0] mux_25725(input [0:0] sel);
    case (sel) 0: mux_25725 = 8'h0; 1: mux_25725 = vout_peek_9020;
    endcase
  endfunction
  wire [7:0] v_25726;
  function [7:0] mux_25726(input [0:0] sel);
    case (sel) 0: mux_25726 = 8'h0; 1: mux_25726 = vout_peek_9011;
    endcase
  endfunction
  wire [7:0] v_25727;
  function [7:0] mux_25727(input [0:0] sel);
    case (sel) 0: mux_25727 = 8'h0; 1: mux_25727 = v_25728;
    endcase
  endfunction
  reg [7:0] v_25728 = 8'h0;
  wire [7:0] v_25729;
  wire [7:0] v_25730;
  function [7:0] mux_25730(input [0:0] sel);
    case (sel) 0: mux_25730 = 8'h0; 1: mux_25730 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25731;
  wire [7:0] v_25732;
  wire [7:0] v_25733;
  function [7:0] mux_25733(input [0:0] sel);
    case (sel) 0: mux_25733 = 8'h0; 1: mux_25733 = v_25734;
    endcase
  endfunction
  reg [7:0] v_25734 = 8'h0;
  wire [7:0] v_25735;
  wire [7:0] v_25736;
  function [7:0] mux_25736(input [0:0] sel);
    case (sel) 0: mux_25736 = 8'h0; 1: mux_25736 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25737;
  wire [7:0] v_25738;
  wire [7:0] v_25739;
  function [7:0] mux_25739(input [0:0] sel);
    case (sel) 0: mux_25739 = 8'h0; 1: mux_25739 = vout_peek_8964;
    endcase
  endfunction
  wire [7:0] v_25740;
  function [7:0] mux_25740(input [0:0] sel);
    case (sel) 0: mux_25740 = 8'h0; 1: mux_25740 = vout_peek_8955;
    endcase
  endfunction
  wire [7:0] v_25741;
  function [7:0] mux_25741(input [0:0] sel);
    case (sel) 0: mux_25741 = 8'h0; 1: mux_25741 = v_25742;
    endcase
  endfunction
  reg [7:0] v_25742 = 8'h0;
  wire [7:0] v_25743;
  wire [7:0] v_25744;
  function [7:0] mux_25744(input [0:0] sel);
    case (sel) 0: mux_25744 = 8'h0; 1: mux_25744 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25745;
  wire [7:0] v_25746;
  wire [7:0] v_25747;
  function [7:0] mux_25747(input [0:0] sel);
    case (sel) 0: mux_25747 = 8'h0; 1: mux_25747 = vout_peek_8927;
    endcase
  endfunction
  wire [7:0] v_25748;
  function [7:0] mux_25748(input [0:0] sel);
    case (sel) 0: mux_25748 = 8'h0; 1: mux_25748 = vout_peek_8918;
    endcase
  endfunction
  wire [7:0] v_25749;
  function [7:0] mux_25749(input [0:0] sel);
    case (sel) 0: mux_25749 = 8'h0; 1: mux_25749 = v_25750;
    endcase
  endfunction
  reg [7:0] v_25750 = 8'h0;
  wire [7:0] v_25751;
  wire [7:0] v_25752;
  function [7:0] mux_25752(input [0:0] sel);
    case (sel) 0: mux_25752 = 8'h0; 1: mux_25752 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25753;
  wire [7:0] v_25754;
  wire [7:0] v_25755;
  function [7:0] mux_25755(input [0:0] sel);
    case (sel) 0: mux_25755 = 8'h0; 1: mux_25755 = v_25756;
    endcase
  endfunction
  reg [7:0] v_25756 = 8'h0;
  wire [7:0] v_25757;
  wire [7:0] v_25758;
  function [7:0] mux_25758(input [0:0] sel);
    case (sel) 0: mux_25758 = 8'h0; 1: mux_25758 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25759;
  wire [7:0] v_25760;
  wire [7:0] v_25761;
  function [7:0] mux_25761(input [0:0] sel);
    case (sel) 0: mux_25761 = 8'h0; 1: mux_25761 = v_25762;
    endcase
  endfunction
  reg [7:0] v_25762 = 8'h0;
  wire [7:0] v_25763;
  wire [7:0] v_25764;
  function [7:0] mux_25764(input [0:0] sel);
    case (sel) 0: mux_25764 = 8'h0; 1: mux_25764 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25765;
  wire [7:0] v_25766;
  wire [7:0] v_25767;
  function [7:0] mux_25767(input [0:0] sel);
    case (sel) 0: mux_25767 = 8'h0; 1: mux_25767 = v_25768;
    endcase
  endfunction
  reg [7:0] v_25768 = 8'h0;
  wire [7:0] v_25769;
  wire [7:0] v_25770;
  function [7:0] mux_25770(input [0:0] sel);
    case (sel) 0: mux_25770 = 8'h0; 1: mux_25770 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25771;
  wire [7:0] v_25772;
  wire [7:0] v_25773;
  function [7:0] mux_25773(input [0:0] sel);
    case (sel) 0: mux_25773 = 8'h0; 1: mux_25773 = v_25774;
    endcase
  endfunction
  reg [7:0] v_25774 = 8'h0;
  wire [7:0] v_25775;
  wire [7:0] v_25776;
  function [7:0] mux_25776(input [0:0] sel);
    case (sel) 0: mux_25776 = 8'h0; 1: mux_25776 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25777;
  wire [7:0] v_25778;
  wire [7:0] v_25779;
  function [7:0] mux_25779(input [0:0] sel);
    case (sel) 0: mux_25779 = 8'h0; 1: mux_25779 = vout_peek_8814;
    endcase
  endfunction
  wire [7:0] v_25780;
  function [7:0] mux_25780(input [0:0] sel);
    case (sel) 0: mux_25780 = 8'h0; 1: mux_25780 = vout_peek_8805;
    endcase
  endfunction
  wire [7:0] v_25781;
  function [7:0] mux_25781(input [0:0] sel);
    case (sel) 0: mux_25781 = 8'h0; 1: mux_25781 = v_25782;
    endcase
  endfunction
  reg [7:0] v_25782 = 8'h0;
  wire [7:0] v_25783;
  wire [7:0] v_25784;
  function [7:0] mux_25784(input [0:0] sel);
    case (sel) 0: mux_25784 = 8'h0; 1: mux_25784 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25785;
  wire [7:0] v_25786;
  wire [7:0] v_25787;
  function [7:0] mux_25787(input [0:0] sel);
    case (sel) 0: mux_25787 = 8'h0; 1: mux_25787 = vout_peek_8777;
    endcase
  endfunction
  wire [7:0] v_25788;
  function [7:0] mux_25788(input [0:0] sel);
    case (sel) 0: mux_25788 = 8'h0; 1: mux_25788 = vout_peek_8768;
    endcase
  endfunction
  wire [7:0] v_25789;
  function [7:0] mux_25789(input [0:0] sel);
    case (sel) 0: mux_25789 = 8'h0; 1: mux_25789 = v_25790;
    endcase
  endfunction
  reg [7:0] v_25790 = 8'h0;
  wire [7:0] v_25791;
  wire [7:0] v_25792;
  function [7:0] mux_25792(input [0:0] sel);
    case (sel) 0: mux_25792 = 8'h0; 1: mux_25792 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25793;
  wire [7:0] v_25794;
  wire [7:0] v_25795;
  function [7:0] mux_25795(input [0:0] sel);
    case (sel) 0: mux_25795 = 8'h0; 1: mux_25795 = v_25796;
    endcase
  endfunction
  reg [7:0] v_25796 = 8'h0;
  wire [7:0] v_25797;
  wire [7:0] v_25798;
  function [7:0] mux_25798(input [0:0] sel);
    case (sel) 0: mux_25798 = 8'h0; 1: mux_25798 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25799;
  wire [7:0] v_25800;
  wire [7:0] v_25801;
  function [7:0] mux_25801(input [0:0] sel);
    case (sel) 0: mux_25801 = 8'h0; 1: mux_25801 = vout_peek_8721;
    endcase
  endfunction
  wire [7:0] v_25802;
  function [7:0] mux_25802(input [0:0] sel);
    case (sel) 0: mux_25802 = 8'h0; 1: mux_25802 = vout_peek_8712;
    endcase
  endfunction
  wire [7:0] v_25803;
  function [7:0] mux_25803(input [0:0] sel);
    case (sel) 0: mux_25803 = 8'h0; 1: mux_25803 = v_25804;
    endcase
  endfunction
  reg [7:0] v_25804 = 8'h0;
  wire [7:0] v_25805;
  wire [7:0] v_25806;
  function [7:0] mux_25806(input [0:0] sel);
    case (sel) 0: mux_25806 = 8'h0; 1: mux_25806 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25807;
  wire [7:0] v_25808;
  wire [7:0] v_25809;
  function [7:0] mux_25809(input [0:0] sel);
    case (sel) 0: mux_25809 = 8'h0; 1: mux_25809 = vout_peek_8684;
    endcase
  endfunction
  wire [7:0] v_25810;
  function [7:0] mux_25810(input [0:0] sel);
    case (sel) 0: mux_25810 = 8'h0; 1: mux_25810 = vout_peek_8675;
    endcase
  endfunction
  wire [7:0] v_25811;
  function [7:0] mux_25811(input [0:0] sel);
    case (sel) 0: mux_25811 = 8'h0; 1: mux_25811 = v_25812;
    endcase
  endfunction
  reg [7:0] v_25812 = 8'h0;
  wire [7:0] v_25813;
  wire [7:0] v_25814;
  function [7:0] mux_25814(input [0:0] sel);
    case (sel) 0: mux_25814 = 8'h0; 1: mux_25814 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25815;
  wire [7:0] v_25816;
  wire [7:0] v_25817;
  function [7:0] mux_25817(input [0:0] sel);
    case (sel) 0: mux_25817 = 8'h0; 1: mux_25817 = v_25818;
    endcase
  endfunction
  reg [7:0] v_25818 = 8'h0;
  wire [7:0] v_25819;
  wire [7:0] v_25820;
  function [7:0] mux_25820(input [0:0] sel);
    case (sel) 0: mux_25820 = 8'h0; 1: mux_25820 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25821;
  wire [7:0] v_25822;
  wire [7:0] v_25823;
  function [7:0] mux_25823(input [0:0] sel);
    case (sel) 0: mux_25823 = 8'h0; 1: mux_25823 = v_25824;
    endcase
  endfunction
  reg [7:0] v_25824 = 8'h0;
  wire [7:0] v_25825;
  wire [7:0] v_25826;
  function [7:0] mux_25826(input [0:0] sel);
    case (sel) 0: mux_25826 = 8'h0; 1: mux_25826 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25827;
  wire [7:0] v_25828;
  wire [7:0] v_25829;
  function [7:0] mux_25829(input [0:0] sel);
    case (sel) 0: mux_25829 = 8'h0; 1: mux_25829 = vout_peek_8609;
    endcase
  endfunction
  wire [7:0] v_25830;
  function [7:0] mux_25830(input [0:0] sel);
    case (sel) 0: mux_25830 = 8'h0; 1: mux_25830 = vout_peek_8600;
    endcase
  endfunction
  wire [7:0] v_25831;
  function [7:0] mux_25831(input [0:0] sel);
    case (sel) 0: mux_25831 = 8'h0; 1: mux_25831 = v_25832;
    endcase
  endfunction
  reg [7:0] v_25832 = 8'h0;
  wire [7:0] v_25833;
  wire [7:0] v_25834;
  function [7:0] mux_25834(input [0:0] sel);
    case (sel) 0: mux_25834 = 8'h0; 1: mux_25834 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25835;
  wire [7:0] v_25836;
  wire [7:0] v_25837;
  function [7:0] mux_25837(input [0:0] sel);
    case (sel) 0: mux_25837 = 8'h0; 1: mux_25837 = vout_peek_8572;
    endcase
  endfunction
  wire [7:0] v_25838;
  function [7:0] mux_25838(input [0:0] sel);
    case (sel) 0: mux_25838 = 8'h0; 1: mux_25838 = vout_peek_8563;
    endcase
  endfunction
  wire [7:0] v_25839;
  function [7:0] mux_25839(input [0:0] sel);
    case (sel) 0: mux_25839 = 8'h0; 1: mux_25839 = v_25840;
    endcase
  endfunction
  reg [7:0] v_25840 = 8'h0;
  wire [7:0] v_25841;
  wire [7:0] v_25842;
  function [7:0] mux_25842(input [0:0] sel);
    case (sel) 0: mux_25842 = 8'h0; 1: mux_25842 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25843;
  wire [7:0] v_25844;
  wire [7:0] v_25845;
  function [7:0] mux_25845(input [0:0] sel);
    case (sel) 0: mux_25845 = 8'h0; 1: mux_25845 = v_25846;
    endcase
  endfunction
  reg [7:0] v_25846 = 8'h0;
  wire [7:0] v_25847;
  wire [7:0] v_25848;
  function [7:0] mux_25848(input [0:0] sel);
    case (sel) 0: mux_25848 = 8'h0; 1: mux_25848 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25849;
  wire [7:0] v_25850;
  wire [7:0] v_25851;
  function [7:0] mux_25851(input [0:0] sel);
    case (sel) 0: mux_25851 = 8'h0; 1: mux_25851 = vout_peek_8516;
    endcase
  endfunction
  wire [7:0] v_25852;
  function [7:0] mux_25852(input [0:0] sel);
    case (sel) 0: mux_25852 = 8'h0; 1: mux_25852 = vout_peek_8507;
    endcase
  endfunction
  wire [7:0] v_25853;
  function [7:0] mux_25853(input [0:0] sel);
    case (sel) 0: mux_25853 = 8'h0; 1: mux_25853 = v_25854;
    endcase
  endfunction
  reg [7:0] v_25854 = 8'h0;
  wire [7:0] v_25855;
  wire [7:0] v_25856;
  function [7:0] mux_25856(input [0:0] sel);
    case (sel) 0: mux_25856 = 8'h0; 1: mux_25856 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25857;
  wire [7:0] v_25858;
  wire [7:0] v_25859;
  function [7:0] mux_25859(input [0:0] sel);
    case (sel) 0: mux_25859 = 8'h0; 1: mux_25859 = vout_peek_8479;
    endcase
  endfunction
  wire [7:0] v_25860;
  function [7:0] mux_25860(input [0:0] sel);
    case (sel) 0: mux_25860 = 8'h0; 1: mux_25860 = vout_peek_8470;
    endcase
  endfunction
  wire [7:0] v_25861;
  function [7:0] mux_25861(input [0:0] sel);
    case (sel) 0: mux_25861 = 8'h0; 1: mux_25861 = v_25862;
    endcase
  endfunction
  reg [7:0] v_25862 = 8'h0;
  wire [7:0] v_25863;
  wire [7:0] v_25864;
  function [7:0] mux_25864(input [0:0] sel);
    case (sel) 0: mux_25864 = 8'h0; 1: mux_25864 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25865;
  wire [7:0] v_25866;
  wire [7:0] v_25867;
  function [7:0] mux_25867(input [0:0] sel);
    case (sel) 0: mux_25867 = 8'h0; 1: mux_25867 = v_25868;
    endcase
  endfunction
  reg [7:0] v_25868 = 8'h0;
  wire [7:0] v_25869;
  wire [7:0] v_25870;
  function [7:0] mux_25870(input [0:0] sel);
    case (sel) 0: mux_25870 = 8'h0; 1: mux_25870 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25871;
  wire [7:0] v_25872;
  wire [7:0] v_25873;
  function [7:0] mux_25873(input [0:0] sel);
    case (sel) 0: mux_25873 = 8'h0; 1: mux_25873 = v_25874;
    endcase
  endfunction
  reg [7:0] v_25874 = 8'h0;
  wire [7:0] v_25875;
  wire [7:0] v_25876;
  function [7:0] mux_25876(input [0:0] sel);
    case (sel) 0: mux_25876 = 8'h0; 1: mux_25876 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25877;
  wire [7:0] v_25878;
  wire [7:0] v_25879;
  function [7:0] mux_25879(input [0:0] sel);
    case (sel) 0: mux_25879 = 8'h0; 1: mux_25879 = v_25880;
    endcase
  endfunction
  reg [7:0] v_25880 = 8'h0;
  wire [7:0] v_25881;
  wire [7:0] v_25882;
  function [7:0] mux_25882(input [0:0] sel);
    case (sel) 0: mux_25882 = 8'h0; 1: mux_25882 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25883;
  wire [7:0] v_25884;
  wire [7:0] v_25885;
  function [7:0] mux_25885(input [0:0] sel);
    case (sel) 0: mux_25885 = 8'h0; 1: mux_25885 = vout_peek_8385;
    endcase
  endfunction
  wire [7:0] v_25886;
  function [7:0] mux_25886(input [0:0] sel);
    case (sel) 0: mux_25886 = 8'h0; 1: mux_25886 = vout_peek_8376;
    endcase
  endfunction
  wire [7:0] v_25887;
  function [7:0] mux_25887(input [0:0] sel);
    case (sel) 0: mux_25887 = 8'h0; 1: mux_25887 = v_25888;
    endcase
  endfunction
  reg [7:0] v_25888 = 8'h0;
  wire [7:0] v_25889;
  wire [7:0] v_25890;
  function [7:0] mux_25890(input [0:0] sel);
    case (sel) 0: mux_25890 = 8'h0; 1: mux_25890 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25891;
  wire [7:0] v_25892;
  wire [7:0] v_25893;
  function [7:0] mux_25893(input [0:0] sel);
    case (sel) 0: mux_25893 = 8'h0; 1: mux_25893 = vout_peek_8348;
    endcase
  endfunction
  wire [7:0] v_25894;
  function [7:0] mux_25894(input [0:0] sel);
    case (sel) 0: mux_25894 = 8'h0; 1: mux_25894 = vout_peek_8339;
    endcase
  endfunction
  wire [7:0] v_25895;
  function [7:0] mux_25895(input [0:0] sel);
    case (sel) 0: mux_25895 = 8'h0; 1: mux_25895 = v_25896;
    endcase
  endfunction
  reg [7:0] v_25896 = 8'h0;
  wire [7:0] v_25897;
  wire [7:0] v_25898;
  function [7:0] mux_25898(input [0:0] sel);
    case (sel) 0: mux_25898 = 8'h0; 1: mux_25898 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25899;
  wire [7:0] v_25900;
  wire [7:0] v_25901;
  function [7:0] mux_25901(input [0:0] sel);
    case (sel) 0: mux_25901 = 8'h0; 1: mux_25901 = v_25902;
    endcase
  endfunction
  reg [7:0] v_25902 = 8'h0;
  wire [7:0] v_25903;
  wire [7:0] v_25904;
  function [7:0] mux_25904(input [0:0] sel);
    case (sel) 0: mux_25904 = 8'h0; 1: mux_25904 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25905;
  wire [7:0] v_25906;
  wire [7:0] v_25907;
  function [7:0] mux_25907(input [0:0] sel);
    case (sel) 0: mux_25907 = 8'h0; 1: mux_25907 = vout_peek_8292;
    endcase
  endfunction
  wire [7:0] v_25908;
  function [7:0] mux_25908(input [0:0] sel);
    case (sel) 0: mux_25908 = 8'h0; 1: mux_25908 = vout_peek_8283;
    endcase
  endfunction
  wire [7:0] v_25909;
  function [7:0] mux_25909(input [0:0] sel);
    case (sel) 0: mux_25909 = 8'h0; 1: mux_25909 = v_25910;
    endcase
  endfunction
  reg [7:0] v_25910 = 8'h0;
  wire [7:0] v_25911;
  wire [7:0] v_25912;
  function [7:0] mux_25912(input [0:0] sel);
    case (sel) 0: mux_25912 = 8'h0; 1: mux_25912 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25913;
  wire [7:0] v_25914;
  wire [7:0] v_25915;
  function [7:0] mux_25915(input [0:0] sel);
    case (sel) 0: mux_25915 = 8'h0; 1: mux_25915 = vout_peek_8255;
    endcase
  endfunction
  wire [7:0] v_25916;
  function [7:0] mux_25916(input [0:0] sel);
    case (sel) 0: mux_25916 = 8'h0; 1: mux_25916 = vout_peek_8246;
    endcase
  endfunction
  wire [7:0] v_25917;
  function [7:0] mux_25917(input [0:0] sel);
    case (sel) 0: mux_25917 = 8'h0; 1: mux_25917 = v_25918;
    endcase
  endfunction
  reg [7:0] v_25918 = 8'h0;
  wire [7:0] v_25919;
  wire [7:0] v_25920;
  function [7:0] mux_25920(input [0:0] sel);
    case (sel) 0: mux_25920 = 8'h0; 1: mux_25920 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25921;
  wire [7:0] v_25922;
  wire [7:0] v_25923;
  function [7:0] mux_25923(input [0:0] sel);
    case (sel) 0: mux_25923 = 8'h0; 1: mux_25923 = v_25924;
    endcase
  endfunction
  reg [7:0] v_25924 = 8'h0;
  wire [7:0] v_25925;
  wire [7:0] v_25926;
  function [7:0] mux_25926(input [0:0] sel);
    case (sel) 0: mux_25926 = 8'h0; 1: mux_25926 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25927;
  wire [7:0] v_25928;
  wire [7:0] v_25929;
  function [7:0] mux_25929(input [0:0] sel);
    case (sel) 0: mux_25929 = 8'h0; 1: mux_25929 = v_25930;
    endcase
  endfunction
  reg [7:0] v_25930 = 8'h0;
  wire [7:0] v_25931;
  wire [7:0] v_25932;
  function [7:0] mux_25932(input [0:0] sel);
    case (sel) 0: mux_25932 = 8'h0; 1: mux_25932 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25933;
  wire [7:0] v_25934;
  wire [7:0] v_25935;
  function [7:0] mux_25935(input [0:0] sel);
    case (sel) 0: mux_25935 = 8'h0; 1: mux_25935 = vout_peek_8180;
    endcase
  endfunction
  wire [7:0] v_25936;
  function [7:0] mux_25936(input [0:0] sel);
    case (sel) 0: mux_25936 = 8'h0; 1: mux_25936 = vout_peek_8171;
    endcase
  endfunction
  wire [7:0] v_25937;
  function [7:0] mux_25937(input [0:0] sel);
    case (sel) 0: mux_25937 = 8'h0; 1: mux_25937 = v_25938;
    endcase
  endfunction
  reg [7:0] v_25938 = 8'h0;
  wire [7:0] v_25939;
  wire [7:0] v_25940;
  function [7:0] mux_25940(input [0:0] sel);
    case (sel) 0: mux_25940 = 8'h0; 1: mux_25940 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25941;
  wire [7:0] v_25942;
  wire [7:0] v_25943;
  function [7:0] mux_25943(input [0:0] sel);
    case (sel) 0: mux_25943 = 8'h0; 1: mux_25943 = vout_peek_8143;
    endcase
  endfunction
  wire [7:0] v_25944;
  function [7:0] mux_25944(input [0:0] sel);
    case (sel) 0: mux_25944 = 8'h0; 1: mux_25944 = vout_peek_8134;
    endcase
  endfunction
  wire [7:0] v_25945;
  function [7:0] mux_25945(input [0:0] sel);
    case (sel) 0: mux_25945 = 8'h0; 1: mux_25945 = v_25946;
    endcase
  endfunction
  reg [7:0] v_25946 = 8'h0;
  wire [7:0] v_25947;
  wire [7:0] v_25948;
  function [7:0] mux_25948(input [0:0] sel);
    case (sel) 0: mux_25948 = 8'h0; 1: mux_25948 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25949;
  wire [7:0] v_25950;
  wire [7:0] v_25951;
  function [7:0] mux_25951(input [0:0] sel);
    case (sel) 0: mux_25951 = 8'h0; 1: mux_25951 = v_25952;
    endcase
  endfunction
  reg [7:0] v_25952 = 8'h0;
  wire [7:0] v_25953;
  wire [7:0] v_25954;
  function [7:0] mux_25954(input [0:0] sel);
    case (sel) 0: mux_25954 = 8'h0; 1: mux_25954 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25955;
  wire [7:0] v_25956;
  wire [7:0] v_25957;
  function [7:0] mux_25957(input [0:0] sel);
    case (sel) 0: mux_25957 = 8'h0; 1: mux_25957 = vout_peek_8087;
    endcase
  endfunction
  wire [7:0] v_25958;
  function [7:0] mux_25958(input [0:0] sel);
    case (sel) 0: mux_25958 = 8'h0; 1: mux_25958 = vout_peek_8078;
    endcase
  endfunction
  wire [7:0] v_25959;
  function [7:0] mux_25959(input [0:0] sel);
    case (sel) 0: mux_25959 = 8'h0; 1: mux_25959 = v_25960;
    endcase
  endfunction
  reg [7:0] v_25960 = 8'h0;
  wire [7:0] v_25961;
  wire [7:0] v_25962;
  function [7:0] mux_25962(input [0:0] sel);
    case (sel) 0: mux_25962 = 8'h0; 1: mux_25962 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25963;
  wire [7:0] v_25964;
  wire [7:0] v_25965;
  function [7:0] mux_25965(input [0:0] sel);
    case (sel) 0: mux_25965 = 8'h0; 1: mux_25965 = vout_peek_8050;
    endcase
  endfunction
  wire [7:0] v_25966;
  function [7:0] mux_25966(input [0:0] sel);
    case (sel) 0: mux_25966 = 8'h0; 1: mux_25966 = vout_peek_8041;
    endcase
  endfunction
  wire [7:0] v_25967;
  function [7:0] mux_25967(input [0:0] sel);
    case (sel) 0: mux_25967 = 8'h0; 1: mux_25967 = v_25968;
    endcase
  endfunction
  reg [7:0] v_25968 = 8'h0;
  wire [7:0] v_25969;
  wire [7:0] v_25970;
  function [7:0] mux_25970(input [0:0] sel);
    case (sel) 0: mux_25970 = 8'h0; 1: mux_25970 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25971;
  wire [7:0] v_25972;
  wire [7:0] v_25973;
  function [7:0] mux_25973(input [0:0] sel);
    case (sel) 0: mux_25973 = 8'h0; 1: mux_25973 = v_25974;
    endcase
  endfunction
  reg [7:0] v_25974 = 8'h0;
  wire [7:0] v_25975;
  wire [7:0] v_25976;
  function [7:0] mux_25976(input [0:0] sel);
    case (sel) 0: mux_25976 = 8'h0; 1: mux_25976 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25977;
  wire [7:0] v_25978;
  wire [7:0] v_25979;
  function [7:0] mux_25979(input [0:0] sel);
    case (sel) 0: mux_25979 = 8'h0; 1: mux_25979 = v_25980;
    endcase
  endfunction
  reg [7:0] v_25980 = 8'h0;
  wire [7:0] v_25981;
  wire [7:0] v_25982;
  function [7:0] mux_25982(input [0:0] sel);
    case (sel) 0: mux_25982 = 8'h0; 1: mux_25982 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25983;
  wire [7:0] v_25984;
  wire [7:0] v_25985;
  function [7:0] mux_25985(input [0:0] sel);
    case (sel) 0: mux_25985 = 8'h0; 1: mux_25985 = v_25986;
    endcase
  endfunction
  reg [7:0] v_25986 = 8'h0;
  wire [7:0] v_25987;
  wire [7:0] v_25988;
  function [7:0] mux_25988(input [0:0] sel);
    case (sel) 0: mux_25988 = 8'h0; 1: mux_25988 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25989;
  wire [7:0] v_25990;
  wire [7:0] v_25991;
  function [7:0] mux_25991(input [0:0] sel);
    case (sel) 0: mux_25991 = 8'h0; 1: mux_25991 = v_25992;
    endcase
  endfunction
  reg [7:0] v_25992 = 8'h0;
  wire [7:0] v_25993;
  wire [7:0] v_25994;
  function [7:0] mux_25994(input [0:0] sel);
    case (sel) 0: mux_25994 = 8'h0; 1: mux_25994 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_25995;
  wire [7:0] v_25996;
  wire [7:0] v_25997;
  function [7:0] mux_25997(input [0:0] sel);
    case (sel) 0: mux_25997 = 8'h0; 1: mux_25997 = v_25998;
    endcase
  endfunction
  reg [7:0] v_25998 = 8'h0;
  wire [7:0] v_25999;
  wire [7:0] v_26000;
  function [7:0] mux_26000(input [0:0] sel);
    case (sel) 0: mux_26000 = 8'h0; 1: mux_26000 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26001;
  wire [7:0] v_26002;
  wire [7:0] v_26003;
  function [7:0] mux_26003(input [0:0] sel);
    case (sel) 0: mux_26003 = 8'h0; 1: mux_26003 = v_26004;
    endcase
  endfunction
  reg [7:0] v_26004 = 8'h0;
  wire [7:0] v_26005;
  wire [7:0] v_26006;
  function [7:0] mux_26006(input [0:0] sel);
    case (sel) 0: mux_26006 = 8'h0; 1: mux_26006 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26007;
  wire [7:0] v_26008;
  wire [7:0] v_26009;
  function [7:0] mux_26009(input [0:0] sel);
    case (sel) 0: mux_26009 = 8'h0; 1: mux_26009 = v_26010;
    endcase
  endfunction
  reg [7:0] v_26010 = 8'h0;
  wire [7:0] v_26011;
  wire [7:0] v_26012;
  function [7:0] mux_26012(input [0:0] sel);
    case (sel) 0: mux_26012 = 8'h0; 1: mux_26012 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26013;
  wire [7:0] v_26014;
  wire [7:0] v_26015;
  function [7:0] mux_26015(input [0:0] sel);
    case (sel) 0: mux_26015 = 8'h0; 1: mux_26015 = v_26016;
    endcase
  endfunction
  reg [7:0] v_26016 = 8'h0;
  wire [7:0] v_26017;
  wire [7:0] v_26018;
  function [7:0] mux_26018(input [0:0] sel);
    case (sel) 0: mux_26018 = 8'h0; 1: mux_26018 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26019;
  wire [7:0] v_26020;
  wire [7:0] v_26021;
  function [7:0] mux_26021(input [0:0] sel);
    case (sel) 0: mux_26021 = 8'h0; 1: mux_26021 = vout_peek_1660;
    endcase
  endfunction
  wire [7:0] v_26022;
  function [7:0] mux_26022(input [0:0] sel);
    case (sel) 0: mux_26022 = 8'h0; 1: mux_26022 = vout_peek_1651;
    endcase
  endfunction
  wire [7:0] v_26023;
  function [7:0] mux_26023(input [0:0] sel);
    case (sel) 0: mux_26023 = 8'h0; 1: mux_26023 = v_26024;
    endcase
  endfunction
  reg [7:0] v_26024 = 8'h0;
  wire [7:0] v_26025;
  wire [7:0] v_26026;
  function [7:0] mux_26026(input [0:0] sel);
    case (sel) 0: mux_26026 = 8'h0; 1: mux_26026 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26027;
  wire [7:0] v_26028;
  wire [7:0] v_26029;
  function [7:0] mux_26029(input [0:0] sel);
    case (sel) 0: mux_26029 = 8'h0; 1: mux_26029 = vout_peek_1623;
    endcase
  endfunction
  wire [7:0] v_26030;
  function [7:0] mux_26030(input [0:0] sel);
    case (sel) 0: mux_26030 = 8'h0; 1: mux_26030 = vout_peek_1614;
    endcase
  endfunction
  wire [7:0] v_26031;
  function [7:0] mux_26031(input [0:0] sel);
    case (sel) 0: mux_26031 = 8'h0; 1: mux_26031 = v_26032;
    endcase
  endfunction
  reg [7:0] v_26032 = 8'h0;
  wire [7:0] v_26033;
  wire [7:0] v_26034;
  function [7:0] mux_26034(input [0:0] sel);
    case (sel) 0: mux_26034 = 8'h0; 1: mux_26034 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26035;
  wire [7:0] v_26036;
  wire [7:0] v_26037;
  function [7:0] mux_26037(input [0:0] sel);
    case (sel) 0: mux_26037 = 8'h0; 1: mux_26037 = v_26038;
    endcase
  endfunction
  reg [7:0] v_26038 = 8'h0;
  wire [7:0] v_26039;
  wire [7:0] v_26040;
  function [7:0] mux_26040(input [0:0] sel);
    case (sel) 0: mux_26040 = 8'h0; 1: mux_26040 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26041;
  wire [7:0] v_26042;
  wire [7:0] v_26043;
  function [7:0] mux_26043(input [0:0] sel);
    case (sel) 0: mux_26043 = 8'h0; 1: mux_26043 = vout_peek_1567;
    endcase
  endfunction
  wire [7:0] v_26044;
  function [7:0] mux_26044(input [0:0] sel);
    case (sel) 0: mux_26044 = 8'h0; 1: mux_26044 = vout_peek_1558;
    endcase
  endfunction
  wire [7:0] v_26045;
  function [7:0] mux_26045(input [0:0] sel);
    case (sel) 0: mux_26045 = 8'h0; 1: mux_26045 = v_26046;
    endcase
  endfunction
  reg [7:0] v_26046 = 8'h0;
  wire [7:0] v_26047;
  wire [7:0] v_26048;
  function [7:0] mux_26048(input [0:0] sel);
    case (sel) 0: mux_26048 = 8'h0; 1: mux_26048 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26049;
  wire [7:0] v_26050;
  wire [7:0] v_26051;
  function [7:0] mux_26051(input [0:0] sel);
    case (sel) 0: mux_26051 = 8'h0; 1: mux_26051 = vout_peek_1530;
    endcase
  endfunction
  wire [7:0] v_26052;
  function [7:0] mux_26052(input [0:0] sel);
    case (sel) 0: mux_26052 = 8'h0; 1: mux_26052 = vout_peek_1521;
    endcase
  endfunction
  wire [7:0] v_26053;
  function [7:0] mux_26053(input [0:0] sel);
    case (sel) 0: mux_26053 = 8'h0; 1: mux_26053 = v_26054;
    endcase
  endfunction
  reg [7:0] v_26054 = 8'h0;
  wire [7:0] v_26055;
  wire [7:0] v_26056;
  function [7:0] mux_26056(input [0:0] sel);
    case (sel) 0: mux_26056 = 8'h0; 1: mux_26056 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26057;
  wire [7:0] v_26058;
  wire [7:0] v_26059;
  function [7:0] mux_26059(input [0:0] sel);
    case (sel) 0: mux_26059 = 8'h0; 1: mux_26059 = v_26060;
    endcase
  endfunction
  reg [7:0] v_26060 = 8'h0;
  wire [7:0] v_26061;
  wire [7:0] v_26062;
  function [7:0] mux_26062(input [0:0] sel);
    case (sel) 0: mux_26062 = 8'h0; 1: mux_26062 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26063;
  wire [7:0] v_26064;
  wire [7:0] v_26065;
  function [7:0] mux_26065(input [0:0] sel);
    case (sel) 0: mux_26065 = 8'h0; 1: mux_26065 = v_26066;
    endcase
  endfunction
  reg [7:0] v_26066 = 8'h0;
  wire [7:0] v_26067;
  wire [7:0] v_26068;
  function [7:0] mux_26068(input [0:0] sel);
    case (sel) 0: mux_26068 = 8'h0; 1: mux_26068 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26069;
  wire [7:0] v_26070;
  wire [7:0] v_26071;
  function [7:0] mux_26071(input [0:0] sel);
    case (sel) 0: mux_26071 = 8'h0; 1: mux_26071 = vout_peek_1455;
    endcase
  endfunction
  wire [7:0] v_26072;
  function [7:0] mux_26072(input [0:0] sel);
    case (sel) 0: mux_26072 = 8'h0; 1: mux_26072 = vout_peek_1446;
    endcase
  endfunction
  wire [7:0] v_26073;
  function [7:0] mux_26073(input [0:0] sel);
    case (sel) 0: mux_26073 = 8'h0; 1: mux_26073 = v_26074;
    endcase
  endfunction
  reg [7:0] v_26074 = 8'h0;
  wire [7:0] v_26075;
  wire [7:0] v_26076;
  function [7:0] mux_26076(input [0:0] sel);
    case (sel) 0: mux_26076 = 8'h0; 1: mux_26076 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26077;
  wire [7:0] v_26078;
  wire [7:0] v_26079;
  function [7:0] mux_26079(input [0:0] sel);
    case (sel) 0: mux_26079 = 8'h0; 1: mux_26079 = vout_peek_1418;
    endcase
  endfunction
  wire [7:0] v_26080;
  function [7:0] mux_26080(input [0:0] sel);
    case (sel) 0: mux_26080 = 8'h0; 1: mux_26080 = vout_peek_1409;
    endcase
  endfunction
  wire [7:0] v_26081;
  function [7:0] mux_26081(input [0:0] sel);
    case (sel) 0: mux_26081 = 8'h0; 1: mux_26081 = v_26082;
    endcase
  endfunction
  reg [7:0] v_26082 = 8'h0;
  wire [7:0] v_26083;
  wire [7:0] v_26084;
  function [7:0] mux_26084(input [0:0] sel);
    case (sel) 0: mux_26084 = 8'h0; 1: mux_26084 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26085;
  wire [7:0] v_26086;
  wire [7:0] v_26087;
  function [7:0] mux_26087(input [0:0] sel);
    case (sel) 0: mux_26087 = 8'h0; 1: mux_26087 = v_26088;
    endcase
  endfunction
  reg [7:0] v_26088 = 8'h0;
  wire [7:0] v_26089;
  wire [7:0] v_26090;
  function [7:0] mux_26090(input [0:0] sel);
    case (sel) 0: mux_26090 = 8'h0; 1: mux_26090 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26091;
  wire [7:0] v_26092;
  wire [7:0] v_26093;
  function [7:0] mux_26093(input [0:0] sel);
    case (sel) 0: mux_26093 = 8'h0; 1: mux_26093 = vout_peek_1362;
    endcase
  endfunction
  wire [7:0] v_26094;
  function [7:0] mux_26094(input [0:0] sel);
    case (sel) 0: mux_26094 = 8'h0; 1: mux_26094 = vout_peek_1353;
    endcase
  endfunction
  wire [7:0] v_26095;
  function [7:0] mux_26095(input [0:0] sel);
    case (sel) 0: mux_26095 = 8'h0; 1: mux_26095 = v_26096;
    endcase
  endfunction
  reg [7:0] v_26096 = 8'h0;
  wire [7:0] v_26097;
  wire [7:0] v_26098;
  function [7:0] mux_26098(input [0:0] sel);
    case (sel) 0: mux_26098 = 8'h0; 1: mux_26098 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26099;
  wire [7:0] v_26100;
  wire [7:0] v_26101;
  function [7:0] mux_26101(input [0:0] sel);
    case (sel) 0: mux_26101 = 8'h0; 1: mux_26101 = vout_peek_1325;
    endcase
  endfunction
  wire [7:0] v_26102;
  function [7:0] mux_26102(input [0:0] sel);
    case (sel) 0: mux_26102 = 8'h0; 1: mux_26102 = vout_peek_1316;
    endcase
  endfunction
  wire [7:0] v_26103;
  function [7:0] mux_26103(input [0:0] sel);
    case (sel) 0: mux_26103 = 8'h0; 1: mux_26103 = v_26104;
    endcase
  endfunction
  reg [7:0] v_26104 = 8'h0;
  wire [7:0] v_26105;
  wire [7:0] v_26106;
  function [7:0] mux_26106(input [0:0] sel);
    case (sel) 0: mux_26106 = 8'h0; 1: mux_26106 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26107;
  wire [7:0] v_26108;
  wire [7:0] v_26109;
  function [7:0] mux_26109(input [0:0] sel);
    case (sel) 0: mux_26109 = 8'h0; 1: mux_26109 = v_26110;
    endcase
  endfunction
  reg [7:0] v_26110 = 8'h0;
  wire [7:0] v_26111;
  wire [7:0] v_26112;
  function [7:0] mux_26112(input [0:0] sel);
    case (sel) 0: mux_26112 = 8'h0; 1: mux_26112 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26113;
  wire [7:0] v_26114;
  wire [7:0] v_26115;
  function [7:0] mux_26115(input [0:0] sel);
    case (sel) 0: mux_26115 = 8'h0; 1: mux_26115 = v_26116;
    endcase
  endfunction
  reg [7:0] v_26116 = 8'h0;
  wire [7:0] v_26117;
  wire [7:0] v_26118;
  function [7:0] mux_26118(input [0:0] sel);
    case (sel) 0: mux_26118 = 8'h0; 1: mux_26118 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26119;
  wire [7:0] v_26120;
  wire [7:0] v_26121;
  function [7:0] mux_26121(input [0:0] sel);
    case (sel) 0: mux_26121 = 8'h0; 1: mux_26121 = v_26122;
    endcase
  endfunction
  reg [7:0] v_26122 = 8'h0;
  wire [7:0] v_26123;
  wire [7:0] v_26124;
  function [7:0] mux_26124(input [0:0] sel);
    case (sel) 0: mux_26124 = 8'h0; 1: mux_26124 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26125;
  wire [7:0] v_26126;
  wire [7:0] v_26127;
  function [7:0] mux_26127(input [0:0] sel);
    case (sel) 0: mux_26127 = 8'h0; 1: mux_26127 = vout_peek_1231;
    endcase
  endfunction
  wire [7:0] v_26128;
  function [7:0] mux_26128(input [0:0] sel);
    case (sel) 0: mux_26128 = 8'h0; 1: mux_26128 = vout_peek_1222;
    endcase
  endfunction
  wire [7:0] v_26129;
  function [7:0] mux_26129(input [0:0] sel);
    case (sel) 0: mux_26129 = 8'h0; 1: mux_26129 = v_26130;
    endcase
  endfunction
  reg [7:0] v_26130 = 8'h0;
  wire [7:0] v_26131;
  wire [7:0] v_26132;
  function [7:0] mux_26132(input [0:0] sel);
    case (sel) 0: mux_26132 = 8'h0; 1: mux_26132 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26133;
  wire [7:0] v_26134;
  wire [7:0] v_26135;
  function [7:0] mux_26135(input [0:0] sel);
    case (sel) 0: mux_26135 = 8'h0; 1: mux_26135 = vout_peek_1194;
    endcase
  endfunction
  wire [7:0] v_26136;
  function [7:0] mux_26136(input [0:0] sel);
    case (sel) 0: mux_26136 = 8'h0; 1: mux_26136 = vout_peek_1185;
    endcase
  endfunction
  wire [7:0] v_26137;
  function [7:0] mux_26137(input [0:0] sel);
    case (sel) 0: mux_26137 = 8'h0; 1: mux_26137 = v_26138;
    endcase
  endfunction
  reg [7:0] v_26138 = 8'h0;
  wire [7:0] v_26139;
  wire [7:0] v_26140;
  function [7:0] mux_26140(input [0:0] sel);
    case (sel) 0: mux_26140 = 8'h0; 1: mux_26140 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26141;
  wire [7:0] v_26142;
  wire [7:0] v_26143;
  function [7:0] mux_26143(input [0:0] sel);
    case (sel) 0: mux_26143 = 8'h0; 1: mux_26143 = v_26144;
    endcase
  endfunction
  reg [7:0] v_26144 = 8'h0;
  wire [7:0] v_26145;
  wire [7:0] v_26146;
  function [7:0] mux_26146(input [0:0] sel);
    case (sel) 0: mux_26146 = 8'h0; 1: mux_26146 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26147;
  wire [7:0] v_26148;
  wire [7:0] v_26149;
  function [7:0] mux_26149(input [0:0] sel);
    case (sel) 0: mux_26149 = 8'h0; 1: mux_26149 = vout_peek_1138;
    endcase
  endfunction
  wire [7:0] v_26150;
  function [7:0] mux_26150(input [0:0] sel);
    case (sel) 0: mux_26150 = 8'h0; 1: mux_26150 = vout_peek_1129;
    endcase
  endfunction
  wire [7:0] v_26151;
  function [7:0] mux_26151(input [0:0] sel);
    case (sel) 0: mux_26151 = 8'h0; 1: mux_26151 = v_26152;
    endcase
  endfunction
  reg [7:0] v_26152 = 8'h0;
  wire [7:0] v_26153;
  wire [7:0] v_26154;
  function [7:0] mux_26154(input [0:0] sel);
    case (sel) 0: mux_26154 = 8'h0; 1: mux_26154 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26155;
  wire [7:0] v_26156;
  wire [7:0] v_26157;
  function [7:0] mux_26157(input [0:0] sel);
    case (sel) 0: mux_26157 = 8'h0; 1: mux_26157 = vout_peek_1101;
    endcase
  endfunction
  wire [7:0] v_26158;
  function [7:0] mux_26158(input [0:0] sel);
    case (sel) 0: mux_26158 = 8'h0; 1: mux_26158 = vout_peek_1092;
    endcase
  endfunction
  wire [7:0] v_26159;
  function [7:0] mux_26159(input [0:0] sel);
    case (sel) 0: mux_26159 = 8'h0; 1: mux_26159 = v_26160;
    endcase
  endfunction
  reg [7:0] v_26160 = 8'h0;
  wire [7:0] v_26161;
  wire [7:0] v_26162;
  function [7:0] mux_26162(input [0:0] sel);
    case (sel) 0: mux_26162 = 8'h0; 1: mux_26162 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26163;
  wire [7:0] v_26164;
  wire [7:0] v_26165;
  function [7:0] mux_26165(input [0:0] sel);
    case (sel) 0: mux_26165 = 8'h0; 1: mux_26165 = v_26166;
    endcase
  endfunction
  reg [7:0] v_26166 = 8'h0;
  wire [7:0] v_26167;
  wire [7:0] v_26168;
  function [7:0] mux_26168(input [0:0] sel);
    case (sel) 0: mux_26168 = 8'h0; 1: mux_26168 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26169;
  wire [7:0] v_26170;
  wire [7:0] v_26171;
  function [7:0] mux_26171(input [0:0] sel);
    case (sel) 0: mux_26171 = 8'h0; 1: mux_26171 = v_26172;
    endcase
  endfunction
  reg [7:0] v_26172 = 8'h0;
  wire [7:0] v_26173;
  wire [7:0] v_26174;
  function [7:0] mux_26174(input [0:0] sel);
    case (sel) 0: mux_26174 = 8'h0; 1: mux_26174 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26175;
  wire [7:0] v_26176;
  wire [7:0] v_26177;
  function [7:0] mux_26177(input [0:0] sel);
    case (sel) 0: mux_26177 = 8'h0; 1: mux_26177 = vout_peek_1026;
    endcase
  endfunction
  wire [7:0] v_26178;
  function [7:0] mux_26178(input [0:0] sel);
    case (sel) 0: mux_26178 = 8'h0; 1: mux_26178 = vout_peek_1017;
    endcase
  endfunction
  wire [7:0] v_26179;
  function [7:0] mux_26179(input [0:0] sel);
    case (sel) 0: mux_26179 = 8'h0; 1: mux_26179 = v_26180;
    endcase
  endfunction
  reg [7:0] v_26180 = 8'h0;
  wire [7:0] v_26181;
  wire [7:0] v_26182;
  function [7:0] mux_26182(input [0:0] sel);
    case (sel) 0: mux_26182 = 8'h0; 1: mux_26182 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26183;
  wire [7:0] v_26184;
  wire [7:0] v_26185;
  function [7:0] mux_26185(input [0:0] sel);
    case (sel) 0: mux_26185 = 8'h0; 1: mux_26185 = vout_peek_989;
    endcase
  endfunction
  wire [7:0] v_26186;
  function [7:0] mux_26186(input [0:0] sel);
    case (sel) 0: mux_26186 = 8'h0; 1: mux_26186 = vout_peek_980;
    endcase
  endfunction
  wire [7:0] v_26187;
  function [7:0] mux_26187(input [0:0] sel);
    case (sel) 0: mux_26187 = 8'h0; 1: mux_26187 = v_26188;
    endcase
  endfunction
  reg [7:0] v_26188 = 8'h0;
  wire [7:0] v_26189;
  wire [7:0] v_26190;
  function [7:0] mux_26190(input [0:0] sel);
    case (sel) 0: mux_26190 = 8'h0; 1: mux_26190 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26191;
  wire [7:0] v_26192;
  wire [7:0] v_26193;
  function [7:0] mux_26193(input [0:0] sel);
    case (sel) 0: mux_26193 = 8'h0; 1: mux_26193 = v_26194;
    endcase
  endfunction
  reg [7:0] v_26194 = 8'h0;
  wire [7:0] v_26195;
  wire [7:0] v_26196;
  function [7:0] mux_26196(input [0:0] sel);
    case (sel) 0: mux_26196 = 8'h0; 1: mux_26196 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26197;
  wire [7:0] v_26198;
  wire [7:0] v_26199;
  function [7:0] mux_26199(input [0:0] sel);
    case (sel) 0: mux_26199 = 8'h0; 1: mux_26199 = vout_peek_933;
    endcase
  endfunction
  wire [7:0] v_26200;
  function [7:0] mux_26200(input [0:0] sel);
    case (sel) 0: mux_26200 = 8'h0; 1: mux_26200 = vout_peek_924;
    endcase
  endfunction
  wire [7:0] v_26201;
  function [7:0] mux_26201(input [0:0] sel);
    case (sel) 0: mux_26201 = 8'h0; 1: mux_26201 = v_26202;
    endcase
  endfunction
  reg [7:0] v_26202 = 8'h0;
  wire [7:0] v_26203;
  wire [7:0] v_26204;
  function [7:0] mux_26204(input [0:0] sel);
    case (sel) 0: mux_26204 = 8'h0; 1: mux_26204 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26205;
  wire [7:0] v_26206;
  wire [7:0] v_26207;
  function [7:0] mux_26207(input [0:0] sel);
    case (sel) 0: mux_26207 = 8'h0; 1: mux_26207 = vout_peek_896;
    endcase
  endfunction
  wire [7:0] v_26208;
  function [7:0] mux_26208(input [0:0] sel);
    case (sel) 0: mux_26208 = 8'h0; 1: mux_26208 = vout_peek_887;
    endcase
  endfunction
  wire [7:0] v_26209;
  function [7:0] mux_26209(input [0:0] sel);
    case (sel) 0: mux_26209 = 8'h0; 1: mux_26209 = v_26210;
    endcase
  endfunction
  reg [7:0] v_26210 = 8'h0;
  wire [7:0] v_26211;
  wire [7:0] v_26212;
  function [7:0] mux_26212(input [0:0] sel);
    case (sel) 0: mux_26212 = 8'h0; 1: mux_26212 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26213;
  wire [7:0] v_26214;
  wire [7:0] v_26215;
  function [7:0] mux_26215(input [0:0] sel);
    case (sel) 0: mux_26215 = 8'h0; 1: mux_26215 = v_26216;
    endcase
  endfunction
  reg [7:0] v_26216 = 8'h0;
  wire [7:0] v_26217;
  wire [7:0] v_26218;
  function [7:0] mux_26218(input [0:0] sel);
    case (sel) 0: mux_26218 = 8'h0; 1: mux_26218 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26219;
  wire [7:0] v_26220;
  wire [7:0] v_26221;
  function [7:0] mux_26221(input [0:0] sel);
    case (sel) 0: mux_26221 = 8'h0; 1: mux_26221 = v_26222;
    endcase
  endfunction
  reg [7:0] v_26222 = 8'h0;
  wire [7:0] v_26223;
  wire [7:0] v_26224;
  function [7:0] mux_26224(input [0:0] sel);
    case (sel) 0: mux_26224 = 8'h0; 1: mux_26224 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26225;
  wire [7:0] v_26226;
  wire [7:0] v_26227;
  function [7:0] mux_26227(input [0:0] sel);
    case (sel) 0: mux_26227 = 8'h0; 1: mux_26227 = v_26228;
    endcase
  endfunction
  reg [7:0] v_26228 = 8'h0;
  wire [7:0] v_26229;
  wire [7:0] v_26230;
  function [7:0] mux_26230(input [0:0] sel);
    case (sel) 0: mux_26230 = 8'h0; 1: mux_26230 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26231;
  wire [7:0] v_26232;
  wire [7:0] v_26233;
  function [7:0] mux_26233(input [0:0] sel);
    case (sel) 0: mux_26233 = 8'h0; 1: mux_26233 = v_26234;
    endcase
  endfunction
  reg [7:0] v_26234 = 8'h0;
  wire [7:0] v_26235;
  wire [7:0] v_26236;
  function [7:0] mux_26236(input [0:0] sel);
    case (sel) 0: mux_26236 = 8'h0; 1: mux_26236 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26237;
  wire [7:0] v_26238;
  wire [7:0] v_26239;
  function [7:0] mux_26239(input [0:0] sel);
    case (sel) 0: mux_26239 = 8'h0; 1: mux_26239 = vout_peek_782;
    endcase
  endfunction
  wire [7:0] v_26240;
  function [7:0] mux_26240(input [0:0] sel);
    case (sel) 0: mux_26240 = 8'h0; 1: mux_26240 = vout_peek_773;
    endcase
  endfunction
  wire [7:0] v_26241;
  function [7:0] mux_26241(input [0:0] sel);
    case (sel) 0: mux_26241 = 8'h0; 1: mux_26241 = v_26242;
    endcase
  endfunction
  reg [7:0] v_26242 = 8'h0;
  wire [7:0] v_26243;
  wire [7:0] v_26244;
  function [7:0] mux_26244(input [0:0] sel);
    case (sel) 0: mux_26244 = 8'h0; 1: mux_26244 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26245;
  wire [7:0] v_26246;
  wire [7:0] v_26247;
  function [7:0] mux_26247(input [0:0] sel);
    case (sel) 0: mux_26247 = 8'h0; 1: mux_26247 = vout_peek_745;
    endcase
  endfunction
  wire [7:0] v_26248;
  function [7:0] mux_26248(input [0:0] sel);
    case (sel) 0: mux_26248 = 8'h0; 1: mux_26248 = vout_peek_736;
    endcase
  endfunction
  wire [7:0] v_26249;
  function [7:0] mux_26249(input [0:0] sel);
    case (sel) 0: mux_26249 = 8'h0; 1: mux_26249 = v_26250;
    endcase
  endfunction
  reg [7:0] v_26250 = 8'h0;
  wire [7:0] v_26251;
  wire [7:0] v_26252;
  function [7:0] mux_26252(input [0:0] sel);
    case (sel) 0: mux_26252 = 8'h0; 1: mux_26252 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26253;
  wire [7:0] v_26254;
  wire [7:0] v_26255;
  function [7:0] mux_26255(input [0:0] sel);
    case (sel) 0: mux_26255 = 8'h0; 1: mux_26255 = v_26256;
    endcase
  endfunction
  reg [7:0] v_26256 = 8'h0;
  wire [7:0] v_26257;
  wire [7:0] v_26258;
  function [7:0] mux_26258(input [0:0] sel);
    case (sel) 0: mux_26258 = 8'h0; 1: mux_26258 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26259;
  wire [7:0] v_26260;
  wire [7:0] v_26261;
  function [7:0] mux_26261(input [0:0] sel);
    case (sel) 0: mux_26261 = 8'h0; 1: mux_26261 = vout_peek_689;
    endcase
  endfunction
  wire [7:0] v_26262;
  function [7:0] mux_26262(input [0:0] sel);
    case (sel) 0: mux_26262 = 8'h0; 1: mux_26262 = vout_peek_680;
    endcase
  endfunction
  wire [7:0] v_26263;
  function [7:0] mux_26263(input [0:0] sel);
    case (sel) 0: mux_26263 = 8'h0; 1: mux_26263 = v_26264;
    endcase
  endfunction
  reg [7:0] v_26264 = 8'h0;
  wire [7:0] v_26265;
  wire [7:0] v_26266;
  function [7:0] mux_26266(input [0:0] sel);
    case (sel) 0: mux_26266 = 8'h0; 1: mux_26266 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26267;
  wire [7:0] v_26268;
  wire [7:0] v_26269;
  function [7:0] mux_26269(input [0:0] sel);
    case (sel) 0: mux_26269 = 8'h0; 1: mux_26269 = vout_peek_652;
    endcase
  endfunction
  wire [7:0] v_26270;
  function [7:0] mux_26270(input [0:0] sel);
    case (sel) 0: mux_26270 = 8'h0; 1: mux_26270 = vout_peek_643;
    endcase
  endfunction
  wire [7:0] v_26271;
  function [7:0] mux_26271(input [0:0] sel);
    case (sel) 0: mux_26271 = 8'h0; 1: mux_26271 = v_26272;
    endcase
  endfunction
  reg [7:0] v_26272 = 8'h0;
  wire [7:0] v_26273;
  wire [7:0] v_26274;
  function [7:0] mux_26274(input [0:0] sel);
    case (sel) 0: mux_26274 = 8'h0; 1: mux_26274 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26275;
  wire [7:0] v_26276;
  wire [7:0] v_26277;
  function [7:0] mux_26277(input [0:0] sel);
    case (sel) 0: mux_26277 = 8'h0; 1: mux_26277 = v_26278;
    endcase
  endfunction
  reg [7:0] v_26278 = 8'h0;
  wire [7:0] v_26279;
  wire [7:0] v_26280;
  function [7:0] mux_26280(input [0:0] sel);
    case (sel) 0: mux_26280 = 8'h0; 1: mux_26280 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26281;
  wire [7:0] v_26282;
  wire [7:0] v_26283;
  function [7:0] mux_26283(input [0:0] sel);
    case (sel) 0: mux_26283 = 8'h0; 1: mux_26283 = v_26284;
    endcase
  endfunction
  reg [7:0] v_26284 = 8'h0;
  wire [7:0] v_26285;
  wire [7:0] v_26286;
  function [7:0] mux_26286(input [0:0] sel);
    case (sel) 0: mux_26286 = 8'h0; 1: mux_26286 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26287;
  wire [7:0] v_26288;
  wire [7:0] v_26289;
  function [7:0] mux_26289(input [0:0] sel);
    case (sel) 0: mux_26289 = 8'h0; 1: mux_26289 = vout_peek_577;
    endcase
  endfunction
  wire [7:0] v_26290;
  function [7:0] mux_26290(input [0:0] sel);
    case (sel) 0: mux_26290 = 8'h0; 1: mux_26290 = vout_peek_568;
    endcase
  endfunction
  wire [7:0] v_26291;
  function [7:0] mux_26291(input [0:0] sel);
    case (sel) 0: mux_26291 = 8'h0; 1: mux_26291 = v_26292;
    endcase
  endfunction
  reg [7:0] v_26292 = 8'h0;
  wire [7:0] v_26293;
  wire [7:0] v_26294;
  function [7:0] mux_26294(input [0:0] sel);
    case (sel) 0: mux_26294 = 8'h0; 1: mux_26294 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26295;
  wire [7:0] v_26296;
  wire [7:0] v_26297;
  function [7:0] mux_26297(input [0:0] sel);
    case (sel) 0: mux_26297 = 8'h0; 1: mux_26297 = vout_peek_540;
    endcase
  endfunction
  wire [7:0] v_26298;
  function [7:0] mux_26298(input [0:0] sel);
    case (sel) 0: mux_26298 = 8'h0; 1: mux_26298 = vout_peek_531;
    endcase
  endfunction
  wire [7:0] v_26299;
  function [7:0] mux_26299(input [0:0] sel);
    case (sel) 0: mux_26299 = 8'h0; 1: mux_26299 = v_26300;
    endcase
  endfunction
  reg [7:0] v_26300 = 8'h0;
  wire [7:0] v_26301;
  wire [7:0] v_26302;
  function [7:0] mux_26302(input [0:0] sel);
    case (sel) 0: mux_26302 = 8'h0; 1: mux_26302 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26303;
  wire [7:0] v_26304;
  wire [7:0] v_26305;
  function [7:0] mux_26305(input [0:0] sel);
    case (sel) 0: mux_26305 = 8'h0; 1: mux_26305 = v_26306;
    endcase
  endfunction
  reg [7:0] v_26306 = 8'h0;
  wire [7:0] v_26307;
  wire [7:0] v_26308;
  function [7:0] mux_26308(input [0:0] sel);
    case (sel) 0: mux_26308 = 8'h0; 1: mux_26308 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26309;
  wire [7:0] v_26310;
  wire [7:0] v_26311;
  function [7:0] mux_26311(input [0:0] sel);
    case (sel) 0: mux_26311 = 8'h0; 1: mux_26311 = vout_peek_484;
    endcase
  endfunction
  wire [7:0] v_26312;
  function [7:0] mux_26312(input [0:0] sel);
    case (sel) 0: mux_26312 = 8'h0; 1: mux_26312 = vout_peek_475;
    endcase
  endfunction
  wire [7:0] v_26313;
  function [7:0] mux_26313(input [0:0] sel);
    case (sel) 0: mux_26313 = 8'h0; 1: mux_26313 = v_26314;
    endcase
  endfunction
  reg [7:0] v_26314 = 8'h0;
  wire [7:0] v_26315;
  wire [7:0] v_26316;
  function [7:0] mux_26316(input [0:0] sel);
    case (sel) 0: mux_26316 = 8'h0; 1: mux_26316 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26317;
  wire [7:0] v_26318;
  wire [7:0] v_26319;
  function [7:0] mux_26319(input [0:0] sel);
    case (sel) 0: mux_26319 = 8'h0; 1: mux_26319 = vout_peek_447;
    endcase
  endfunction
  wire [7:0] v_26320;
  function [7:0] mux_26320(input [0:0] sel);
    case (sel) 0: mux_26320 = 8'h0; 1: mux_26320 = vout_peek_438;
    endcase
  endfunction
  wire [7:0] v_26321;
  function [7:0] mux_26321(input [0:0] sel);
    case (sel) 0: mux_26321 = 8'h0; 1: mux_26321 = v_26322;
    endcase
  endfunction
  reg [7:0] v_26322 = 8'h0;
  wire [7:0] v_26323;
  wire [7:0] v_26324;
  function [7:0] mux_26324(input [0:0] sel);
    case (sel) 0: mux_26324 = 8'h0; 1: mux_26324 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26325;
  wire [7:0] v_26326;
  wire [7:0] v_26327;
  function [7:0] mux_26327(input [0:0] sel);
    case (sel) 0: mux_26327 = 8'h0; 1: mux_26327 = v_26328;
    endcase
  endfunction
  reg [7:0] v_26328 = 8'h0;
  wire [7:0] v_26329;
  wire [7:0] v_26330;
  function [7:0] mux_26330(input [0:0] sel);
    case (sel) 0: mux_26330 = 8'h0; 1: mux_26330 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26331;
  wire [7:0] v_26332;
  wire [7:0] v_26333;
  function [7:0] mux_26333(input [0:0] sel);
    case (sel) 0: mux_26333 = 8'h0; 1: mux_26333 = v_26334;
    endcase
  endfunction
  reg [7:0] v_26334 = 8'h0;
  wire [7:0] v_26335;
  wire [7:0] v_26336;
  function [7:0] mux_26336(input [0:0] sel);
    case (sel) 0: mux_26336 = 8'h0; 1: mux_26336 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26337;
  wire [7:0] v_26338;
  wire [7:0] v_26339;
  function [7:0] mux_26339(input [0:0] sel);
    case (sel) 0: mux_26339 = 8'h0; 1: mux_26339 = v_26340;
    endcase
  endfunction
  reg [7:0] v_26340 = 8'h0;
  wire [7:0] v_26341;
  wire [7:0] v_26342;
  function [7:0] mux_26342(input [0:0] sel);
    case (sel) 0: mux_26342 = 8'h0; 1: mux_26342 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26343;
  wire [7:0] v_26344;
  wire [7:0] v_26345;
  function [7:0] mux_26345(input [0:0] sel);
    case (sel) 0: mux_26345 = 8'h0; 1: mux_26345 = vout_peek_352;
    endcase
  endfunction
  wire [7:0] v_26346;
  function [7:0] mux_26346(input [0:0] sel);
    case (sel) 0: mux_26346 = 8'h0; 1: mux_26346 = vout_peek_343;
    endcase
  endfunction
  wire [7:0] v_26347;
  function [7:0] mux_26347(input [0:0] sel);
    case (sel) 0: mux_26347 = 8'h0; 1: mux_26347 = v_26348;
    endcase
  endfunction
  reg [7:0] v_26348 = 8'h0;
  wire [7:0] v_26349;
  wire [7:0] v_26350;
  function [7:0] mux_26350(input [0:0] sel);
    case (sel) 0: mux_26350 = 8'h0; 1: mux_26350 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26351;
  wire [7:0] v_26352;
  wire [7:0] v_26353;
  function [7:0] mux_26353(input [0:0] sel);
    case (sel) 0: mux_26353 = 8'h0; 1: mux_26353 = vout_peek_315;
    endcase
  endfunction
  wire [7:0] v_26354;
  function [7:0] mux_26354(input [0:0] sel);
    case (sel) 0: mux_26354 = 8'h0; 1: mux_26354 = vout_peek_306;
    endcase
  endfunction
  wire [7:0] v_26355;
  function [7:0] mux_26355(input [0:0] sel);
    case (sel) 0: mux_26355 = 8'h0; 1: mux_26355 = v_26356;
    endcase
  endfunction
  reg [7:0] v_26356 = 8'h0;
  wire [7:0] v_26357;
  wire [7:0] v_26358;
  function [7:0] mux_26358(input [0:0] sel);
    case (sel) 0: mux_26358 = 8'h0; 1: mux_26358 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26359;
  wire [7:0] v_26360;
  wire [7:0] v_26361;
  function [7:0] mux_26361(input [0:0] sel);
    case (sel) 0: mux_26361 = 8'h0; 1: mux_26361 = v_26362;
    endcase
  endfunction
  reg [7:0] v_26362 = 8'h0;
  wire [7:0] v_26363;
  wire [7:0] v_26364;
  function [7:0] mux_26364(input [0:0] sel);
    case (sel) 0: mux_26364 = 8'h0; 1: mux_26364 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26365;
  wire [7:0] v_26366;
  wire [7:0] v_26367;
  function [7:0] mux_26367(input [0:0] sel);
    case (sel) 0: mux_26367 = 8'h0; 1: mux_26367 = vout_peek_259;
    endcase
  endfunction
  wire [7:0] v_26368;
  function [7:0] mux_26368(input [0:0] sel);
    case (sel) 0: mux_26368 = 8'h0; 1: mux_26368 = vout_peek_250;
    endcase
  endfunction
  wire [7:0] v_26369;
  function [7:0] mux_26369(input [0:0] sel);
    case (sel) 0: mux_26369 = 8'h0; 1: mux_26369 = v_26370;
    endcase
  endfunction
  reg [7:0] v_26370 = 8'h0;
  wire [7:0] v_26371;
  wire [7:0] v_26372;
  function [7:0] mux_26372(input [0:0] sel);
    case (sel) 0: mux_26372 = 8'h0; 1: mux_26372 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26373;
  wire [7:0] v_26374;
  wire [7:0] v_26375;
  function [7:0] mux_26375(input [0:0] sel);
    case (sel) 0: mux_26375 = 8'h0; 1: mux_26375 = vout_peek_222;
    endcase
  endfunction
  wire [7:0] v_26376;
  function [7:0] mux_26376(input [0:0] sel);
    case (sel) 0: mux_26376 = 8'h0; 1: mux_26376 = vout_peek_213;
    endcase
  endfunction
  wire [7:0] v_26377;
  function [7:0] mux_26377(input [0:0] sel);
    case (sel) 0: mux_26377 = 8'h0; 1: mux_26377 = v_26378;
    endcase
  endfunction
  reg [7:0] v_26378 = 8'h0;
  wire [7:0] v_26379;
  wire [7:0] v_26380;
  function [7:0] mux_26380(input [0:0] sel);
    case (sel) 0: mux_26380 = 8'h0; 1: mux_26380 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26381;
  wire [7:0] v_26382;
  wire [7:0] v_26383;
  function [7:0] mux_26383(input [0:0] sel);
    case (sel) 0: mux_26383 = 8'h0; 1: mux_26383 = v_26384;
    endcase
  endfunction
  reg [7:0] v_26384 = 8'h0;
  wire [7:0] v_26385;
  wire [7:0] v_26386;
  function [7:0] mux_26386(input [0:0] sel);
    case (sel) 0: mux_26386 = 8'h0; 1: mux_26386 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26387;
  wire [7:0] v_26388;
  wire [7:0] v_26389;
  function [7:0] mux_26389(input [0:0] sel);
    case (sel) 0: mux_26389 = 8'h0; 1: mux_26389 = v_26390;
    endcase
  endfunction
  reg [7:0] v_26390 = 8'h0;
  wire [7:0] v_26391;
  wire [7:0] v_26392;
  function [7:0] mux_26392(input [0:0] sel);
    case (sel) 0: mux_26392 = 8'h0; 1: mux_26392 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26393;
  wire [7:0] v_26394;
  wire [7:0] v_26395;
  function [7:0] mux_26395(input [0:0] sel);
    case (sel) 0: mux_26395 = 8'h0; 1: mux_26395 = vout_peek_146;
    endcase
  endfunction
  wire [7:0] v_26396;
  function [7:0] mux_26396(input [0:0] sel);
    case (sel) 0: mux_26396 = 8'h0; 1: mux_26396 = vout_peek_137;
    endcase
  endfunction
  wire [7:0] v_26397;
  function [7:0] mux_26397(input [0:0] sel);
    case (sel) 0: mux_26397 = 8'h0; 1: mux_26397 = v_26398;
    endcase
  endfunction
  reg [7:0] v_26398 = 8'h0;
  wire [7:0] v_26399;
  wire [7:0] v_26400;
  function [7:0] mux_26400(input [0:0] sel);
    case (sel) 0: mux_26400 = 8'h0; 1: mux_26400 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26401;
  wire [7:0] v_26402;
  wire [7:0] v_26403;
  function [7:0] mux_26403(input [0:0] sel);
    case (sel) 0: mux_26403 = 8'h0; 1: mux_26403 = vout_peek_109;
    endcase
  endfunction
  wire [7:0] v_26404;
  function [7:0] mux_26404(input [0:0] sel);
    case (sel) 0: mux_26404 = 8'h0; 1: mux_26404 = vout_peek_100;
    endcase
  endfunction
  wire [7:0] v_26405;
  function [7:0] mux_26405(input [0:0] sel);
    case (sel) 0: mux_26405 = 8'h0; 1: mux_26405 = v_26406;
    endcase
  endfunction
  reg [7:0] v_26406 = 8'h0;
  wire [7:0] v_26407;
  wire [7:0] v_26408;
  function [7:0] mux_26408(input [0:0] sel);
    case (sel) 0: mux_26408 = 8'h0; 1: mux_26408 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26409;
  wire [7:0] v_26410;
  wire [7:0] v_26411;
  function [7:0] mux_26411(input [0:0] sel);
    case (sel) 0: mux_26411 = 8'h0; 1: mux_26411 = v_26412;
    endcase
  endfunction
  reg [7:0] v_26412 = 8'h0;
  wire [7:0] v_26413;
  wire [7:0] v_26414;
  function [7:0] mux_26414(input [0:0] sel);
    case (sel) 0: mux_26414 = 8'h0; 1: mux_26414 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26415;
  wire [7:0] v_26416;
  wire [7:0] v_26417;
  function [7:0] mux_26417(input [0:0] sel);
    case (sel) 0: mux_26417 = 8'h0; 1: mux_26417 = vout_peek_52;
    endcase
  endfunction
  wire [7:0] v_26418;
  function [7:0] mux_26418(input [0:0] sel);
    case (sel) 0: mux_26418 = 8'h0; 1: mux_26418 = vout_peek_43;
    endcase
  endfunction
  wire [7:0] v_26419;
  function [7:0] mux_26419(input [0:0] sel);
    case (sel) 0: mux_26419 = 8'h0; 1: mux_26419 = v_26420;
    endcase
  endfunction
  reg [7:0] v_26420 = 8'h0;
  wire [7:0] v_26421;
  wire [7:0] v_26422;
  function [7:0] mux_26422(input [0:0] sel);
    case (sel) 0: mux_26422 = 8'h0; 1: mux_26422 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26423;
  wire [7:0] v_26424;
  wire [7:0] v_26425;
  function [7:0] mux_26425(input [0:0] sel);
    case (sel) 0: mux_26425 = 8'h0; 1: mux_26425 = vout_peek_14;
    endcase
  endfunction
  wire [7:0] v_26426;
  function [7:0] mux_26426(input [0:0] sel);
    case (sel) 0: mux_26426 = 8'h0; 1: mux_26426 = vout_peek_3;
    endcase
  endfunction
  wire [7:0] v_26427;
  function [7:0] mux_26427(input [0:0] sel);
    case (sel) 0: mux_26427 = 8'h0; 1: mux_26427 = v_26428;
    endcase
  endfunction
  reg [7:0] v_26428 = 8'h0;
  wire [7:0] v_26429;
  wire [7:0] v_26430;
  function [7:0] mux_26430(input [0:0] sel);
    case (sel) 0: mux_26430 = 8'h0; 1: mux_26430 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26431;
  wire [7:0] v_26432;
  wire [7:0] v_26433;
  function [7:0] mux_26433(input [0:0] sel);
    case (sel) 0: mux_26433 = 8'h0; 1: mux_26433 = v_26434;
    endcase
  endfunction
  reg [7:0] v_26434 = 8'h0;
  wire [7:0] v_26435;
  wire [7:0] v_26436;
  function [7:0] mux_26436(input [0:0] sel);
    case (sel) 0: mux_26436 = 8'h0; 1: mux_26436 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26437;
  wire [7:0] v_26438;
  wire [7:0] v_26439;
  function [7:0] mux_26439(input [0:0] sel);
    case (sel) 0: mux_26439 = 8'h0; 1: mux_26439 = v_26440;
    endcase
  endfunction
  reg [7:0] v_26440 = 8'h0;
  wire [7:0] v_26441;
  wire [7:0] v_26442;
  function [7:0] mux_26442(input [0:0] sel);
    case (sel) 0: mux_26442 = 8'h0; 1: mux_26442 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26443;
  wire [7:0] v_26444;
  wire [7:0] v_26445;
  function [7:0] mux_26445(input [0:0] sel);
    case (sel) 0: mux_26445 = 8'h0; 1: mux_26445 = v_26446;
    endcase
  endfunction
  reg [7:0] v_26446 = 8'h0;
  wire [7:0] v_26447;
  wire [7:0] v_26448;
  function [7:0] mux_26448(input [0:0] sel);
    case (sel) 0: mux_26448 = 8'h0; 1: mux_26448 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26449;
  wire [7:0] v_26450;
  wire [7:0] v_26451;
  function [7:0] mux_26451(input [0:0] sel);
    case (sel) 0: mux_26451 = 8'h0; 1: mux_26451 = v_26452;
    endcase
  endfunction
  reg [7:0] v_26452 = 8'h0;
  wire [7:0] v_26453;
  wire [7:0] v_26454;
  function [7:0] mux_26454(input [0:0] sel);
    case (sel) 0: mux_26454 = 8'h0; 1: mux_26454 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26455;
  wire [7:0] v_26456;
  wire [7:0] v_26457;
  function [7:0] mux_26457(input [0:0] sel);
    case (sel) 0: mux_26457 = 8'h0; 1: mux_26457 = vout_peek_2542;
    endcase
  endfunction
  wire [7:0] v_26458;
  function [7:0] mux_26458(input [0:0] sel);
    case (sel) 0: mux_26458 = 8'h0; 1: mux_26458 = vout_peek_2533;
    endcase
  endfunction
  wire [7:0] v_26459;
  function [7:0] mux_26459(input [0:0] sel);
    case (sel) 0: mux_26459 = 8'h0; 1: mux_26459 = v_26460;
    endcase
  endfunction
  reg [7:0] v_26460 = 8'h0;
  wire [7:0] v_26461;
  wire [7:0] v_26462;
  function [7:0] mux_26462(input [0:0] sel);
    case (sel) 0: mux_26462 = 8'h0; 1: mux_26462 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26463;
  wire [7:0] v_26464;
  wire [7:0] v_26465;
  function [7:0] mux_26465(input [0:0] sel);
    case (sel) 0: mux_26465 = 8'h0; 1: mux_26465 = vout_peek_2505;
    endcase
  endfunction
  wire [7:0] v_26466;
  function [7:0] mux_26466(input [0:0] sel);
    case (sel) 0: mux_26466 = 8'h0; 1: mux_26466 = vout_peek_2496;
    endcase
  endfunction
  wire [7:0] v_26467;
  function [7:0] mux_26467(input [0:0] sel);
    case (sel) 0: mux_26467 = 8'h0; 1: mux_26467 = v_26468;
    endcase
  endfunction
  reg [7:0] v_26468 = 8'h0;
  wire [7:0] v_26469;
  wire [7:0] v_26470;
  function [7:0] mux_26470(input [0:0] sel);
    case (sel) 0: mux_26470 = 8'h0; 1: mux_26470 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26471;
  wire [7:0] v_26472;
  wire [7:0] v_26473;
  function [7:0] mux_26473(input [0:0] sel);
    case (sel) 0: mux_26473 = 8'h0; 1: mux_26473 = v_26474;
    endcase
  endfunction
  reg [7:0] v_26474 = 8'h0;
  wire [7:0] v_26475;
  wire [7:0] v_26476;
  function [7:0] mux_26476(input [0:0] sel);
    case (sel) 0: mux_26476 = 8'h0; 1: mux_26476 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26477;
  wire [7:0] v_26478;
  wire [7:0] v_26479;
  function [7:0] mux_26479(input [0:0] sel);
    case (sel) 0: mux_26479 = 8'h0; 1: mux_26479 = vout_peek_2449;
    endcase
  endfunction
  wire [7:0] v_26480;
  function [7:0] mux_26480(input [0:0] sel);
    case (sel) 0: mux_26480 = 8'h0; 1: mux_26480 = vout_peek_2440;
    endcase
  endfunction
  wire [7:0] v_26481;
  function [7:0] mux_26481(input [0:0] sel);
    case (sel) 0: mux_26481 = 8'h0; 1: mux_26481 = v_26482;
    endcase
  endfunction
  reg [7:0] v_26482 = 8'h0;
  wire [7:0] v_26483;
  wire [7:0] v_26484;
  function [7:0] mux_26484(input [0:0] sel);
    case (sel) 0: mux_26484 = 8'h0; 1: mux_26484 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26485;
  wire [7:0] v_26486;
  wire [7:0] v_26487;
  function [7:0] mux_26487(input [0:0] sel);
    case (sel) 0: mux_26487 = 8'h0; 1: mux_26487 = vout_peek_2412;
    endcase
  endfunction
  wire [7:0] v_26488;
  function [7:0] mux_26488(input [0:0] sel);
    case (sel) 0: mux_26488 = 8'h0; 1: mux_26488 = vout_peek_2403;
    endcase
  endfunction
  wire [7:0] v_26489;
  function [7:0] mux_26489(input [0:0] sel);
    case (sel) 0: mux_26489 = 8'h0; 1: mux_26489 = v_26490;
    endcase
  endfunction
  reg [7:0] v_26490 = 8'h0;
  wire [7:0] v_26491;
  wire [7:0] v_26492;
  function [7:0] mux_26492(input [0:0] sel);
    case (sel) 0: mux_26492 = 8'h0; 1: mux_26492 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26493;
  wire [7:0] v_26494;
  wire [7:0] v_26495;
  function [7:0] mux_26495(input [0:0] sel);
    case (sel) 0: mux_26495 = 8'h0; 1: mux_26495 = v_26496;
    endcase
  endfunction
  reg [7:0] v_26496 = 8'h0;
  wire [7:0] v_26497;
  wire [7:0] v_26498;
  function [7:0] mux_26498(input [0:0] sel);
    case (sel) 0: mux_26498 = 8'h0; 1: mux_26498 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26499;
  wire [7:0] v_26500;
  wire [7:0] v_26501;
  function [7:0] mux_26501(input [0:0] sel);
    case (sel) 0: mux_26501 = 8'h0; 1: mux_26501 = v_26502;
    endcase
  endfunction
  reg [7:0] v_26502 = 8'h0;
  wire [7:0] v_26503;
  wire [7:0] v_26504;
  function [7:0] mux_26504(input [0:0] sel);
    case (sel) 0: mux_26504 = 8'h0; 1: mux_26504 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26505;
  wire [7:0] v_26506;
  wire [7:0] v_26507;
  function [7:0] mux_26507(input [0:0] sel);
    case (sel) 0: mux_26507 = 8'h0; 1: mux_26507 = vout_peek_2337;
    endcase
  endfunction
  wire [7:0] v_26508;
  function [7:0] mux_26508(input [0:0] sel);
    case (sel) 0: mux_26508 = 8'h0; 1: mux_26508 = vout_peek_2328;
    endcase
  endfunction
  wire [7:0] v_26509;
  function [7:0] mux_26509(input [0:0] sel);
    case (sel) 0: mux_26509 = 8'h0; 1: mux_26509 = v_26510;
    endcase
  endfunction
  reg [7:0] v_26510 = 8'h0;
  wire [7:0] v_26511;
  wire [7:0] v_26512;
  function [7:0] mux_26512(input [0:0] sel);
    case (sel) 0: mux_26512 = 8'h0; 1: mux_26512 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26513;
  wire [7:0] v_26514;
  wire [7:0] v_26515;
  function [7:0] mux_26515(input [0:0] sel);
    case (sel) 0: mux_26515 = 8'h0; 1: mux_26515 = vout_peek_2300;
    endcase
  endfunction
  wire [7:0] v_26516;
  function [7:0] mux_26516(input [0:0] sel);
    case (sel) 0: mux_26516 = 8'h0; 1: mux_26516 = vout_peek_2291;
    endcase
  endfunction
  wire [7:0] v_26517;
  function [7:0] mux_26517(input [0:0] sel);
    case (sel) 0: mux_26517 = 8'h0; 1: mux_26517 = v_26518;
    endcase
  endfunction
  reg [7:0] v_26518 = 8'h0;
  wire [7:0] v_26519;
  wire [7:0] v_26520;
  function [7:0] mux_26520(input [0:0] sel);
    case (sel) 0: mux_26520 = 8'h0; 1: mux_26520 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26521;
  wire [7:0] v_26522;
  wire [7:0] v_26523;
  function [7:0] mux_26523(input [0:0] sel);
    case (sel) 0: mux_26523 = 8'h0; 1: mux_26523 = v_26524;
    endcase
  endfunction
  reg [7:0] v_26524 = 8'h0;
  wire [7:0] v_26525;
  wire [7:0] v_26526;
  function [7:0] mux_26526(input [0:0] sel);
    case (sel) 0: mux_26526 = 8'h0; 1: mux_26526 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26527;
  wire [7:0] v_26528;
  wire [7:0] v_26529;
  function [7:0] mux_26529(input [0:0] sel);
    case (sel) 0: mux_26529 = 8'h0; 1: mux_26529 = vout_peek_2244;
    endcase
  endfunction
  wire [7:0] v_26530;
  function [7:0] mux_26530(input [0:0] sel);
    case (sel) 0: mux_26530 = 8'h0; 1: mux_26530 = vout_peek_2235;
    endcase
  endfunction
  wire [7:0] v_26531;
  function [7:0] mux_26531(input [0:0] sel);
    case (sel) 0: mux_26531 = 8'h0; 1: mux_26531 = v_26532;
    endcase
  endfunction
  reg [7:0] v_26532 = 8'h0;
  wire [7:0] v_26533;
  wire [7:0] v_26534;
  function [7:0] mux_26534(input [0:0] sel);
    case (sel) 0: mux_26534 = 8'h0; 1: mux_26534 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26535;
  wire [7:0] v_26536;
  wire [7:0] v_26537;
  function [7:0] mux_26537(input [0:0] sel);
    case (sel) 0: mux_26537 = 8'h0; 1: mux_26537 = vout_peek_2207;
    endcase
  endfunction
  wire [7:0] v_26538;
  function [7:0] mux_26538(input [0:0] sel);
    case (sel) 0: mux_26538 = 8'h0; 1: mux_26538 = vout_peek_2198;
    endcase
  endfunction
  wire [7:0] v_26539;
  function [7:0] mux_26539(input [0:0] sel);
    case (sel) 0: mux_26539 = 8'h0; 1: mux_26539 = v_26540;
    endcase
  endfunction
  reg [7:0] v_26540 = 8'h0;
  wire [7:0] v_26541;
  wire [7:0] v_26542;
  function [7:0] mux_26542(input [0:0] sel);
    case (sel) 0: mux_26542 = 8'h0; 1: mux_26542 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26543;
  wire [7:0] v_26544;
  wire [7:0] v_26545;
  function [7:0] mux_26545(input [0:0] sel);
    case (sel) 0: mux_26545 = 8'h0; 1: mux_26545 = v_26546;
    endcase
  endfunction
  reg [7:0] v_26546 = 8'h0;
  wire [7:0] v_26547;
  wire [7:0] v_26548;
  function [7:0] mux_26548(input [0:0] sel);
    case (sel) 0: mux_26548 = 8'h0; 1: mux_26548 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26549;
  wire [7:0] v_26550;
  wire [7:0] v_26551;
  function [7:0] mux_26551(input [0:0] sel);
    case (sel) 0: mux_26551 = 8'h0; 1: mux_26551 = v_26552;
    endcase
  endfunction
  reg [7:0] v_26552 = 8'h0;
  wire [7:0] v_26553;
  wire [7:0] v_26554;
  function [7:0] mux_26554(input [0:0] sel);
    case (sel) 0: mux_26554 = 8'h0; 1: mux_26554 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26555;
  wire [7:0] v_26556;
  wire [7:0] v_26557;
  function [7:0] mux_26557(input [0:0] sel);
    case (sel) 0: mux_26557 = 8'h0; 1: mux_26557 = v_26558;
    endcase
  endfunction
  reg [7:0] v_26558 = 8'h0;
  wire [7:0] v_26559;
  wire [7:0] v_26560;
  function [7:0] mux_26560(input [0:0] sel);
    case (sel) 0: mux_26560 = 8'h0; 1: mux_26560 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26561;
  wire [7:0] v_26562;
  wire [7:0] v_26563;
  function [7:0] mux_26563(input [0:0] sel);
    case (sel) 0: mux_26563 = 8'h0; 1: mux_26563 = vout_peek_2113;
    endcase
  endfunction
  wire [7:0] v_26564;
  function [7:0] mux_26564(input [0:0] sel);
    case (sel) 0: mux_26564 = 8'h0; 1: mux_26564 = vout_peek_2104;
    endcase
  endfunction
  wire [7:0] v_26565;
  function [7:0] mux_26565(input [0:0] sel);
    case (sel) 0: mux_26565 = 8'h0; 1: mux_26565 = v_26566;
    endcase
  endfunction
  reg [7:0] v_26566 = 8'h0;
  wire [7:0] v_26567;
  wire [7:0] v_26568;
  function [7:0] mux_26568(input [0:0] sel);
    case (sel) 0: mux_26568 = 8'h0; 1: mux_26568 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26569;
  wire [7:0] v_26570;
  wire [7:0] v_26571;
  function [7:0] mux_26571(input [0:0] sel);
    case (sel) 0: mux_26571 = 8'h0; 1: mux_26571 = vout_peek_2076;
    endcase
  endfunction
  wire [7:0] v_26572;
  function [7:0] mux_26572(input [0:0] sel);
    case (sel) 0: mux_26572 = 8'h0; 1: mux_26572 = vout_peek_2067;
    endcase
  endfunction
  wire [7:0] v_26573;
  function [7:0] mux_26573(input [0:0] sel);
    case (sel) 0: mux_26573 = 8'h0; 1: mux_26573 = v_26574;
    endcase
  endfunction
  reg [7:0] v_26574 = 8'h0;
  wire [7:0] v_26575;
  wire [7:0] v_26576;
  function [7:0] mux_26576(input [0:0] sel);
    case (sel) 0: mux_26576 = 8'h0; 1: mux_26576 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26577;
  wire [7:0] v_26578;
  wire [7:0] v_26579;
  function [7:0] mux_26579(input [0:0] sel);
    case (sel) 0: mux_26579 = 8'h0; 1: mux_26579 = v_26580;
    endcase
  endfunction
  reg [7:0] v_26580 = 8'h0;
  wire [7:0] v_26581;
  wire [7:0] v_26582;
  function [7:0] mux_26582(input [0:0] sel);
    case (sel) 0: mux_26582 = 8'h0; 1: mux_26582 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26583;
  wire [7:0] v_26584;
  wire [7:0] v_26585;
  function [7:0] mux_26585(input [0:0] sel);
    case (sel) 0: mux_26585 = 8'h0; 1: mux_26585 = vout_peek_2020;
    endcase
  endfunction
  wire [7:0] v_26586;
  function [7:0] mux_26586(input [0:0] sel);
    case (sel) 0: mux_26586 = 8'h0; 1: mux_26586 = vout_peek_2011;
    endcase
  endfunction
  wire [7:0] v_26587;
  function [7:0] mux_26587(input [0:0] sel);
    case (sel) 0: mux_26587 = 8'h0; 1: mux_26587 = v_26588;
    endcase
  endfunction
  reg [7:0] v_26588 = 8'h0;
  wire [7:0] v_26589;
  wire [7:0] v_26590;
  function [7:0] mux_26590(input [0:0] sel);
    case (sel) 0: mux_26590 = 8'h0; 1: mux_26590 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26591;
  wire [7:0] v_26592;
  wire [7:0] v_26593;
  function [7:0] mux_26593(input [0:0] sel);
    case (sel) 0: mux_26593 = 8'h0; 1: mux_26593 = vout_peek_1983;
    endcase
  endfunction
  wire [7:0] v_26594;
  function [7:0] mux_26594(input [0:0] sel);
    case (sel) 0: mux_26594 = 8'h0; 1: mux_26594 = vout_peek_1974;
    endcase
  endfunction
  wire [7:0] v_26595;
  function [7:0] mux_26595(input [0:0] sel);
    case (sel) 0: mux_26595 = 8'h0; 1: mux_26595 = v_26596;
    endcase
  endfunction
  reg [7:0] v_26596 = 8'h0;
  wire [7:0] v_26597;
  wire [7:0] v_26598;
  function [7:0] mux_26598(input [0:0] sel);
    case (sel) 0: mux_26598 = 8'h0; 1: mux_26598 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26599;
  wire [7:0] v_26600;
  wire [7:0] v_26601;
  function [7:0] mux_26601(input [0:0] sel);
    case (sel) 0: mux_26601 = 8'h0; 1: mux_26601 = v_26602;
    endcase
  endfunction
  reg [7:0] v_26602 = 8'h0;
  wire [7:0] v_26603;
  wire [7:0] v_26604;
  function [7:0] mux_26604(input [0:0] sel);
    case (sel) 0: mux_26604 = 8'h0; 1: mux_26604 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26605;
  wire [7:0] v_26606;
  wire [7:0] v_26607;
  function [7:0] mux_26607(input [0:0] sel);
    case (sel) 0: mux_26607 = 8'h0; 1: mux_26607 = v_26608;
    endcase
  endfunction
  reg [7:0] v_26608 = 8'h0;
  wire [7:0] v_26609;
  wire [7:0] v_26610;
  function [7:0] mux_26610(input [0:0] sel);
    case (sel) 0: mux_26610 = 8'h0; 1: mux_26610 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26611;
  wire [7:0] v_26612;
  wire [7:0] v_26613;
  function [7:0] mux_26613(input [0:0] sel);
    case (sel) 0: mux_26613 = 8'h0; 1: mux_26613 = vout_peek_1908;
    endcase
  endfunction
  wire [7:0] v_26614;
  function [7:0] mux_26614(input [0:0] sel);
    case (sel) 0: mux_26614 = 8'h0; 1: mux_26614 = vout_peek_1899;
    endcase
  endfunction
  wire [7:0] v_26615;
  function [7:0] mux_26615(input [0:0] sel);
    case (sel) 0: mux_26615 = 8'h0; 1: mux_26615 = v_26616;
    endcase
  endfunction
  reg [7:0] v_26616 = 8'h0;
  wire [7:0] v_26617;
  wire [7:0] v_26618;
  function [7:0] mux_26618(input [0:0] sel);
    case (sel) 0: mux_26618 = 8'h0; 1: mux_26618 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26619;
  wire [7:0] v_26620;
  wire [7:0] v_26621;
  function [7:0] mux_26621(input [0:0] sel);
    case (sel) 0: mux_26621 = 8'h0; 1: mux_26621 = vout_peek_1871;
    endcase
  endfunction
  wire [7:0] v_26622;
  function [7:0] mux_26622(input [0:0] sel);
    case (sel) 0: mux_26622 = 8'h0; 1: mux_26622 = vout_peek_1862;
    endcase
  endfunction
  wire [7:0] v_26623;
  function [7:0] mux_26623(input [0:0] sel);
    case (sel) 0: mux_26623 = 8'h0; 1: mux_26623 = v_26624;
    endcase
  endfunction
  reg [7:0] v_26624 = 8'h0;
  wire [7:0] v_26625;
  wire [7:0] v_26626;
  function [7:0] mux_26626(input [0:0] sel);
    case (sel) 0: mux_26626 = 8'h0; 1: mux_26626 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26627;
  wire [7:0] v_26628;
  wire [7:0] v_26629;
  function [7:0] mux_26629(input [0:0] sel);
    case (sel) 0: mux_26629 = 8'h0; 1: mux_26629 = v_26630;
    endcase
  endfunction
  reg [7:0] v_26630 = 8'h0;
  wire [7:0] v_26631;
  wire [7:0] v_26632;
  function [7:0] mux_26632(input [0:0] sel);
    case (sel) 0: mux_26632 = 8'h0; 1: mux_26632 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26633;
  wire [7:0] v_26634;
  wire [7:0] v_26635;
  function [7:0] mux_26635(input [0:0] sel);
    case (sel) 0: mux_26635 = 8'h0; 1: mux_26635 = vout_peek_1815;
    endcase
  endfunction
  wire [7:0] v_26636;
  function [7:0] mux_26636(input [0:0] sel);
    case (sel) 0: mux_26636 = 8'h0; 1: mux_26636 = vout_peek_1806;
    endcase
  endfunction
  wire [7:0] v_26637;
  function [7:0] mux_26637(input [0:0] sel);
    case (sel) 0: mux_26637 = 8'h0; 1: mux_26637 = v_26638;
    endcase
  endfunction
  reg [7:0] v_26638 = 8'h0;
  wire [7:0] v_26639;
  wire [7:0] v_26640;
  function [7:0] mux_26640(input [0:0] sel);
    case (sel) 0: mux_26640 = 8'h0; 1: mux_26640 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26641;
  wire [7:0] v_26642;
  wire [7:0] v_26643;
  function [7:0] mux_26643(input [0:0] sel);
    case (sel) 0: mux_26643 = 8'h0; 1: mux_26643 = vout_peek_1778;
    endcase
  endfunction
  wire [7:0] v_26644;
  function [7:0] mux_26644(input [0:0] sel);
    case (sel) 0: mux_26644 = 8'h0; 1: mux_26644 = vout_peek_1769;
    endcase
  endfunction
  wire [7:0] v_26645;
  function [7:0] mux_26645(input [0:0] sel);
    case (sel) 0: mux_26645 = 8'h0; 1: mux_26645 = v_26646;
    endcase
  endfunction
  reg [7:0] v_26646 = 8'h0;
  wire [7:0] v_26647;
  wire [7:0] v_26648;
  function [7:0] mux_26648(input [0:0] sel);
    case (sel) 0: mux_26648 = 8'h0; 1: mux_26648 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26649;
  wire [7:0] v_26650;
  wire [7:0] v_26651;
  function [7:0] mux_26651(input [0:0] sel);
    case (sel) 0: mux_26651 = 8'h0; 1: mux_26651 = v_26652;
    endcase
  endfunction
  reg [7:0] v_26652 = 8'h0;
  wire [7:0] v_26653;
  wire [7:0] v_26654;
  function [7:0] mux_26654(input [0:0] sel);
    case (sel) 0: mux_26654 = 8'h0; 1: mux_26654 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26655;
  wire [7:0] v_26656;
  wire [7:0] v_26657;
  function [7:0] mux_26657(input [0:0] sel);
    case (sel) 0: mux_26657 = 8'h0; 1: mux_26657 = v_26658;
    endcase
  endfunction
  reg [7:0] v_26658 = 8'h0;
  wire [7:0] v_26659;
  wire [7:0] v_26660;
  function [7:0] mux_26660(input [0:0] sel);
    case (sel) 0: mux_26660 = 8'h0; 1: mux_26660 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26661;
  wire [7:0] v_26662;
  wire [7:0] v_26663;
  function [7:0] mux_26663(input [0:0] sel);
    case (sel) 0: mux_26663 = 8'h0; 1: mux_26663 = v_26664;
    endcase
  endfunction
  reg [7:0] v_26664 = 8'h0;
  wire [7:0] v_26665;
  wire [7:0] v_26666;
  function [7:0] mux_26666(input [0:0] sel);
    case (sel) 0: mux_26666 = 8'h0; 1: mux_26666 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26667;
  wire [7:0] v_26668;
  wire [7:0] v_26669;
  function [7:0] mux_26669(input [0:0] sel);
    case (sel) 0: mux_26669 = 8'h0; 1: mux_26669 = v_26670;
    endcase
  endfunction
  reg [7:0] v_26670 = 8'h0;
  wire [7:0] v_26671;
  wire [7:0] v_26672;
  function [7:0] mux_26672(input [0:0] sel);
    case (sel) 0: mux_26672 = 8'h0; 1: mux_26672 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26673;
  wire [7:0] v_26674;
  wire [7:0] v_26675;
  function [7:0] mux_26675(input [0:0] sel);
    case (sel) 0: mux_26675 = 8'h0; 1: mux_26675 = v_26676;
    endcase
  endfunction
  reg [7:0] v_26676 = 8'h0;
  wire [7:0] v_26677;
  wire [7:0] v_26678;
  function [7:0] mux_26678(input [0:0] sel);
    case (sel) 0: mux_26678 = 8'h0; 1: mux_26678 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26679;
  wire [7:0] v_26680;
  wire [7:0] v_26681;
  function [7:0] mux_26681(input [0:0] sel);
    case (sel) 0: mux_26681 = 8'h0; 1: mux_26681 = vout_peek_4310;
    endcase
  endfunction
  wire [7:0] v_26682;
  function [7:0] mux_26682(input [0:0] sel);
    case (sel) 0: mux_26682 = 8'h0; 1: mux_26682 = vout_peek_4301;
    endcase
  endfunction
  wire [7:0] v_26683;
  function [7:0] mux_26683(input [0:0] sel);
    case (sel) 0: mux_26683 = 8'h0; 1: mux_26683 = v_26684;
    endcase
  endfunction
  reg [7:0] v_26684 = 8'h0;
  wire [7:0] v_26685;
  wire [7:0] v_26686;
  function [7:0] mux_26686(input [0:0] sel);
    case (sel) 0: mux_26686 = 8'h0; 1: mux_26686 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26687;
  wire [7:0] v_26688;
  wire [7:0] v_26689;
  function [7:0] mux_26689(input [0:0] sel);
    case (sel) 0: mux_26689 = 8'h0; 1: mux_26689 = vout_peek_4273;
    endcase
  endfunction
  wire [7:0] v_26690;
  function [7:0] mux_26690(input [0:0] sel);
    case (sel) 0: mux_26690 = 8'h0; 1: mux_26690 = vout_peek_4264;
    endcase
  endfunction
  wire [7:0] v_26691;
  function [7:0] mux_26691(input [0:0] sel);
    case (sel) 0: mux_26691 = 8'h0; 1: mux_26691 = v_26692;
    endcase
  endfunction
  reg [7:0] v_26692 = 8'h0;
  wire [7:0] v_26693;
  wire [7:0] v_26694;
  function [7:0] mux_26694(input [0:0] sel);
    case (sel) 0: mux_26694 = 8'h0; 1: mux_26694 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26695;
  wire [7:0] v_26696;
  wire [7:0] v_26697;
  function [7:0] mux_26697(input [0:0] sel);
    case (sel) 0: mux_26697 = 8'h0; 1: mux_26697 = v_26698;
    endcase
  endfunction
  reg [7:0] v_26698 = 8'h0;
  wire [7:0] v_26699;
  wire [7:0] v_26700;
  function [7:0] mux_26700(input [0:0] sel);
    case (sel) 0: mux_26700 = 8'h0; 1: mux_26700 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26701;
  wire [7:0] v_26702;
  wire [7:0] v_26703;
  function [7:0] mux_26703(input [0:0] sel);
    case (sel) 0: mux_26703 = 8'h0; 1: mux_26703 = vout_peek_4217;
    endcase
  endfunction
  wire [7:0] v_26704;
  function [7:0] mux_26704(input [0:0] sel);
    case (sel) 0: mux_26704 = 8'h0; 1: mux_26704 = vout_peek_4208;
    endcase
  endfunction
  wire [7:0] v_26705;
  function [7:0] mux_26705(input [0:0] sel);
    case (sel) 0: mux_26705 = 8'h0; 1: mux_26705 = v_26706;
    endcase
  endfunction
  reg [7:0] v_26706 = 8'h0;
  wire [7:0] v_26707;
  wire [7:0] v_26708;
  function [7:0] mux_26708(input [0:0] sel);
    case (sel) 0: mux_26708 = 8'h0; 1: mux_26708 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26709;
  wire [7:0] v_26710;
  wire [7:0] v_26711;
  function [7:0] mux_26711(input [0:0] sel);
    case (sel) 0: mux_26711 = 8'h0; 1: mux_26711 = vout_peek_4180;
    endcase
  endfunction
  wire [7:0] v_26712;
  function [7:0] mux_26712(input [0:0] sel);
    case (sel) 0: mux_26712 = 8'h0; 1: mux_26712 = vout_peek_4171;
    endcase
  endfunction
  wire [7:0] v_26713;
  function [7:0] mux_26713(input [0:0] sel);
    case (sel) 0: mux_26713 = 8'h0; 1: mux_26713 = v_26714;
    endcase
  endfunction
  reg [7:0] v_26714 = 8'h0;
  wire [7:0] v_26715;
  wire [7:0] v_26716;
  function [7:0] mux_26716(input [0:0] sel);
    case (sel) 0: mux_26716 = 8'h0; 1: mux_26716 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26717;
  wire [7:0] v_26718;
  wire [7:0] v_26719;
  function [7:0] mux_26719(input [0:0] sel);
    case (sel) 0: mux_26719 = 8'h0; 1: mux_26719 = v_26720;
    endcase
  endfunction
  reg [7:0] v_26720 = 8'h0;
  wire [7:0] v_26721;
  wire [7:0] v_26722;
  function [7:0] mux_26722(input [0:0] sel);
    case (sel) 0: mux_26722 = 8'h0; 1: mux_26722 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26723;
  wire [7:0] v_26724;
  wire [7:0] v_26725;
  function [7:0] mux_26725(input [0:0] sel);
    case (sel) 0: mux_26725 = 8'h0; 1: mux_26725 = v_26726;
    endcase
  endfunction
  reg [7:0] v_26726 = 8'h0;
  wire [7:0] v_26727;
  wire [7:0] v_26728;
  function [7:0] mux_26728(input [0:0] sel);
    case (sel) 0: mux_26728 = 8'h0; 1: mux_26728 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26729;
  wire [7:0] v_26730;
  wire [7:0] v_26731;
  function [7:0] mux_26731(input [0:0] sel);
    case (sel) 0: mux_26731 = 8'h0; 1: mux_26731 = vout_peek_4105;
    endcase
  endfunction
  wire [7:0] v_26732;
  function [7:0] mux_26732(input [0:0] sel);
    case (sel) 0: mux_26732 = 8'h0; 1: mux_26732 = vout_peek_4096;
    endcase
  endfunction
  wire [7:0] v_26733;
  function [7:0] mux_26733(input [0:0] sel);
    case (sel) 0: mux_26733 = 8'h0; 1: mux_26733 = v_26734;
    endcase
  endfunction
  reg [7:0] v_26734 = 8'h0;
  wire [7:0] v_26735;
  wire [7:0] v_26736;
  function [7:0] mux_26736(input [0:0] sel);
    case (sel) 0: mux_26736 = 8'h0; 1: mux_26736 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26737;
  wire [7:0] v_26738;
  wire [7:0] v_26739;
  function [7:0] mux_26739(input [0:0] sel);
    case (sel) 0: mux_26739 = 8'h0; 1: mux_26739 = vout_peek_4068;
    endcase
  endfunction
  wire [7:0] v_26740;
  function [7:0] mux_26740(input [0:0] sel);
    case (sel) 0: mux_26740 = 8'h0; 1: mux_26740 = vout_peek_4059;
    endcase
  endfunction
  wire [7:0] v_26741;
  function [7:0] mux_26741(input [0:0] sel);
    case (sel) 0: mux_26741 = 8'h0; 1: mux_26741 = v_26742;
    endcase
  endfunction
  reg [7:0] v_26742 = 8'h0;
  wire [7:0] v_26743;
  wire [7:0] v_26744;
  function [7:0] mux_26744(input [0:0] sel);
    case (sel) 0: mux_26744 = 8'h0; 1: mux_26744 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26745;
  wire [7:0] v_26746;
  wire [7:0] v_26747;
  function [7:0] mux_26747(input [0:0] sel);
    case (sel) 0: mux_26747 = 8'h0; 1: mux_26747 = v_26748;
    endcase
  endfunction
  reg [7:0] v_26748 = 8'h0;
  wire [7:0] v_26749;
  wire [7:0] v_26750;
  function [7:0] mux_26750(input [0:0] sel);
    case (sel) 0: mux_26750 = 8'h0; 1: mux_26750 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26751;
  wire [7:0] v_26752;
  wire [7:0] v_26753;
  function [7:0] mux_26753(input [0:0] sel);
    case (sel) 0: mux_26753 = 8'h0; 1: mux_26753 = vout_peek_4012;
    endcase
  endfunction
  wire [7:0] v_26754;
  function [7:0] mux_26754(input [0:0] sel);
    case (sel) 0: mux_26754 = 8'h0; 1: mux_26754 = vout_peek_4003;
    endcase
  endfunction
  wire [7:0] v_26755;
  function [7:0] mux_26755(input [0:0] sel);
    case (sel) 0: mux_26755 = 8'h0; 1: mux_26755 = v_26756;
    endcase
  endfunction
  reg [7:0] v_26756 = 8'h0;
  wire [7:0] v_26757;
  wire [7:0] v_26758;
  function [7:0] mux_26758(input [0:0] sel);
    case (sel) 0: mux_26758 = 8'h0; 1: mux_26758 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26759;
  wire [7:0] v_26760;
  wire [7:0] v_26761;
  function [7:0] mux_26761(input [0:0] sel);
    case (sel) 0: mux_26761 = 8'h0; 1: mux_26761 = vout_peek_3975;
    endcase
  endfunction
  wire [7:0] v_26762;
  function [7:0] mux_26762(input [0:0] sel);
    case (sel) 0: mux_26762 = 8'h0; 1: mux_26762 = vout_peek_3966;
    endcase
  endfunction
  wire [7:0] v_26763;
  function [7:0] mux_26763(input [0:0] sel);
    case (sel) 0: mux_26763 = 8'h0; 1: mux_26763 = v_26764;
    endcase
  endfunction
  reg [7:0] v_26764 = 8'h0;
  wire [7:0] v_26765;
  wire [7:0] v_26766;
  function [7:0] mux_26766(input [0:0] sel);
    case (sel) 0: mux_26766 = 8'h0; 1: mux_26766 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26767;
  wire [7:0] v_26768;
  wire [7:0] v_26769;
  function [7:0] mux_26769(input [0:0] sel);
    case (sel) 0: mux_26769 = 8'h0; 1: mux_26769 = v_26770;
    endcase
  endfunction
  reg [7:0] v_26770 = 8'h0;
  wire [7:0] v_26771;
  wire [7:0] v_26772;
  function [7:0] mux_26772(input [0:0] sel);
    case (sel) 0: mux_26772 = 8'h0; 1: mux_26772 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26773;
  wire [7:0] v_26774;
  wire [7:0] v_26775;
  function [7:0] mux_26775(input [0:0] sel);
    case (sel) 0: mux_26775 = 8'h0; 1: mux_26775 = v_26776;
    endcase
  endfunction
  reg [7:0] v_26776 = 8'h0;
  wire [7:0] v_26777;
  wire [7:0] v_26778;
  function [7:0] mux_26778(input [0:0] sel);
    case (sel) 0: mux_26778 = 8'h0; 1: mux_26778 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26779;
  wire [7:0] v_26780;
  wire [7:0] v_26781;
  function [7:0] mux_26781(input [0:0] sel);
    case (sel) 0: mux_26781 = 8'h0; 1: mux_26781 = v_26782;
    endcase
  endfunction
  reg [7:0] v_26782 = 8'h0;
  wire [7:0] v_26783;
  wire [7:0] v_26784;
  function [7:0] mux_26784(input [0:0] sel);
    case (sel) 0: mux_26784 = 8'h0; 1: mux_26784 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26785;
  wire [7:0] v_26786;
  wire [7:0] v_26787;
  function [7:0] mux_26787(input [0:0] sel);
    case (sel) 0: mux_26787 = 8'h0; 1: mux_26787 = vout_peek_3881;
    endcase
  endfunction
  wire [7:0] v_26788;
  function [7:0] mux_26788(input [0:0] sel);
    case (sel) 0: mux_26788 = 8'h0; 1: mux_26788 = vout_peek_3872;
    endcase
  endfunction
  wire [7:0] v_26789;
  function [7:0] mux_26789(input [0:0] sel);
    case (sel) 0: mux_26789 = 8'h0; 1: mux_26789 = v_26790;
    endcase
  endfunction
  reg [7:0] v_26790 = 8'h0;
  wire [7:0] v_26791;
  wire [7:0] v_26792;
  function [7:0] mux_26792(input [0:0] sel);
    case (sel) 0: mux_26792 = 8'h0; 1: mux_26792 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26793;
  wire [7:0] v_26794;
  wire [7:0] v_26795;
  function [7:0] mux_26795(input [0:0] sel);
    case (sel) 0: mux_26795 = 8'h0; 1: mux_26795 = vout_peek_3844;
    endcase
  endfunction
  wire [7:0] v_26796;
  function [7:0] mux_26796(input [0:0] sel);
    case (sel) 0: mux_26796 = 8'h0; 1: mux_26796 = vout_peek_3835;
    endcase
  endfunction
  wire [7:0] v_26797;
  function [7:0] mux_26797(input [0:0] sel);
    case (sel) 0: mux_26797 = 8'h0; 1: mux_26797 = v_26798;
    endcase
  endfunction
  reg [7:0] v_26798 = 8'h0;
  wire [7:0] v_26799;
  wire [7:0] v_26800;
  function [7:0] mux_26800(input [0:0] sel);
    case (sel) 0: mux_26800 = 8'h0; 1: mux_26800 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26801;
  wire [7:0] v_26802;
  wire [7:0] v_26803;
  function [7:0] mux_26803(input [0:0] sel);
    case (sel) 0: mux_26803 = 8'h0; 1: mux_26803 = v_26804;
    endcase
  endfunction
  reg [7:0] v_26804 = 8'h0;
  wire [7:0] v_26805;
  wire [7:0] v_26806;
  function [7:0] mux_26806(input [0:0] sel);
    case (sel) 0: mux_26806 = 8'h0; 1: mux_26806 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26807;
  wire [7:0] v_26808;
  wire [7:0] v_26809;
  function [7:0] mux_26809(input [0:0] sel);
    case (sel) 0: mux_26809 = 8'h0; 1: mux_26809 = vout_peek_3788;
    endcase
  endfunction
  wire [7:0] v_26810;
  function [7:0] mux_26810(input [0:0] sel);
    case (sel) 0: mux_26810 = 8'h0; 1: mux_26810 = vout_peek_3779;
    endcase
  endfunction
  wire [7:0] v_26811;
  function [7:0] mux_26811(input [0:0] sel);
    case (sel) 0: mux_26811 = 8'h0; 1: mux_26811 = v_26812;
    endcase
  endfunction
  reg [7:0] v_26812 = 8'h0;
  wire [7:0] v_26813;
  wire [7:0] v_26814;
  function [7:0] mux_26814(input [0:0] sel);
    case (sel) 0: mux_26814 = 8'h0; 1: mux_26814 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26815;
  wire [7:0] v_26816;
  wire [7:0] v_26817;
  function [7:0] mux_26817(input [0:0] sel);
    case (sel) 0: mux_26817 = 8'h0; 1: mux_26817 = vout_peek_3751;
    endcase
  endfunction
  wire [7:0] v_26818;
  function [7:0] mux_26818(input [0:0] sel);
    case (sel) 0: mux_26818 = 8'h0; 1: mux_26818 = vout_peek_3742;
    endcase
  endfunction
  wire [7:0] v_26819;
  function [7:0] mux_26819(input [0:0] sel);
    case (sel) 0: mux_26819 = 8'h0; 1: mux_26819 = v_26820;
    endcase
  endfunction
  reg [7:0] v_26820 = 8'h0;
  wire [7:0] v_26821;
  wire [7:0] v_26822;
  function [7:0] mux_26822(input [0:0] sel);
    case (sel) 0: mux_26822 = 8'h0; 1: mux_26822 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26823;
  wire [7:0] v_26824;
  wire [7:0] v_26825;
  function [7:0] mux_26825(input [0:0] sel);
    case (sel) 0: mux_26825 = 8'h0; 1: mux_26825 = v_26826;
    endcase
  endfunction
  reg [7:0] v_26826 = 8'h0;
  wire [7:0] v_26827;
  wire [7:0] v_26828;
  function [7:0] mux_26828(input [0:0] sel);
    case (sel) 0: mux_26828 = 8'h0; 1: mux_26828 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26829;
  wire [7:0] v_26830;
  wire [7:0] v_26831;
  function [7:0] mux_26831(input [0:0] sel);
    case (sel) 0: mux_26831 = 8'h0; 1: mux_26831 = v_26832;
    endcase
  endfunction
  reg [7:0] v_26832 = 8'h0;
  wire [7:0] v_26833;
  wire [7:0] v_26834;
  function [7:0] mux_26834(input [0:0] sel);
    case (sel) 0: mux_26834 = 8'h0; 1: mux_26834 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26835;
  wire [7:0] v_26836;
  wire [7:0] v_26837;
  function [7:0] mux_26837(input [0:0] sel);
    case (sel) 0: mux_26837 = 8'h0; 1: mux_26837 = vout_peek_3676;
    endcase
  endfunction
  wire [7:0] v_26838;
  function [7:0] mux_26838(input [0:0] sel);
    case (sel) 0: mux_26838 = 8'h0; 1: mux_26838 = vout_peek_3667;
    endcase
  endfunction
  wire [7:0] v_26839;
  function [7:0] mux_26839(input [0:0] sel);
    case (sel) 0: mux_26839 = 8'h0; 1: mux_26839 = v_26840;
    endcase
  endfunction
  reg [7:0] v_26840 = 8'h0;
  wire [7:0] v_26841;
  wire [7:0] v_26842;
  function [7:0] mux_26842(input [0:0] sel);
    case (sel) 0: mux_26842 = 8'h0; 1: mux_26842 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26843;
  wire [7:0] v_26844;
  wire [7:0] v_26845;
  function [7:0] mux_26845(input [0:0] sel);
    case (sel) 0: mux_26845 = 8'h0; 1: mux_26845 = vout_peek_3639;
    endcase
  endfunction
  wire [7:0] v_26846;
  function [7:0] mux_26846(input [0:0] sel);
    case (sel) 0: mux_26846 = 8'h0; 1: mux_26846 = vout_peek_3630;
    endcase
  endfunction
  wire [7:0] v_26847;
  function [7:0] mux_26847(input [0:0] sel);
    case (sel) 0: mux_26847 = 8'h0; 1: mux_26847 = v_26848;
    endcase
  endfunction
  reg [7:0] v_26848 = 8'h0;
  wire [7:0] v_26849;
  wire [7:0] v_26850;
  function [7:0] mux_26850(input [0:0] sel);
    case (sel) 0: mux_26850 = 8'h0; 1: mux_26850 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26851;
  wire [7:0] v_26852;
  wire [7:0] v_26853;
  function [7:0] mux_26853(input [0:0] sel);
    case (sel) 0: mux_26853 = 8'h0; 1: mux_26853 = v_26854;
    endcase
  endfunction
  reg [7:0] v_26854 = 8'h0;
  wire [7:0] v_26855;
  wire [7:0] v_26856;
  function [7:0] mux_26856(input [0:0] sel);
    case (sel) 0: mux_26856 = 8'h0; 1: mux_26856 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26857;
  wire [7:0] v_26858;
  wire [7:0] v_26859;
  function [7:0] mux_26859(input [0:0] sel);
    case (sel) 0: mux_26859 = 8'h0; 1: mux_26859 = vout_peek_3583;
    endcase
  endfunction
  wire [7:0] v_26860;
  function [7:0] mux_26860(input [0:0] sel);
    case (sel) 0: mux_26860 = 8'h0; 1: mux_26860 = vout_peek_3574;
    endcase
  endfunction
  wire [7:0] v_26861;
  function [7:0] mux_26861(input [0:0] sel);
    case (sel) 0: mux_26861 = 8'h0; 1: mux_26861 = v_26862;
    endcase
  endfunction
  reg [7:0] v_26862 = 8'h0;
  wire [7:0] v_26863;
  wire [7:0] v_26864;
  function [7:0] mux_26864(input [0:0] sel);
    case (sel) 0: mux_26864 = 8'h0; 1: mux_26864 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26865;
  wire [7:0] v_26866;
  wire [7:0] v_26867;
  function [7:0] mux_26867(input [0:0] sel);
    case (sel) 0: mux_26867 = 8'h0; 1: mux_26867 = vout_peek_3546;
    endcase
  endfunction
  wire [7:0] v_26868;
  function [7:0] mux_26868(input [0:0] sel);
    case (sel) 0: mux_26868 = 8'h0; 1: mux_26868 = vout_peek_3537;
    endcase
  endfunction
  wire [7:0] v_26869;
  function [7:0] mux_26869(input [0:0] sel);
    case (sel) 0: mux_26869 = 8'h0; 1: mux_26869 = v_26870;
    endcase
  endfunction
  reg [7:0] v_26870 = 8'h0;
  wire [7:0] v_26871;
  wire [7:0] v_26872;
  function [7:0] mux_26872(input [0:0] sel);
    case (sel) 0: mux_26872 = 8'h0; 1: mux_26872 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26873;
  wire [7:0] v_26874;
  wire [7:0] v_26875;
  function [7:0] mux_26875(input [0:0] sel);
    case (sel) 0: mux_26875 = 8'h0; 1: mux_26875 = v_26876;
    endcase
  endfunction
  reg [7:0] v_26876 = 8'h0;
  wire [7:0] v_26877;
  wire [7:0] v_26878;
  function [7:0] mux_26878(input [0:0] sel);
    case (sel) 0: mux_26878 = 8'h0; 1: mux_26878 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26879;
  wire [7:0] v_26880;
  wire [7:0] v_26881;
  function [7:0] mux_26881(input [0:0] sel);
    case (sel) 0: mux_26881 = 8'h0; 1: mux_26881 = v_26882;
    endcase
  endfunction
  reg [7:0] v_26882 = 8'h0;
  wire [7:0] v_26883;
  wire [7:0] v_26884;
  function [7:0] mux_26884(input [0:0] sel);
    case (sel) 0: mux_26884 = 8'h0; 1: mux_26884 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26885;
  wire [7:0] v_26886;
  wire [7:0] v_26887;
  function [7:0] mux_26887(input [0:0] sel);
    case (sel) 0: mux_26887 = 8'h0; 1: mux_26887 = v_26888;
    endcase
  endfunction
  reg [7:0] v_26888 = 8'h0;
  wire [7:0] v_26889;
  wire [7:0] v_26890;
  function [7:0] mux_26890(input [0:0] sel);
    case (sel) 0: mux_26890 = 8'h0; 1: mux_26890 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26891;
  wire [7:0] v_26892;
  wire [7:0] v_26893;
  function [7:0] mux_26893(input [0:0] sel);
    case (sel) 0: mux_26893 = 8'h0; 1: mux_26893 = v_26894;
    endcase
  endfunction
  reg [7:0] v_26894 = 8'h0;
  wire [7:0] v_26895;
  wire [7:0] v_26896;
  function [7:0] mux_26896(input [0:0] sel);
    case (sel) 0: mux_26896 = 8'h0; 1: mux_26896 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26897;
  wire [7:0] v_26898;
  wire [7:0] v_26899;
  function [7:0] mux_26899(input [0:0] sel);
    case (sel) 0: mux_26899 = 8'h0; 1: mux_26899 = vout_peek_3433;
    endcase
  endfunction
  wire [7:0] v_26900;
  function [7:0] mux_26900(input [0:0] sel);
    case (sel) 0: mux_26900 = 8'h0; 1: mux_26900 = vout_peek_3424;
    endcase
  endfunction
  wire [7:0] v_26901;
  function [7:0] mux_26901(input [0:0] sel);
    case (sel) 0: mux_26901 = 8'h0; 1: mux_26901 = v_26902;
    endcase
  endfunction
  reg [7:0] v_26902 = 8'h0;
  wire [7:0] v_26903;
  wire [7:0] v_26904;
  function [7:0] mux_26904(input [0:0] sel);
    case (sel) 0: mux_26904 = 8'h0; 1: mux_26904 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26905;
  wire [7:0] v_26906;
  wire [7:0] v_26907;
  function [7:0] mux_26907(input [0:0] sel);
    case (sel) 0: mux_26907 = 8'h0; 1: mux_26907 = vout_peek_3396;
    endcase
  endfunction
  wire [7:0] v_26908;
  function [7:0] mux_26908(input [0:0] sel);
    case (sel) 0: mux_26908 = 8'h0; 1: mux_26908 = vout_peek_3387;
    endcase
  endfunction
  wire [7:0] v_26909;
  function [7:0] mux_26909(input [0:0] sel);
    case (sel) 0: mux_26909 = 8'h0; 1: mux_26909 = v_26910;
    endcase
  endfunction
  reg [7:0] v_26910 = 8'h0;
  wire [7:0] v_26911;
  wire [7:0] v_26912;
  function [7:0] mux_26912(input [0:0] sel);
    case (sel) 0: mux_26912 = 8'h0; 1: mux_26912 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26913;
  wire [7:0] v_26914;
  wire [7:0] v_26915;
  function [7:0] mux_26915(input [0:0] sel);
    case (sel) 0: mux_26915 = 8'h0; 1: mux_26915 = v_26916;
    endcase
  endfunction
  reg [7:0] v_26916 = 8'h0;
  wire [7:0] v_26917;
  wire [7:0] v_26918;
  function [7:0] mux_26918(input [0:0] sel);
    case (sel) 0: mux_26918 = 8'h0; 1: mux_26918 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26919;
  wire [7:0] v_26920;
  wire [7:0] v_26921;
  function [7:0] mux_26921(input [0:0] sel);
    case (sel) 0: mux_26921 = 8'h0; 1: mux_26921 = vout_peek_3340;
    endcase
  endfunction
  wire [7:0] v_26922;
  function [7:0] mux_26922(input [0:0] sel);
    case (sel) 0: mux_26922 = 8'h0; 1: mux_26922 = vout_peek_3331;
    endcase
  endfunction
  wire [7:0] v_26923;
  function [7:0] mux_26923(input [0:0] sel);
    case (sel) 0: mux_26923 = 8'h0; 1: mux_26923 = v_26924;
    endcase
  endfunction
  reg [7:0] v_26924 = 8'h0;
  wire [7:0] v_26925;
  wire [7:0] v_26926;
  function [7:0] mux_26926(input [0:0] sel);
    case (sel) 0: mux_26926 = 8'h0; 1: mux_26926 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26927;
  wire [7:0] v_26928;
  wire [7:0] v_26929;
  function [7:0] mux_26929(input [0:0] sel);
    case (sel) 0: mux_26929 = 8'h0; 1: mux_26929 = vout_peek_3303;
    endcase
  endfunction
  wire [7:0] v_26930;
  function [7:0] mux_26930(input [0:0] sel);
    case (sel) 0: mux_26930 = 8'h0; 1: mux_26930 = vout_peek_3294;
    endcase
  endfunction
  wire [7:0] v_26931;
  function [7:0] mux_26931(input [0:0] sel);
    case (sel) 0: mux_26931 = 8'h0; 1: mux_26931 = v_26932;
    endcase
  endfunction
  reg [7:0] v_26932 = 8'h0;
  wire [7:0] v_26933;
  wire [7:0] v_26934;
  function [7:0] mux_26934(input [0:0] sel);
    case (sel) 0: mux_26934 = 8'h0; 1: mux_26934 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26935;
  wire [7:0] v_26936;
  wire [7:0] v_26937;
  function [7:0] mux_26937(input [0:0] sel);
    case (sel) 0: mux_26937 = 8'h0; 1: mux_26937 = v_26938;
    endcase
  endfunction
  reg [7:0] v_26938 = 8'h0;
  wire [7:0] v_26939;
  wire [7:0] v_26940;
  function [7:0] mux_26940(input [0:0] sel);
    case (sel) 0: mux_26940 = 8'h0; 1: mux_26940 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26941;
  wire [7:0] v_26942;
  wire [7:0] v_26943;
  function [7:0] mux_26943(input [0:0] sel);
    case (sel) 0: mux_26943 = 8'h0; 1: mux_26943 = v_26944;
    endcase
  endfunction
  reg [7:0] v_26944 = 8'h0;
  wire [7:0] v_26945;
  wire [7:0] v_26946;
  function [7:0] mux_26946(input [0:0] sel);
    case (sel) 0: mux_26946 = 8'h0; 1: mux_26946 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26947;
  wire [7:0] v_26948;
  wire [7:0] v_26949;
  function [7:0] mux_26949(input [0:0] sel);
    case (sel) 0: mux_26949 = 8'h0; 1: mux_26949 = vout_peek_3228;
    endcase
  endfunction
  wire [7:0] v_26950;
  function [7:0] mux_26950(input [0:0] sel);
    case (sel) 0: mux_26950 = 8'h0; 1: mux_26950 = vout_peek_3219;
    endcase
  endfunction
  wire [7:0] v_26951;
  function [7:0] mux_26951(input [0:0] sel);
    case (sel) 0: mux_26951 = 8'h0; 1: mux_26951 = v_26952;
    endcase
  endfunction
  reg [7:0] v_26952 = 8'h0;
  wire [7:0] v_26953;
  wire [7:0] v_26954;
  function [7:0] mux_26954(input [0:0] sel);
    case (sel) 0: mux_26954 = 8'h0; 1: mux_26954 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26955;
  wire [7:0] v_26956;
  wire [7:0] v_26957;
  function [7:0] mux_26957(input [0:0] sel);
    case (sel) 0: mux_26957 = 8'h0; 1: mux_26957 = vout_peek_3191;
    endcase
  endfunction
  wire [7:0] v_26958;
  function [7:0] mux_26958(input [0:0] sel);
    case (sel) 0: mux_26958 = 8'h0; 1: mux_26958 = vout_peek_3182;
    endcase
  endfunction
  wire [7:0] v_26959;
  function [7:0] mux_26959(input [0:0] sel);
    case (sel) 0: mux_26959 = 8'h0; 1: mux_26959 = v_26960;
    endcase
  endfunction
  reg [7:0] v_26960 = 8'h0;
  wire [7:0] v_26961;
  wire [7:0] v_26962;
  function [7:0] mux_26962(input [0:0] sel);
    case (sel) 0: mux_26962 = 8'h0; 1: mux_26962 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26963;
  wire [7:0] v_26964;
  wire [7:0] v_26965;
  function [7:0] mux_26965(input [0:0] sel);
    case (sel) 0: mux_26965 = 8'h0; 1: mux_26965 = v_26966;
    endcase
  endfunction
  reg [7:0] v_26966 = 8'h0;
  wire [7:0] v_26967;
  wire [7:0] v_26968;
  function [7:0] mux_26968(input [0:0] sel);
    case (sel) 0: mux_26968 = 8'h0; 1: mux_26968 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26969;
  wire [7:0] v_26970;
  wire [7:0] v_26971;
  function [7:0] mux_26971(input [0:0] sel);
    case (sel) 0: mux_26971 = 8'h0; 1: mux_26971 = vout_peek_3135;
    endcase
  endfunction
  wire [7:0] v_26972;
  function [7:0] mux_26972(input [0:0] sel);
    case (sel) 0: mux_26972 = 8'h0; 1: mux_26972 = vout_peek_3126;
    endcase
  endfunction
  wire [7:0] v_26973;
  function [7:0] mux_26973(input [0:0] sel);
    case (sel) 0: mux_26973 = 8'h0; 1: mux_26973 = v_26974;
    endcase
  endfunction
  reg [7:0] v_26974 = 8'h0;
  wire [7:0] v_26975;
  wire [7:0] v_26976;
  function [7:0] mux_26976(input [0:0] sel);
    case (sel) 0: mux_26976 = 8'h0; 1: mux_26976 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26977;
  wire [7:0] v_26978;
  wire [7:0] v_26979;
  function [7:0] mux_26979(input [0:0] sel);
    case (sel) 0: mux_26979 = 8'h0; 1: mux_26979 = vout_peek_3098;
    endcase
  endfunction
  wire [7:0] v_26980;
  function [7:0] mux_26980(input [0:0] sel);
    case (sel) 0: mux_26980 = 8'h0; 1: mux_26980 = vout_peek_3089;
    endcase
  endfunction
  wire [7:0] v_26981;
  function [7:0] mux_26981(input [0:0] sel);
    case (sel) 0: mux_26981 = 8'h0; 1: mux_26981 = v_26982;
    endcase
  endfunction
  reg [7:0] v_26982 = 8'h0;
  wire [7:0] v_26983;
  wire [7:0] v_26984;
  function [7:0] mux_26984(input [0:0] sel);
    case (sel) 0: mux_26984 = 8'h0; 1: mux_26984 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26985;
  wire [7:0] v_26986;
  wire [7:0] v_26987;
  function [7:0] mux_26987(input [0:0] sel);
    case (sel) 0: mux_26987 = 8'h0; 1: mux_26987 = v_26988;
    endcase
  endfunction
  reg [7:0] v_26988 = 8'h0;
  wire [7:0] v_26989;
  wire [7:0] v_26990;
  function [7:0] mux_26990(input [0:0] sel);
    case (sel) 0: mux_26990 = 8'h0; 1: mux_26990 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26991;
  wire [7:0] v_26992;
  wire [7:0] v_26993;
  function [7:0] mux_26993(input [0:0] sel);
    case (sel) 0: mux_26993 = 8'h0; 1: mux_26993 = v_26994;
    endcase
  endfunction
  reg [7:0] v_26994 = 8'h0;
  wire [7:0] v_26995;
  wire [7:0] v_26996;
  function [7:0] mux_26996(input [0:0] sel);
    case (sel) 0: mux_26996 = 8'h0; 1: mux_26996 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_26997;
  wire [7:0] v_26998;
  wire [7:0] v_26999;
  function [7:0] mux_26999(input [0:0] sel);
    case (sel) 0: mux_26999 = 8'h0; 1: mux_26999 = v_27000;
    endcase
  endfunction
  reg [7:0] v_27000 = 8'h0;
  wire [7:0] v_27001;
  wire [7:0] v_27002;
  function [7:0] mux_27002(input [0:0] sel);
    case (sel) 0: mux_27002 = 8'h0; 1: mux_27002 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27003;
  wire [7:0] v_27004;
  wire [7:0] v_27005;
  function [7:0] mux_27005(input [0:0] sel);
    case (sel) 0: mux_27005 = 8'h0; 1: mux_27005 = vout_peek_3004;
    endcase
  endfunction
  wire [7:0] v_27006;
  function [7:0] mux_27006(input [0:0] sel);
    case (sel) 0: mux_27006 = 8'h0; 1: mux_27006 = vout_peek_2995;
    endcase
  endfunction
  wire [7:0] v_27007;
  function [7:0] mux_27007(input [0:0] sel);
    case (sel) 0: mux_27007 = 8'h0; 1: mux_27007 = v_27008;
    endcase
  endfunction
  reg [7:0] v_27008 = 8'h0;
  wire [7:0] v_27009;
  wire [7:0] v_27010;
  function [7:0] mux_27010(input [0:0] sel);
    case (sel) 0: mux_27010 = 8'h0; 1: mux_27010 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27011;
  wire [7:0] v_27012;
  wire [7:0] v_27013;
  function [7:0] mux_27013(input [0:0] sel);
    case (sel) 0: mux_27013 = 8'h0; 1: mux_27013 = vout_peek_2967;
    endcase
  endfunction
  wire [7:0] v_27014;
  function [7:0] mux_27014(input [0:0] sel);
    case (sel) 0: mux_27014 = 8'h0; 1: mux_27014 = vout_peek_2958;
    endcase
  endfunction
  wire [7:0] v_27015;
  function [7:0] mux_27015(input [0:0] sel);
    case (sel) 0: mux_27015 = 8'h0; 1: mux_27015 = v_27016;
    endcase
  endfunction
  reg [7:0] v_27016 = 8'h0;
  wire [7:0] v_27017;
  wire [7:0] v_27018;
  function [7:0] mux_27018(input [0:0] sel);
    case (sel) 0: mux_27018 = 8'h0; 1: mux_27018 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27019;
  wire [7:0] v_27020;
  wire [7:0] v_27021;
  function [7:0] mux_27021(input [0:0] sel);
    case (sel) 0: mux_27021 = 8'h0; 1: mux_27021 = v_27022;
    endcase
  endfunction
  reg [7:0] v_27022 = 8'h0;
  wire [7:0] v_27023;
  wire [7:0] v_27024;
  function [7:0] mux_27024(input [0:0] sel);
    case (sel) 0: mux_27024 = 8'h0; 1: mux_27024 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27025;
  wire [7:0] v_27026;
  wire [7:0] v_27027;
  function [7:0] mux_27027(input [0:0] sel);
    case (sel) 0: mux_27027 = 8'h0; 1: mux_27027 = vout_peek_2911;
    endcase
  endfunction
  wire [7:0] v_27028;
  function [7:0] mux_27028(input [0:0] sel);
    case (sel) 0: mux_27028 = 8'h0; 1: mux_27028 = vout_peek_2902;
    endcase
  endfunction
  wire [7:0] v_27029;
  function [7:0] mux_27029(input [0:0] sel);
    case (sel) 0: mux_27029 = 8'h0; 1: mux_27029 = v_27030;
    endcase
  endfunction
  reg [7:0] v_27030 = 8'h0;
  wire [7:0] v_27031;
  wire [7:0] v_27032;
  function [7:0] mux_27032(input [0:0] sel);
    case (sel) 0: mux_27032 = 8'h0; 1: mux_27032 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27033;
  wire [7:0] v_27034;
  wire [7:0] v_27035;
  function [7:0] mux_27035(input [0:0] sel);
    case (sel) 0: mux_27035 = 8'h0; 1: mux_27035 = vout_peek_2874;
    endcase
  endfunction
  wire [7:0] v_27036;
  function [7:0] mux_27036(input [0:0] sel);
    case (sel) 0: mux_27036 = 8'h0; 1: mux_27036 = vout_peek_2865;
    endcase
  endfunction
  wire [7:0] v_27037;
  function [7:0] mux_27037(input [0:0] sel);
    case (sel) 0: mux_27037 = 8'h0; 1: mux_27037 = v_27038;
    endcase
  endfunction
  reg [7:0] v_27038 = 8'h0;
  wire [7:0] v_27039;
  wire [7:0] v_27040;
  function [7:0] mux_27040(input [0:0] sel);
    case (sel) 0: mux_27040 = 8'h0; 1: mux_27040 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27041;
  wire [7:0] v_27042;
  wire [7:0] v_27043;
  function [7:0] mux_27043(input [0:0] sel);
    case (sel) 0: mux_27043 = 8'h0; 1: mux_27043 = v_27044;
    endcase
  endfunction
  reg [7:0] v_27044 = 8'h0;
  wire [7:0] v_27045;
  wire [7:0] v_27046;
  function [7:0] mux_27046(input [0:0] sel);
    case (sel) 0: mux_27046 = 8'h0; 1: mux_27046 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27047;
  wire [7:0] v_27048;
  wire [7:0] v_27049;
  function [7:0] mux_27049(input [0:0] sel);
    case (sel) 0: mux_27049 = 8'h0; 1: mux_27049 = v_27050;
    endcase
  endfunction
  reg [7:0] v_27050 = 8'h0;
  wire [7:0] v_27051;
  wire [7:0] v_27052;
  function [7:0] mux_27052(input [0:0] sel);
    case (sel) 0: mux_27052 = 8'h0; 1: mux_27052 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27053;
  wire [7:0] v_27054;
  wire [7:0] v_27055;
  function [7:0] mux_27055(input [0:0] sel);
    case (sel) 0: mux_27055 = 8'h0; 1: mux_27055 = vout_peek_2799;
    endcase
  endfunction
  wire [7:0] v_27056;
  function [7:0] mux_27056(input [0:0] sel);
    case (sel) 0: mux_27056 = 8'h0; 1: mux_27056 = vout_peek_2790;
    endcase
  endfunction
  wire [7:0] v_27057;
  function [7:0] mux_27057(input [0:0] sel);
    case (sel) 0: mux_27057 = 8'h0; 1: mux_27057 = v_27058;
    endcase
  endfunction
  reg [7:0] v_27058 = 8'h0;
  wire [7:0] v_27059;
  wire [7:0] v_27060;
  function [7:0] mux_27060(input [0:0] sel);
    case (sel) 0: mux_27060 = 8'h0; 1: mux_27060 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27061;
  wire [7:0] v_27062;
  wire [7:0] v_27063;
  function [7:0] mux_27063(input [0:0] sel);
    case (sel) 0: mux_27063 = 8'h0; 1: mux_27063 = vout_peek_2762;
    endcase
  endfunction
  wire [7:0] v_27064;
  function [7:0] mux_27064(input [0:0] sel);
    case (sel) 0: mux_27064 = 8'h0; 1: mux_27064 = vout_peek_2753;
    endcase
  endfunction
  wire [7:0] v_27065;
  function [7:0] mux_27065(input [0:0] sel);
    case (sel) 0: mux_27065 = 8'h0; 1: mux_27065 = v_27066;
    endcase
  endfunction
  reg [7:0] v_27066 = 8'h0;
  wire [7:0] v_27067;
  wire [7:0] v_27068;
  function [7:0] mux_27068(input [0:0] sel);
    case (sel) 0: mux_27068 = 8'h0; 1: mux_27068 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27069;
  wire [7:0] v_27070;
  wire [7:0] v_27071;
  function [7:0] mux_27071(input [0:0] sel);
    case (sel) 0: mux_27071 = 8'h0; 1: mux_27071 = v_27072;
    endcase
  endfunction
  reg [7:0] v_27072 = 8'h0;
  wire [7:0] v_27073;
  wire [7:0] v_27074;
  function [7:0] mux_27074(input [0:0] sel);
    case (sel) 0: mux_27074 = 8'h0; 1: mux_27074 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27075;
  wire [7:0] v_27076;
  wire [7:0] v_27077;
  function [7:0] mux_27077(input [0:0] sel);
    case (sel) 0: mux_27077 = 8'h0; 1: mux_27077 = vout_peek_2706;
    endcase
  endfunction
  wire [7:0] v_27078;
  function [7:0] mux_27078(input [0:0] sel);
    case (sel) 0: mux_27078 = 8'h0; 1: mux_27078 = vout_peek_2697;
    endcase
  endfunction
  wire [7:0] v_27079;
  function [7:0] mux_27079(input [0:0] sel);
    case (sel) 0: mux_27079 = 8'h0; 1: mux_27079 = v_27080;
    endcase
  endfunction
  reg [7:0] v_27080 = 8'h0;
  wire [7:0] v_27081;
  wire [7:0] v_27082;
  function [7:0] mux_27082(input [0:0] sel);
    case (sel) 0: mux_27082 = 8'h0; 1: mux_27082 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27083;
  wire [7:0] v_27084;
  wire [7:0] v_27085;
  function [7:0] mux_27085(input [0:0] sel);
    case (sel) 0: mux_27085 = 8'h0; 1: mux_27085 = vout_peek_2669;
    endcase
  endfunction
  wire [7:0] v_27086;
  function [7:0] mux_27086(input [0:0] sel);
    case (sel) 0: mux_27086 = 8'h0; 1: mux_27086 = vout_peek_2660;
    endcase
  endfunction
  wire [7:0] v_27087;
  function [7:0] mux_27087(input [0:0] sel);
    case (sel) 0: mux_27087 = 8'h0; 1: mux_27087 = v_27088;
    endcase
  endfunction
  reg [7:0] v_27088 = 8'h0;
  wire [7:0] v_27089;
  wire [7:0] v_27090;
  function [7:0] mux_27090(input [0:0] sel);
    case (sel) 0: mux_27090 = 8'h0; 1: mux_27090 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27091;
  wire [7:0] v_27092;
  wire [7:0] v_27093;
  function [7:0] mux_27093(input [0:0] sel);
    case (sel) 0: mux_27093 = 8'h0; 1: mux_27093 = v_27094;
    endcase
  endfunction
  reg [7:0] v_27094 = 8'h0;
  wire [7:0] v_27095;
  wire [7:0] v_27096;
  function [7:0] mux_27096(input [0:0] sel);
    case (sel) 0: mux_27096 = 8'h0; 1: mux_27096 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27097;
  wire [7:0] v_27098;
  wire [7:0] v_27099;
  function [7:0] mux_27099(input [0:0] sel);
    case (sel) 0: mux_27099 = 8'h0; 1: mux_27099 = v_27100;
    endcase
  endfunction
  reg [7:0] v_27100 = 8'h0;
  wire [7:0] v_27101;
  wire [7:0] v_27102;
  function [7:0] mux_27102(input [0:0] sel);
    case (sel) 0: mux_27102 = 8'h0; 1: mux_27102 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27103;
  wire [7:0] v_27104;
  wire [7:0] v_27105;
  function [7:0] mux_27105(input [0:0] sel);
    case (sel) 0: mux_27105 = 8'h0; 1: mux_27105 = v_27106;
    endcase
  endfunction
  reg [7:0] v_27106 = 8'h0;
  wire [7:0] v_27107;
  wire [7:0] v_27108;
  function [7:0] mux_27108(input [0:0] sel);
    case (sel) 0: mux_27108 = 8'h0; 1: mux_27108 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27109;
  wire [7:0] v_27110;
  wire [7:0] v_27111;
  function [7:0] mux_27111(input [0:0] sel);
    case (sel) 0: mux_27111 = 8'h0; 1: mux_27111 = v_27112;
    endcase
  endfunction
  reg [7:0] v_27112 = 8'h0;
  wire [7:0] v_27113;
  wire [7:0] v_27114;
  function [7:0] mux_27114(input [0:0] sel);
    case (sel) 0: mux_27114 = 8'h0; 1: mux_27114 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27115;
  wire [7:0] v_27116;
  wire [7:0] v_27117;
  function [7:0] mux_27117(input [0:0] sel);
    case (sel) 0: mux_27117 = 8'h0; 1: mux_27117 = v_27118;
    endcase
  endfunction
  reg [7:0] v_27118 = 8'h0;
  wire [7:0] v_27119;
  wire [7:0] v_27120;
  function [7:0] mux_27120(input [0:0] sel);
    case (sel) 0: mux_27120 = 8'h0; 1: mux_27120 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27121;
  wire [7:0] v_27122;
  wire [7:0] v_27123;
  function [7:0] mux_27123(input [0:0] sel);
    case (sel) 0: mux_27123 = 8'h0; 1: mux_27123 = v_27124;
    endcase
  endfunction
  reg [7:0] v_27124 = 8'h0;
  wire [7:0] v_27125;
  wire [7:0] v_27126;
  function [7:0] mux_27126(input [0:0] sel);
    case (sel) 0: mux_27126 = 8'h0; 1: mux_27126 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27127;
  wire [7:0] v_27128;
  wire [7:0] v_27129;
  function [7:0] mux_27129(input [0:0] sel);
    case (sel) 0: mux_27129 = 8'h0; 1: mux_27129 = vout_peek_7870;
    endcase
  endfunction
  wire [7:0] v_27130;
  function [7:0] mux_27130(input [0:0] sel);
    case (sel) 0: mux_27130 = 8'h0; 1: mux_27130 = vout_peek_7861;
    endcase
  endfunction
  wire [7:0] v_27131;
  function [7:0] mux_27131(input [0:0] sel);
    case (sel) 0: mux_27131 = 8'h0; 1: mux_27131 = v_27132;
    endcase
  endfunction
  reg [7:0] v_27132 = 8'h0;
  wire [7:0] v_27133;
  wire [7:0] v_27134;
  function [7:0] mux_27134(input [0:0] sel);
    case (sel) 0: mux_27134 = 8'h0; 1: mux_27134 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27135;
  wire [7:0] v_27136;
  wire [7:0] v_27137;
  function [7:0] mux_27137(input [0:0] sel);
    case (sel) 0: mux_27137 = 8'h0; 1: mux_27137 = vout_peek_7833;
    endcase
  endfunction
  wire [7:0] v_27138;
  function [7:0] mux_27138(input [0:0] sel);
    case (sel) 0: mux_27138 = 8'h0; 1: mux_27138 = vout_peek_7824;
    endcase
  endfunction
  wire [7:0] v_27139;
  function [7:0] mux_27139(input [0:0] sel);
    case (sel) 0: mux_27139 = 8'h0; 1: mux_27139 = v_27140;
    endcase
  endfunction
  reg [7:0] v_27140 = 8'h0;
  wire [7:0] v_27141;
  wire [7:0] v_27142;
  function [7:0] mux_27142(input [0:0] sel);
    case (sel) 0: mux_27142 = 8'h0; 1: mux_27142 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27143;
  wire [7:0] v_27144;
  wire [7:0] v_27145;
  function [7:0] mux_27145(input [0:0] sel);
    case (sel) 0: mux_27145 = 8'h0; 1: mux_27145 = v_27146;
    endcase
  endfunction
  reg [7:0] v_27146 = 8'h0;
  wire [7:0] v_27147;
  wire [7:0] v_27148;
  function [7:0] mux_27148(input [0:0] sel);
    case (sel) 0: mux_27148 = 8'h0; 1: mux_27148 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27149;
  wire [7:0] v_27150;
  wire [7:0] v_27151;
  function [7:0] mux_27151(input [0:0] sel);
    case (sel) 0: mux_27151 = 8'h0; 1: mux_27151 = vout_peek_7777;
    endcase
  endfunction
  wire [7:0] v_27152;
  function [7:0] mux_27152(input [0:0] sel);
    case (sel) 0: mux_27152 = 8'h0; 1: mux_27152 = vout_peek_7768;
    endcase
  endfunction
  wire [7:0] v_27153;
  function [7:0] mux_27153(input [0:0] sel);
    case (sel) 0: mux_27153 = 8'h0; 1: mux_27153 = v_27154;
    endcase
  endfunction
  reg [7:0] v_27154 = 8'h0;
  wire [7:0] v_27155;
  wire [7:0] v_27156;
  function [7:0] mux_27156(input [0:0] sel);
    case (sel) 0: mux_27156 = 8'h0; 1: mux_27156 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27157;
  wire [7:0] v_27158;
  wire [7:0] v_27159;
  function [7:0] mux_27159(input [0:0] sel);
    case (sel) 0: mux_27159 = 8'h0; 1: mux_27159 = vout_peek_7740;
    endcase
  endfunction
  wire [7:0] v_27160;
  function [7:0] mux_27160(input [0:0] sel);
    case (sel) 0: mux_27160 = 8'h0; 1: mux_27160 = vout_peek_7731;
    endcase
  endfunction
  wire [7:0] v_27161;
  function [7:0] mux_27161(input [0:0] sel);
    case (sel) 0: mux_27161 = 8'h0; 1: mux_27161 = v_27162;
    endcase
  endfunction
  reg [7:0] v_27162 = 8'h0;
  wire [7:0] v_27163;
  wire [7:0] v_27164;
  function [7:0] mux_27164(input [0:0] sel);
    case (sel) 0: mux_27164 = 8'h0; 1: mux_27164 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27165;
  wire [7:0] v_27166;
  wire [7:0] v_27167;
  function [7:0] mux_27167(input [0:0] sel);
    case (sel) 0: mux_27167 = 8'h0; 1: mux_27167 = v_27168;
    endcase
  endfunction
  reg [7:0] v_27168 = 8'h0;
  wire [7:0] v_27169;
  wire [7:0] v_27170;
  function [7:0] mux_27170(input [0:0] sel);
    case (sel) 0: mux_27170 = 8'h0; 1: mux_27170 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27171;
  wire [7:0] v_27172;
  wire [7:0] v_27173;
  function [7:0] mux_27173(input [0:0] sel);
    case (sel) 0: mux_27173 = 8'h0; 1: mux_27173 = v_27174;
    endcase
  endfunction
  reg [7:0] v_27174 = 8'h0;
  wire [7:0] v_27175;
  wire [7:0] v_27176;
  function [7:0] mux_27176(input [0:0] sel);
    case (sel) 0: mux_27176 = 8'h0; 1: mux_27176 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27177;
  wire [7:0] v_27178;
  wire [7:0] v_27179;
  function [7:0] mux_27179(input [0:0] sel);
    case (sel) 0: mux_27179 = 8'h0; 1: mux_27179 = vout_peek_7665;
    endcase
  endfunction
  wire [7:0] v_27180;
  function [7:0] mux_27180(input [0:0] sel);
    case (sel) 0: mux_27180 = 8'h0; 1: mux_27180 = vout_peek_7656;
    endcase
  endfunction
  wire [7:0] v_27181;
  function [7:0] mux_27181(input [0:0] sel);
    case (sel) 0: mux_27181 = 8'h0; 1: mux_27181 = v_27182;
    endcase
  endfunction
  reg [7:0] v_27182 = 8'h0;
  wire [7:0] v_27183;
  wire [7:0] v_27184;
  function [7:0] mux_27184(input [0:0] sel);
    case (sel) 0: mux_27184 = 8'h0; 1: mux_27184 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27185;
  wire [7:0] v_27186;
  wire [7:0] v_27187;
  function [7:0] mux_27187(input [0:0] sel);
    case (sel) 0: mux_27187 = 8'h0; 1: mux_27187 = vout_peek_7628;
    endcase
  endfunction
  wire [7:0] v_27188;
  function [7:0] mux_27188(input [0:0] sel);
    case (sel) 0: mux_27188 = 8'h0; 1: mux_27188 = vout_peek_7619;
    endcase
  endfunction
  wire [7:0] v_27189;
  function [7:0] mux_27189(input [0:0] sel);
    case (sel) 0: mux_27189 = 8'h0; 1: mux_27189 = v_27190;
    endcase
  endfunction
  reg [7:0] v_27190 = 8'h0;
  wire [7:0] v_27191;
  wire [7:0] v_27192;
  function [7:0] mux_27192(input [0:0] sel);
    case (sel) 0: mux_27192 = 8'h0; 1: mux_27192 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27193;
  wire [7:0] v_27194;
  wire [7:0] v_27195;
  function [7:0] mux_27195(input [0:0] sel);
    case (sel) 0: mux_27195 = 8'h0; 1: mux_27195 = v_27196;
    endcase
  endfunction
  reg [7:0] v_27196 = 8'h0;
  wire [7:0] v_27197;
  wire [7:0] v_27198;
  function [7:0] mux_27198(input [0:0] sel);
    case (sel) 0: mux_27198 = 8'h0; 1: mux_27198 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27199;
  wire [7:0] v_27200;
  wire [7:0] v_27201;
  function [7:0] mux_27201(input [0:0] sel);
    case (sel) 0: mux_27201 = 8'h0; 1: mux_27201 = vout_peek_7572;
    endcase
  endfunction
  wire [7:0] v_27202;
  function [7:0] mux_27202(input [0:0] sel);
    case (sel) 0: mux_27202 = 8'h0; 1: mux_27202 = vout_peek_7563;
    endcase
  endfunction
  wire [7:0] v_27203;
  function [7:0] mux_27203(input [0:0] sel);
    case (sel) 0: mux_27203 = 8'h0; 1: mux_27203 = v_27204;
    endcase
  endfunction
  reg [7:0] v_27204 = 8'h0;
  wire [7:0] v_27205;
  wire [7:0] v_27206;
  function [7:0] mux_27206(input [0:0] sel);
    case (sel) 0: mux_27206 = 8'h0; 1: mux_27206 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27207;
  wire [7:0] v_27208;
  wire [7:0] v_27209;
  function [7:0] mux_27209(input [0:0] sel);
    case (sel) 0: mux_27209 = 8'h0; 1: mux_27209 = vout_peek_7535;
    endcase
  endfunction
  wire [7:0] v_27210;
  function [7:0] mux_27210(input [0:0] sel);
    case (sel) 0: mux_27210 = 8'h0; 1: mux_27210 = vout_peek_7526;
    endcase
  endfunction
  wire [7:0] v_27211;
  function [7:0] mux_27211(input [0:0] sel);
    case (sel) 0: mux_27211 = 8'h0; 1: mux_27211 = v_27212;
    endcase
  endfunction
  reg [7:0] v_27212 = 8'h0;
  wire [7:0] v_27213;
  wire [7:0] v_27214;
  function [7:0] mux_27214(input [0:0] sel);
    case (sel) 0: mux_27214 = 8'h0; 1: mux_27214 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27215;
  wire [7:0] v_27216;
  wire [7:0] v_27217;
  function [7:0] mux_27217(input [0:0] sel);
    case (sel) 0: mux_27217 = 8'h0; 1: mux_27217 = v_27218;
    endcase
  endfunction
  reg [7:0] v_27218 = 8'h0;
  wire [7:0] v_27219;
  wire [7:0] v_27220;
  function [7:0] mux_27220(input [0:0] sel);
    case (sel) 0: mux_27220 = 8'h0; 1: mux_27220 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27221;
  wire [7:0] v_27222;
  wire [7:0] v_27223;
  function [7:0] mux_27223(input [0:0] sel);
    case (sel) 0: mux_27223 = 8'h0; 1: mux_27223 = v_27224;
    endcase
  endfunction
  reg [7:0] v_27224 = 8'h0;
  wire [7:0] v_27225;
  wire [7:0] v_27226;
  function [7:0] mux_27226(input [0:0] sel);
    case (sel) 0: mux_27226 = 8'h0; 1: mux_27226 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27227;
  wire [7:0] v_27228;
  wire [7:0] v_27229;
  function [7:0] mux_27229(input [0:0] sel);
    case (sel) 0: mux_27229 = 8'h0; 1: mux_27229 = v_27230;
    endcase
  endfunction
  reg [7:0] v_27230 = 8'h0;
  wire [7:0] v_27231;
  wire [7:0] v_27232;
  function [7:0] mux_27232(input [0:0] sel);
    case (sel) 0: mux_27232 = 8'h0; 1: mux_27232 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27233;
  wire [7:0] v_27234;
  wire [7:0] v_27235;
  function [7:0] mux_27235(input [0:0] sel);
    case (sel) 0: mux_27235 = 8'h0; 1: mux_27235 = vout_peek_7441;
    endcase
  endfunction
  wire [7:0] v_27236;
  function [7:0] mux_27236(input [0:0] sel);
    case (sel) 0: mux_27236 = 8'h0; 1: mux_27236 = vout_peek_7432;
    endcase
  endfunction
  wire [7:0] v_27237;
  function [7:0] mux_27237(input [0:0] sel);
    case (sel) 0: mux_27237 = 8'h0; 1: mux_27237 = v_27238;
    endcase
  endfunction
  reg [7:0] v_27238 = 8'h0;
  wire [7:0] v_27239;
  wire [7:0] v_27240;
  function [7:0] mux_27240(input [0:0] sel);
    case (sel) 0: mux_27240 = 8'h0; 1: mux_27240 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27241;
  wire [7:0] v_27242;
  wire [7:0] v_27243;
  function [7:0] mux_27243(input [0:0] sel);
    case (sel) 0: mux_27243 = 8'h0; 1: mux_27243 = vout_peek_7404;
    endcase
  endfunction
  wire [7:0] v_27244;
  function [7:0] mux_27244(input [0:0] sel);
    case (sel) 0: mux_27244 = 8'h0; 1: mux_27244 = vout_peek_7395;
    endcase
  endfunction
  wire [7:0] v_27245;
  function [7:0] mux_27245(input [0:0] sel);
    case (sel) 0: mux_27245 = 8'h0; 1: mux_27245 = v_27246;
    endcase
  endfunction
  reg [7:0] v_27246 = 8'h0;
  wire [7:0] v_27247;
  wire [7:0] v_27248;
  function [7:0] mux_27248(input [0:0] sel);
    case (sel) 0: mux_27248 = 8'h0; 1: mux_27248 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27249;
  wire [7:0] v_27250;
  wire [7:0] v_27251;
  function [7:0] mux_27251(input [0:0] sel);
    case (sel) 0: mux_27251 = 8'h0; 1: mux_27251 = v_27252;
    endcase
  endfunction
  reg [7:0] v_27252 = 8'h0;
  wire [7:0] v_27253;
  wire [7:0] v_27254;
  function [7:0] mux_27254(input [0:0] sel);
    case (sel) 0: mux_27254 = 8'h0; 1: mux_27254 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27255;
  wire [7:0] v_27256;
  wire [7:0] v_27257;
  function [7:0] mux_27257(input [0:0] sel);
    case (sel) 0: mux_27257 = 8'h0; 1: mux_27257 = vout_peek_7348;
    endcase
  endfunction
  wire [7:0] v_27258;
  function [7:0] mux_27258(input [0:0] sel);
    case (sel) 0: mux_27258 = 8'h0; 1: mux_27258 = vout_peek_7339;
    endcase
  endfunction
  wire [7:0] v_27259;
  function [7:0] mux_27259(input [0:0] sel);
    case (sel) 0: mux_27259 = 8'h0; 1: mux_27259 = v_27260;
    endcase
  endfunction
  reg [7:0] v_27260 = 8'h0;
  wire [7:0] v_27261;
  wire [7:0] v_27262;
  function [7:0] mux_27262(input [0:0] sel);
    case (sel) 0: mux_27262 = 8'h0; 1: mux_27262 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27263;
  wire [7:0] v_27264;
  wire [7:0] v_27265;
  function [7:0] mux_27265(input [0:0] sel);
    case (sel) 0: mux_27265 = 8'h0; 1: mux_27265 = vout_peek_7311;
    endcase
  endfunction
  wire [7:0] v_27266;
  function [7:0] mux_27266(input [0:0] sel);
    case (sel) 0: mux_27266 = 8'h0; 1: mux_27266 = vout_peek_7302;
    endcase
  endfunction
  wire [7:0] v_27267;
  function [7:0] mux_27267(input [0:0] sel);
    case (sel) 0: mux_27267 = 8'h0; 1: mux_27267 = v_27268;
    endcase
  endfunction
  reg [7:0] v_27268 = 8'h0;
  wire [7:0] v_27269;
  wire [7:0] v_27270;
  function [7:0] mux_27270(input [0:0] sel);
    case (sel) 0: mux_27270 = 8'h0; 1: mux_27270 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27271;
  wire [7:0] v_27272;
  wire [7:0] v_27273;
  function [7:0] mux_27273(input [0:0] sel);
    case (sel) 0: mux_27273 = 8'h0; 1: mux_27273 = v_27274;
    endcase
  endfunction
  reg [7:0] v_27274 = 8'h0;
  wire [7:0] v_27275;
  wire [7:0] v_27276;
  function [7:0] mux_27276(input [0:0] sel);
    case (sel) 0: mux_27276 = 8'h0; 1: mux_27276 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27277;
  wire [7:0] v_27278;
  wire [7:0] v_27279;
  function [7:0] mux_27279(input [0:0] sel);
    case (sel) 0: mux_27279 = 8'h0; 1: mux_27279 = v_27280;
    endcase
  endfunction
  reg [7:0] v_27280 = 8'h0;
  wire [7:0] v_27281;
  wire [7:0] v_27282;
  function [7:0] mux_27282(input [0:0] sel);
    case (sel) 0: mux_27282 = 8'h0; 1: mux_27282 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27283;
  wire [7:0] v_27284;
  wire [7:0] v_27285;
  function [7:0] mux_27285(input [0:0] sel);
    case (sel) 0: mux_27285 = 8'h0; 1: mux_27285 = vout_peek_7236;
    endcase
  endfunction
  wire [7:0] v_27286;
  function [7:0] mux_27286(input [0:0] sel);
    case (sel) 0: mux_27286 = 8'h0; 1: mux_27286 = vout_peek_7227;
    endcase
  endfunction
  wire [7:0] v_27287;
  function [7:0] mux_27287(input [0:0] sel);
    case (sel) 0: mux_27287 = 8'h0; 1: mux_27287 = v_27288;
    endcase
  endfunction
  reg [7:0] v_27288 = 8'h0;
  wire [7:0] v_27289;
  wire [7:0] v_27290;
  function [7:0] mux_27290(input [0:0] sel);
    case (sel) 0: mux_27290 = 8'h0; 1: mux_27290 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27291;
  wire [7:0] v_27292;
  wire [7:0] v_27293;
  function [7:0] mux_27293(input [0:0] sel);
    case (sel) 0: mux_27293 = 8'h0; 1: mux_27293 = vout_peek_7199;
    endcase
  endfunction
  wire [7:0] v_27294;
  function [7:0] mux_27294(input [0:0] sel);
    case (sel) 0: mux_27294 = 8'h0; 1: mux_27294 = vout_peek_7190;
    endcase
  endfunction
  wire [7:0] v_27295;
  function [7:0] mux_27295(input [0:0] sel);
    case (sel) 0: mux_27295 = 8'h0; 1: mux_27295 = v_27296;
    endcase
  endfunction
  reg [7:0] v_27296 = 8'h0;
  wire [7:0] v_27297;
  wire [7:0] v_27298;
  function [7:0] mux_27298(input [0:0] sel);
    case (sel) 0: mux_27298 = 8'h0; 1: mux_27298 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27299;
  wire [7:0] v_27300;
  wire [7:0] v_27301;
  function [7:0] mux_27301(input [0:0] sel);
    case (sel) 0: mux_27301 = 8'h0; 1: mux_27301 = v_27302;
    endcase
  endfunction
  reg [7:0] v_27302 = 8'h0;
  wire [7:0] v_27303;
  wire [7:0] v_27304;
  function [7:0] mux_27304(input [0:0] sel);
    case (sel) 0: mux_27304 = 8'h0; 1: mux_27304 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27305;
  wire [7:0] v_27306;
  wire [7:0] v_27307;
  function [7:0] mux_27307(input [0:0] sel);
    case (sel) 0: mux_27307 = 8'h0; 1: mux_27307 = vout_peek_7143;
    endcase
  endfunction
  wire [7:0] v_27308;
  function [7:0] mux_27308(input [0:0] sel);
    case (sel) 0: mux_27308 = 8'h0; 1: mux_27308 = vout_peek_7134;
    endcase
  endfunction
  wire [7:0] v_27309;
  function [7:0] mux_27309(input [0:0] sel);
    case (sel) 0: mux_27309 = 8'h0; 1: mux_27309 = v_27310;
    endcase
  endfunction
  reg [7:0] v_27310 = 8'h0;
  wire [7:0] v_27311;
  wire [7:0] v_27312;
  function [7:0] mux_27312(input [0:0] sel);
    case (sel) 0: mux_27312 = 8'h0; 1: mux_27312 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27313;
  wire [7:0] v_27314;
  wire [7:0] v_27315;
  function [7:0] mux_27315(input [0:0] sel);
    case (sel) 0: mux_27315 = 8'h0; 1: mux_27315 = vout_peek_7106;
    endcase
  endfunction
  wire [7:0] v_27316;
  function [7:0] mux_27316(input [0:0] sel);
    case (sel) 0: mux_27316 = 8'h0; 1: mux_27316 = vout_peek_7097;
    endcase
  endfunction
  wire [7:0] v_27317;
  function [7:0] mux_27317(input [0:0] sel);
    case (sel) 0: mux_27317 = 8'h0; 1: mux_27317 = v_27318;
    endcase
  endfunction
  reg [7:0] v_27318 = 8'h0;
  wire [7:0] v_27319;
  wire [7:0] v_27320;
  function [7:0] mux_27320(input [0:0] sel);
    case (sel) 0: mux_27320 = 8'h0; 1: mux_27320 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27321;
  wire [7:0] v_27322;
  wire [7:0] v_27323;
  function [7:0] mux_27323(input [0:0] sel);
    case (sel) 0: mux_27323 = 8'h0; 1: mux_27323 = v_27324;
    endcase
  endfunction
  reg [7:0] v_27324 = 8'h0;
  wire [7:0] v_27325;
  wire [7:0] v_27326;
  function [7:0] mux_27326(input [0:0] sel);
    case (sel) 0: mux_27326 = 8'h0; 1: mux_27326 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27327;
  wire [7:0] v_27328;
  wire [7:0] v_27329;
  function [7:0] mux_27329(input [0:0] sel);
    case (sel) 0: mux_27329 = 8'h0; 1: mux_27329 = v_27330;
    endcase
  endfunction
  reg [7:0] v_27330 = 8'h0;
  wire [7:0] v_27331;
  wire [7:0] v_27332;
  function [7:0] mux_27332(input [0:0] sel);
    case (sel) 0: mux_27332 = 8'h0; 1: mux_27332 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27333;
  wire [7:0] v_27334;
  wire [7:0] v_27335;
  function [7:0] mux_27335(input [0:0] sel);
    case (sel) 0: mux_27335 = 8'h0; 1: mux_27335 = v_27336;
    endcase
  endfunction
  reg [7:0] v_27336 = 8'h0;
  wire [7:0] v_27337;
  wire [7:0] v_27338;
  function [7:0] mux_27338(input [0:0] sel);
    case (sel) 0: mux_27338 = 8'h0; 1: mux_27338 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27339;
  wire [7:0] v_27340;
  wire [7:0] v_27341;
  function [7:0] mux_27341(input [0:0] sel);
    case (sel) 0: mux_27341 = 8'h0; 1: mux_27341 = v_27342;
    endcase
  endfunction
  reg [7:0] v_27342 = 8'h0;
  wire [7:0] v_27343;
  wire [7:0] v_27344;
  function [7:0] mux_27344(input [0:0] sel);
    case (sel) 0: mux_27344 = 8'h0; 1: mux_27344 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27345;
  wire [7:0] v_27346;
  wire [7:0] v_27347;
  function [7:0] mux_27347(input [0:0] sel);
    case (sel) 0: mux_27347 = 8'h0; 1: mux_27347 = vout_peek_6993;
    endcase
  endfunction
  wire [7:0] v_27348;
  function [7:0] mux_27348(input [0:0] sel);
    case (sel) 0: mux_27348 = 8'h0; 1: mux_27348 = vout_peek_6984;
    endcase
  endfunction
  wire [7:0] v_27349;
  function [7:0] mux_27349(input [0:0] sel);
    case (sel) 0: mux_27349 = 8'h0; 1: mux_27349 = v_27350;
    endcase
  endfunction
  reg [7:0] v_27350 = 8'h0;
  wire [7:0] v_27351;
  wire [7:0] v_27352;
  function [7:0] mux_27352(input [0:0] sel);
    case (sel) 0: mux_27352 = 8'h0; 1: mux_27352 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27353;
  wire [7:0] v_27354;
  wire [7:0] v_27355;
  function [7:0] mux_27355(input [0:0] sel);
    case (sel) 0: mux_27355 = 8'h0; 1: mux_27355 = vout_peek_6956;
    endcase
  endfunction
  wire [7:0] v_27356;
  function [7:0] mux_27356(input [0:0] sel);
    case (sel) 0: mux_27356 = 8'h0; 1: mux_27356 = vout_peek_6947;
    endcase
  endfunction
  wire [7:0] v_27357;
  function [7:0] mux_27357(input [0:0] sel);
    case (sel) 0: mux_27357 = 8'h0; 1: mux_27357 = v_27358;
    endcase
  endfunction
  reg [7:0] v_27358 = 8'h0;
  wire [7:0] v_27359;
  wire [7:0] v_27360;
  function [7:0] mux_27360(input [0:0] sel);
    case (sel) 0: mux_27360 = 8'h0; 1: mux_27360 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27361;
  wire [7:0] v_27362;
  wire [7:0] v_27363;
  function [7:0] mux_27363(input [0:0] sel);
    case (sel) 0: mux_27363 = 8'h0; 1: mux_27363 = v_27364;
    endcase
  endfunction
  reg [7:0] v_27364 = 8'h0;
  wire [7:0] v_27365;
  wire [7:0] v_27366;
  function [7:0] mux_27366(input [0:0] sel);
    case (sel) 0: mux_27366 = 8'h0; 1: mux_27366 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27367;
  wire [7:0] v_27368;
  wire [7:0] v_27369;
  function [7:0] mux_27369(input [0:0] sel);
    case (sel) 0: mux_27369 = 8'h0; 1: mux_27369 = vout_peek_6900;
    endcase
  endfunction
  wire [7:0] v_27370;
  function [7:0] mux_27370(input [0:0] sel);
    case (sel) 0: mux_27370 = 8'h0; 1: mux_27370 = vout_peek_6891;
    endcase
  endfunction
  wire [7:0] v_27371;
  function [7:0] mux_27371(input [0:0] sel);
    case (sel) 0: mux_27371 = 8'h0; 1: mux_27371 = v_27372;
    endcase
  endfunction
  reg [7:0] v_27372 = 8'h0;
  wire [7:0] v_27373;
  wire [7:0] v_27374;
  function [7:0] mux_27374(input [0:0] sel);
    case (sel) 0: mux_27374 = 8'h0; 1: mux_27374 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27375;
  wire [7:0] v_27376;
  wire [7:0] v_27377;
  function [7:0] mux_27377(input [0:0] sel);
    case (sel) 0: mux_27377 = 8'h0; 1: mux_27377 = vout_peek_6863;
    endcase
  endfunction
  wire [7:0] v_27378;
  function [7:0] mux_27378(input [0:0] sel);
    case (sel) 0: mux_27378 = 8'h0; 1: mux_27378 = vout_peek_6854;
    endcase
  endfunction
  wire [7:0] v_27379;
  function [7:0] mux_27379(input [0:0] sel);
    case (sel) 0: mux_27379 = 8'h0; 1: mux_27379 = v_27380;
    endcase
  endfunction
  reg [7:0] v_27380 = 8'h0;
  wire [7:0] v_27381;
  wire [7:0] v_27382;
  function [7:0] mux_27382(input [0:0] sel);
    case (sel) 0: mux_27382 = 8'h0; 1: mux_27382 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27383;
  wire [7:0] v_27384;
  wire [7:0] v_27385;
  function [7:0] mux_27385(input [0:0] sel);
    case (sel) 0: mux_27385 = 8'h0; 1: mux_27385 = v_27386;
    endcase
  endfunction
  reg [7:0] v_27386 = 8'h0;
  wire [7:0] v_27387;
  wire [7:0] v_27388;
  function [7:0] mux_27388(input [0:0] sel);
    case (sel) 0: mux_27388 = 8'h0; 1: mux_27388 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27389;
  wire [7:0] v_27390;
  wire [7:0] v_27391;
  function [7:0] mux_27391(input [0:0] sel);
    case (sel) 0: mux_27391 = 8'h0; 1: mux_27391 = v_27392;
    endcase
  endfunction
  reg [7:0] v_27392 = 8'h0;
  wire [7:0] v_27393;
  wire [7:0] v_27394;
  function [7:0] mux_27394(input [0:0] sel);
    case (sel) 0: mux_27394 = 8'h0; 1: mux_27394 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27395;
  wire [7:0] v_27396;
  wire [7:0] v_27397;
  function [7:0] mux_27397(input [0:0] sel);
    case (sel) 0: mux_27397 = 8'h0; 1: mux_27397 = vout_peek_6788;
    endcase
  endfunction
  wire [7:0] v_27398;
  function [7:0] mux_27398(input [0:0] sel);
    case (sel) 0: mux_27398 = 8'h0; 1: mux_27398 = vout_peek_6779;
    endcase
  endfunction
  wire [7:0] v_27399;
  function [7:0] mux_27399(input [0:0] sel);
    case (sel) 0: mux_27399 = 8'h0; 1: mux_27399 = v_27400;
    endcase
  endfunction
  reg [7:0] v_27400 = 8'h0;
  wire [7:0] v_27401;
  wire [7:0] v_27402;
  function [7:0] mux_27402(input [0:0] sel);
    case (sel) 0: mux_27402 = 8'h0; 1: mux_27402 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27403;
  wire [7:0] v_27404;
  wire [7:0] v_27405;
  function [7:0] mux_27405(input [0:0] sel);
    case (sel) 0: mux_27405 = 8'h0; 1: mux_27405 = vout_peek_6751;
    endcase
  endfunction
  wire [7:0] v_27406;
  function [7:0] mux_27406(input [0:0] sel);
    case (sel) 0: mux_27406 = 8'h0; 1: mux_27406 = vout_peek_6742;
    endcase
  endfunction
  wire [7:0] v_27407;
  function [7:0] mux_27407(input [0:0] sel);
    case (sel) 0: mux_27407 = 8'h0; 1: mux_27407 = v_27408;
    endcase
  endfunction
  reg [7:0] v_27408 = 8'h0;
  wire [7:0] v_27409;
  wire [7:0] v_27410;
  function [7:0] mux_27410(input [0:0] sel);
    case (sel) 0: mux_27410 = 8'h0; 1: mux_27410 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27411;
  wire [7:0] v_27412;
  wire [7:0] v_27413;
  function [7:0] mux_27413(input [0:0] sel);
    case (sel) 0: mux_27413 = 8'h0; 1: mux_27413 = v_27414;
    endcase
  endfunction
  reg [7:0] v_27414 = 8'h0;
  wire [7:0] v_27415;
  wire [7:0] v_27416;
  function [7:0] mux_27416(input [0:0] sel);
    case (sel) 0: mux_27416 = 8'h0; 1: mux_27416 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27417;
  wire [7:0] v_27418;
  wire [7:0] v_27419;
  function [7:0] mux_27419(input [0:0] sel);
    case (sel) 0: mux_27419 = 8'h0; 1: mux_27419 = vout_peek_6695;
    endcase
  endfunction
  wire [7:0] v_27420;
  function [7:0] mux_27420(input [0:0] sel);
    case (sel) 0: mux_27420 = 8'h0; 1: mux_27420 = vout_peek_6686;
    endcase
  endfunction
  wire [7:0] v_27421;
  function [7:0] mux_27421(input [0:0] sel);
    case (sel) 0: mux_27421 = 8'h0; 1: mux_27421 = v_27422;
    endcase
  endfunction
  reg [7:0] v_27422 = 8'h0;
  wire [7:0] v_27423;
  wire [7:0] v_27424;
  function [7:0] mux_27424(input [0:0] sel);
    case (sel) 0: mux_27424 = 8'h0; 1: mux_27424 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27425;
  wire [7:0] v_27426;
  wire [7:0] v_27427;
  function [7:0] mux_27427(input [0:0] sel);
    case (sel) 0: mux_27427 = 8'h0; 1: mux_27427 = vout_peek_6658;
    endcase
  endfunction
  wire [7:0] v_27428;
  function [7:0] mux_27428(input [0:0] sel);
    case (sel) 0: mux_27428 = 8'h0; 1: mux_27428 = vout_peek_6649;
    endcase
  endfunction
  wire [7:0] v_27429;
  function [7:0] mux_27429(input [0:0] sel);
    case (sel) 0: mux_27429 = 8'h0; 1: mux_27429 = v_27430;
    endcase
  endfunction
  reg [7:0] v_27430 = 8'h0;
  wire [7:0] v_27431;
  wire [7:0] v_27432;
  function [7:0] mux_27432(input [0:0] sel);
    case (sel) 0: mux_27432 = 8'h0; 1: mux_27432 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27433;
  wire [7:0] v_27434;
  wire [7:0] v_27435;
  function [7:0] mux_27435(input [0:0] sel);
    case (sel) 0: mux_27435 = 8'h0; 1: mux_27435 = v_27436;
    endcase
  endfunction
  reg [7:0] v_27436 = 8'h0;
  wire [7:0] v_27437;
  wire [7:0] v_27438;
  function [7:0] mux_27438(input [0:0] sel);
    case (sel) 0: mux_27438 = 8'h0; 1: mux_27438 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27439;
  wire [7:0] v_27440;
  wire [7:0] v_27441;
  function [7:0] mux_27441(input [0:0] sel);
    case (sel) 0: mux_27441 = 8'h0; 1: mux_27441 = v_27442;
    endcase
  endfunction
  reg [7:0] v_27442 = 8'h0;
  wire [7:0] v_27443;
  wire [7:0] v_27444;
  function [7:0] mux_27444(input [0:0] sel);
    case (sel) 0: mux_27444 = 8'h0; 1: mux_27444 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27445;
  wire [7:0] v_27446;
  wire [7:0] v_27447;
  function [7:0] mux_27447(input [0:0] sel);
    case (sel) 0: mux_27447 = 8'h0; 1: mux_27447 = v_27448;
    endcase
  endfunction
  reg [7:0] v_27448 = 8'h0;
  wire [7:0] v_27449;
  wire [7:0] v_27450;
  function [7:0] mux_27450(input [0:0] sel);
    case (sel) 0: mux_27450 = 8'h0; 1: mux_27450 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27451;
  wire [7:0] v_27452;
  wire [7:0] v_27453;
  function [7:0] mux_27453(input [0:0] sel);
    case (sel) 0: mux_27453 = 8'h0; 1: mux_27453 = vout_peek_6564;
    endcase
  endfunction
  wire [7:0] v_27454;
  function [7:0] mux_27454(input [0:0] sel);
    case (sel) 0: mux_27454 = 8'h0; 1: mux_27454 = vout_peek_6555;
    endcase
  endfunction
  wire [7:0] v_27455;
  function [7:0] mux_27455(input [0:0] sel);
    case (sel) 0: mux_27455 = 8'h0; 1: mux_27455 = v_27456;
    endcase
  endfunction
  reg [7:0] v_27456 = 8'h0;
  wire [7:0] v_27457;
  wire [7:0] v_27458;
  function [7:0] mux_27458(input [0:0] sel);
    case (sel) 0: mux_27458 = 8'h0; 1: mux_27458 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27459;
  wire [7:0] v_27460;
  wire [7:0] v_27461;
  function [7:0] mux_27461(input [0:0] sel);
    case (sel) 0: mux_27461 = 8'h0; 1: mux_27461 = vout_peek_6527;
    endcase
  endfunction
  wire [7:0] v_27462;
  function [7:0] mux_27462(input [0:0] sel);
    case (sel) 0: mux_27462 = 8'h0; 1: mux_27462 = vout_peek_6518;
    endcase
  endfunction
  wire [7:0] v_27463;
  function [7:0] mux_27463(input [0:0] sel);
    case (sel) 0: mux_27463 = 8'h0; 1: mux_27463 = v_27464;
    endcase
  endfunction
  reg [7:0] v_27464 = 8'h0;
  wire [7:0] v_27465;
  wire [7:0] v_27466;
  function [7:0] mux_27466(input [0:0] sel);
    case (sel) 0: mux_27466 = 8'h0; 1: mux_27466 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27467;
  wire [7:0] v_27468;
  wire [7:0] v_27469;
  function [7:0] mux_27469(input [0:0] sel);
    case (sel) 0: mux_27469 = 8'h0; 1: mux_27469 = v_27470;
    endcase
  endfunction
  reg [7:0] v_27470 = 8'h0;
  wire [7:0] v_27471;
  wire [7:0] v_27472;
  function [7:0] mux_27472(input [0:0] sel);
    case (sel) 0: mux_27472 = 8'h0; 1: mux_27472 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27473;
  wire [7:0] v_27474;
  wire [7:0] v_27475;
  function [7:0] mux_27475(input [0:0] sel);
    case (sel) 0: mux_27475 = 8'h0; 1: mux_27475 = vout_peek_6471;
    endcase
  endfunction
  wire [7:0] v_27476;
  function [7:0] mux_27476(input [0:0] sel);
    case (sel) 0: mux_27476 = 8'h0; 1: mux_27476 = vout_peek_6462;
    endcase
  endfunction
  wire [7:0] v_27477;
  function [7:0] mux_27477(input [0:0] sel);
    case (sel) 0: mux_27477 = 8'h0; 1: mux_27477 = v_27478;
    endcase
  endfunction
  reg [7:0] v_27478 = 8'h0;
  wire [7:0] v_27479;
  wire [7:0] v_27480;
  function [7:0] mux_27480(input [0:0] sel);
    case (sel) 0: mux_27480 = 8'h0; 1: mux_27480 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27481;
  wire [7:0] v_27482;
  wire [7:0] v_27483;
  function [7:0] mux_27483(input [0:0] sel);
    case (sel) 0: mux_27483 = 8'h0; 1: mux_27483 = vout_peek_6434;
    endcase
  endfunction
  wire [7:0] v_27484;
  function [7:0] mux_27484(input [0:0] sel);
    case (sel) 0: mux_27484 = 8'h0; 1: mux_27484 = vout_peek_6425;
    endcase
  endfunction
  wire [7:0] v_27485;
  function [7:0] mux_27485(input [0:0] sel);
    case (sel) 0: mux_27485 = 8'h0; 1: mux_27485 = v_27486;
    endcase
  endfunction
  reg [7:0] v_27486 = 8'h0;
  wire [7:0] v_27487;
  wire [7:0] v_27488;
  function [7:0] mux_27488(input [0:0] sel);
    case (sel) 0: mux_27488 = 8'h0; 1: mux_27488 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27489;
  wire [7:0] v_27490;
  wire [7:0] v_27491;
  function [7:0] mux_27491(input [0:0] sel);
    case (sel) 0: mux_27491 = 8'h0; 1: mux_27491 = v_27492;
    endcase
  endfunction
  reg [7:0] v_27492 = 8'h0;
  wire [7:0] v_27493;
  wire [7:0] v_27494;
  function [7:0] mux_27494(input [0:0] sel);
    case (sel) 0: mux_27494 = 8'h0; 1: mux_27494 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27495;
  wire [7:0] v_27496;
  wire [7:0] v_27497;
  function [7:0] mux_27497(input [0:0] sel);
    case (sel) 0: mux_27497 = 8'h0; 1: mux_27497 = v_27498;
    endcase
  endfunction
  reg [7:0] v_27498 = 8'h0;
  wire [7:0] v_27499;
  wire [7:0] v_27500;
  function [7:0] mux_27500(input [0:0] sel);
    case (sel) 0: mux_27500 = 8'h0; 1: mux_27500 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27501;
  wire [7:0] v_27502;
  wire [7:0] v_27503;
  function [7:0] mux_27503(input [0:0] sel);
    case (sel) 0: mux_27503 = 8'h0; 1: mux_27503 = vout_peek_6359;
    endcase
  endfunction
  wire [7:0] v_27504;
  function [7:0] mux_27504(input [0:0] sel);
    case (sel) 0: mux_27504 = 8'h0; 1: mux_27504 = vout_peek_6350;
    endcase
  endfunction
  wire [7:0] v_27505;
  function [7:0] mux_27505(input [0:0] sel);
    case (sel) 0: mux_27505 = 8'h0; 1: mux_27505 = v_27506;
    endcase
  endfunction
  reg [7:0] v_27506 = 8'h0;
  wire [7:0] v_27507;
  wire [7:0] v_27508;
  function [7:0] mux_27508(input [0:0] sel);
    case (sel) 0: mux_27508 = 8'h0; 1: mux_27508 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27509;
  wire [7:0] v_27510;
  wire [7:0] v_27511;
  function [7:0] mux_27511(input [0:0] sel);
    case (sel) 0: mux_27511 = 8'h0; 1: mux_27511 = vout_peek_6322;
    endcase
  endfunction
  wire [7:0] v_27512;
  function [7:0] mux_27512(input [0:0] sel);
    case (sel) 0: mux_27512 = 8'h0; 1: mux_27512 = vout_peek_6313;
    endcase
  endfunction
  wire [7:0] v_27513;
  function [7:0] mux_27513(input [0:0] sel);
    case (sel) 0: mux_27513 = 8'h0; 1: mux_27513 = v_27514;
    endcase
  endfunction
  reg [7:0] v_27514 = 8'h0;
  wire [7:0] v_27515;
  wire [7:0] v_27516;
  function [7:0] mux_27516(input [0:0] sel);
    case (sel) 0: mux_27516 = 8'h0; 1: mux_27516 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27517;
  wire [7:0] v_27518;
  wire [7:0] v_27519;
  function [7:0] mux_27519(input [0:0] sel);
    case (sel) 0: mux_27519 = 8'h0; 1: mux_27519 = v_27520;
    endcase
  endfunction
  reg [7:0] v_27520 = 8'h0;
  wire [7:0] v_27521;
  wire [7:0] v_27522;
  function [7:0] mux_27522(input [0:0] sel);
    case (sel) 0: mux_27522 = 8'h0; 1: mux_27522 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27523;
  wire [7:0] v_27524;
  wire [7:0] v_27525;
  function [7:0] mux_27525(input [0:0] sel);
    case (sel) 0: mux_27525 = 8'h0; 1: mux_27525 = vout_peek_6266;
    endcase
  endfunction
  wire [7:0] v_27526;
  function [7:0] mux_27526(input [0:0] sel);
    case (sel) 0: mux_27526 = 8'h0; 1: mux_27526 = vout_peek_6257;
    endcase
  endfunction
  wire [7:0] v_27527;
  function [7:0] mux_27527(input [0:0] sel);
    case (sel) 0: mux_27527 = 8'h0; 1: mux_27527 = v_27528;
    endcase
  endfunction
  reg [7:0] v_27528 = 8'h0;
  wire [7:0] v_27529;
  wire [7:0] v_27530;
  function [7:0] mux_27530(input [0:0] sel);
    case (sel) 0: mux_27530 = 8'h0; 1: mux_27530 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27531;
  wire [7:0] v_27532;
  wire [7:0] v_27533;
  function [7:0] mux_27533(input [0:0] sel);
    case (sel) 0: mux_27533 = 8'h0; 1: mux_27533 = vout_peek_6229;
    endcase
  endfunction
  wire [7:0] v_27534;
  function [7:0] mux_27534(input [0:0] sel);
    case (sel) 0: mux_27534 = 8'h0; 1: mux_27534 = vout_peek_6220;
    endcase
  endfunction
  wire [7:0] v_27535;
  function [7:0] mux_27535(input [0:0] sel);
    case (sel) 0: mux_27535 = 8'h0; 1: mux_27535 = v_27536;
    endcase
  endfunction
  reg [7:0] v_27536 = 8'h0;
  wire [7:0] v_27537;
  wire [7:0] v_27538;
  function [7:0] mux_27538(input [0:0] sel);
    case (sel) 0: mux_27538 = 8'h0; 1: mux_27538 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27539;
  wire [7:0] v_27540;
  wire [7:0] v_27541;
  function [7:0] mux_27541(input [0:0] sel);
    case (sel) 0: mux_27541 = 8'h0; 1: mux_27541 = v_27542;
    endcase
  endfunction
  reg [7:0] v_27542 = 8'h0;
  wire [7:0] v_27543;
  wire [7:0] v_27544;
  function [7:0] mux_27544(input [0:0] sel);
    case (sel) 0: mux_27544 = 8'h0; 1: mux_27544 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27545;
  wire [7:0] v_27546;
  wire [7:0] v_27547;
  function [7:0] mux_27547(input [0:0] sel);
    case (sel) 0: mux_27547 = 8'h0; 1: mux_27547 = v_27548;
    endcase
  endfunction
  reg [7:0] v_27548 = 8'h0;
  wire [7:0] v_27549;
  wire [7:0] v_27550;
  function [7:0] mux_27550(input [0:0] sel);
    case (sel) 0: mux_27550 = 8'h0; 1: mux_27550 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27551;
  wire [7:0] v_27552;
  wire [7:0] v_27553;
  function [7:0] mux_27553(input [0:0] sel);
    case (sel) 0: mux_27553 = 8'h0; 1: mux_27553 = v_27554;
    endcase
  endfunction
  reg [7:0] v_27554 = 8'h0;
  wire [7:0] v_27555;
  wire [7:0] v_27556;
  function [7:0] mux_27556(input [0:0] sel);
    case (sel) 0: mux_27556 = 8'h0; 1: mux_27556 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27557;
  wire [7:0] v_27558;
  wire [7:0] v_27559;
  function [7:0] mux_27559(input [0:0] sel);
    case (sel) 0: mux_27559 = 8'h0; 1: mux_27559 = v_27560;
    endcase
  endfunction
  reg [7:0] v_27560 = 8'h0;
  wire [7:0] v_27561;
  wire [7:0] v_27562;
  function [7:0] mux_27562(input [0:0] sel);
    case (sel) 0: mux_27562 = 8'h0; 1: mux_27562 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27563;
  wire [7:0] v_27564;
  wire [7:0] v_27565;
  function [7:0] mux_27565(input [0:0] sel);
    case (sel) 0: mux_27565 = 8'h0; 1: mux_27565 = v_27566;
    endcase
  endfunction
  reg [7:0] v_27566 = 8'h0;
  wire [7:0] v_27567;
  wire [7:0] v_27568;
  function [7:0] mux_27568(input [0:0] sel);
    case (sel) 0: mux_27568 = 8'h0; 1: mux_27568 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27569;
  wire [7:0] v_27570;
  wire [7:0] v_27571;
  function [7:0] mux_27571(input [0:0] sel);
    case (sel) 0: mux_27571 = 8'h0; 1: mux_27571 = vout_peek_6097;
    endcase
  endfunction
  wire [7:0] v_27572;
  function [7:0] mux_27572(input [0:0] sel);
    case (sel) 0: mux_27572 = 8'h0; 1: mux_27572 = vout_peek_6088;
    endcase
  endfunction
  wire [7:0] v_27573;
  function [7:0] mux_27573(input [0:0] sel);
    case (sel) 0: mux_27573 = 8'h0; 1: mux_27573 = v_27574;
    endcase
  endfunction
  reg [7:0] v_27574 = 8'h0;
  wire [7:0] v_27575;
  wire [7:0] v_27576;
  function [7:0] mux_27576(input [0:0] sel);
    case (sel) 0: mux_27576 = 8'h0; 1: mux_27576 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27577;
  wire [7:0] v_27578;
  wire [7:0] v_27579;
  function [7:0] mux_27579(input [0:0] sel);
    case (sel) 0: mux_27579 = 8'h0; 1: mux_27579 = vout_peek_6060;
    endcase
  endfunction
  wire [7:0] v_27580;
  function [7:0] mux_27580(input [0:0] sel);
    case (sel) 0: mux_27580 = 8'h0; 1: mux_27580 = vout_peek_6051;
    endcase
  endfunction
  wire [7:0] v_27581;
  function [7:0] mux_27581(input [0:0] sel);
    case (sel) 0: mux_27581 = 8'h0; 1: mux_27581 = v_27582;
    endcase
  endfunction
  reg [7:0] v_27582 = 8'h0;
  wire [7:0] v_27583;
  wire [7:0] v_27584;
  function [7:0] mux_27584(input [0:0] sel);
    case (sel) 0: mux_27584 = 8'h0; 1: mux_27584 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27585;
  wire [7:0] v_27586;
  wire [7:0] v_27587;
  function [7:0] mux_27587(input [0:0] sel);
    case (sel) 0: mux_27587 = 8'h0; 1: mux_27587 = v_27588;
    endcase
  endfunction
  reg [7:0] v_27588 = 8'h0;
  wire [7:0] v_27589;
  wire [7:0] v_27590;
  function [7:0] mux_27590(input [0:0] sel);
    case (sel) 0: mux_27590 = 8'h0; 1: mux_27590 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27591;
  wire [7:0] v_27592;
  wire [7:0] v_27593;
  function [7:0] mux_27593(input [0:0] sel);
    case (sel) 0: mux_27593 = 8'h0; 1: mux_27593 = vout_peek_6004;
    endcase
  endfunction
  wire [7:0] v_27594;
  function [7:0] mux_27594(input [0:0] sel);
    case (sel) 0: mux_27594 = 8'h0; 1: mux_27594 = vout_peek_5995;
    endcase
  endfunction
  wire [7:0] v_27595;
  function [7:0] mux_27595(input [0:0] sel);
    case (sel) 0: mux_27595 = 8'h0; 1: mux_27595 = v_27596;
    endcase
  endfunction
  reg [7:0] v_27596 = 8'h0;
  wire [7:0] v_27597;
  wire [7:0] v_27598;
  function [7:0] mux_27598(input [0:0] sel);
    case (sel) 0: mux_27598 = 8'h0; 1: mux_27598 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27599;
  wire [7:0] v_27600;
  wire [7:0] v_27601;
  function [7:0] mux_27601(input [0:0] sel);
    case (sel) 0: mux_27601 = 8'h0; 1: mux_27601 = vout_peek_5967;
    endcase
  endfunction
  wire [7:0] v_27602;
  function [7:0] mux_27602(input [0:0] sel);
    case (sel) 0: mux_27602 = 8'h0; 1: mux_27602 = vout_peek_5958;
    endcase
  endfunction
  wire [7:0] v_27603;
  function [7:0] mux_27603(input [0:0] sel);
    case (sel) 0: mux_27603 = 8'h0; 1: mux_27603 = v_27604;
    endcase
  endfunction
  reg [7:0] v_27604 = 8'h0;
  wire [7:0] v_27605;
  wire [7:0] v_27606;
  function [7:0] mux_27606(input [0:0] sel);
    case (sel) 0: mux_27606 = 8'h0; 1: mux_27606 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27607;
  wire [7:0] v_27608;
  wire [7:0] v_27609;
  function [7:0] mux_27609(input [0:0] sel);
    case (sel) 0: mux_27609 = 8'h0; 1: mux_27609 = v_27610;
    endcase
  endfunction
  reg [7:0] v_27610 = 8'h0;
  wire [7:0] v_27611;
  wire [7:0] v_27612;
  function [7:0] mux_27612(input [0:0] sel);
    case (sel) 0: mux_27612 = 8'h0; 1: mux_27612 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27613;
  wire [7:0] v_27614;
  wire [7:0] v_27615;
  function [7:0] mux_27615(input [0:0] sel);
    case (sel) 0: mux_27615 = 8'h0; 1: mux_27615 = v_27616;
    endcase
  endfunction
  reg [7:0] v_27616 = 8'h0;
  wire [7:0] v_27617;
  wire [7:0] v_27618;
  function [7:0] mux_27618(input [0:0] sel);
    case (sel) 0: mux_27618 = 8'h0; 1: mux_27618 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27619;
  wire [7:0] v_27620;
  wire [7:0] v_27621;
  function [7:0] mux_27621(input [0:0] sel);
    case (sel) 0: mux_27621 = 8'h0; 1: mux_27621 = vout_peek_5892;
    endcase
  endfunction
  wire [7:0] v_27622;
  function [7:0] mux_27622(input [0:0] sel);
    case (sel) 0: mux_27622 = 8'h0; 1: mux_27622 = vout_peek_5883;
    endcase
  endfunction
  wire [7:0] v_27623;
  function [7:0] mux_27623(input [0:0] sel);
    case (sel) 0: mux_27623 = 8'h0; 1: mux_27623 = v_27624;
    endcase
  endfunction
  reg [7:0] v_27624 = 8'h0;
  wire [7:0] v_27625;
  wire [7:0] v_27626;
  function [7:0] mux_27626(input [0:0] sel);
    case (sel) 0: mux_27626 = 8'h0; 1: mux_27626 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27627;
  wire [7:0] v_27628;
  wire [7:0] v_27629;
  function [7:0] mux_27629(input [0:0] sel);
    case (sel) 0: mux_27629 = 8'h0; 1: mux_27629 = vout_peek_5855;
    endcase
  endfunction
  wire [7:0] v_27630;
  function [7:0] mux_27630(input [0:0] sel);
    case (sel) 0: mux_27630 = 8'h0; 1: mux_27630 = vout_peek_5846;
    endcase
  endfunction
  wire [7:0] v_27631;
  function [7:0] mux_27631(input [0:0] sel);
    case (sel) 0: mux_27631 = 8'h0; 1: mux_27631 = v_27632;
    endcase
  endfunction
  reg [7:0] v_27632 = 8'h0;
  wire [7:0] v_27633;
  wire [7:0] v_27634;
  function [7:0] mux_27634(input [0:0] sel);
    case (sel) 0: mux_27634 = 8'h0; 1: mux_27634 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27635;
  wire [7:0] v_27636;
  wire [7:0] v_27637;
  function [7:0] mux_27637(input [0:0] sel);
    case (sel) 0: mux_27637 = 8'h0; 1: mux_27637 = v_27638;
    endcase
  endfunction
  reg [7:0] v_27638 = 8'h0;
  wire [7:0] v_27639;
  wire [7:0] v_27640;
  function [7:0] mux_27640(input [0:0] sel);
    case (sel) 0: mux_27640 = 8'h0; 1: mux_27640 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27641;
  wire [7:0] v_27642;
  wire [7:0] v_27643;
  function [7:0] mux_27643(input [0:0] sel);
    case (sel) 0: mux_27643 = 8'h0; 1: mux_27643 = vout_peek_5799;
    endcase
  endfunction
  wire [7:0] v_27644;
  function [7:0] mux_27644(input [0:0] sel);
    case (sel) 0: mux_27644 = 8'h0; 1: mux_27644 = vout_peek_5790;
    endcase
  endfunction
  wire [7:0] v_27645;
  function [7:0] mux_27645(input [0:0] sel);
    case (sel) 0: mux_27645 = 8'h0; 1: mux_27645 = v_27646;
    endcase
  endfunction
  reg [7:0] v_27646 = 8'h0;
  wire [7:0] v_27647;
  wire [7:0] v_27648;
  function [7:0] mux_27648(input [0:0] sel);
    case (sel) 0: mux_27648 = 8'h0; 1: mux_27648 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27649;
  wire [7:0] v_27650;
  wire [7:0] v_27651;
  function [7:0] mux_27651(input [0:0] sel);
    case (sel) 0: mux_27651 = 8'h0; 1: mux_27651 = vout_peek_5762;
    endcase
  endfunction
  wire [7:0] v_27652;
  function [7:0] mux_27652(input [0:0] sel);
    case (sel) 0: mux_27652 = 8'h0; 1: mux_27652 = vout_peek_5753;
    endcase
  endfunction
  wire [7:0] v_27653;
  function [7:0] mux_27653(input [0:0] sel);
    case (sel) 0: mux_27653 = 8'h0; 1: mux_27653 = v_27654;
    endcase
  endfunction
  reg [7:0] v_27654 = 8'h0;
  wire [7:0] v_27655;
  wire [7:0] v_27656;
  function [7:0] mux_27656(input [0:0] sel);
    case (sel) 0: mux_27656 = 8'h0; 1: mux_27656 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27657;
  wire [7:0] v_27658;
  wire [7:0] v_27659;
  function [7:0] mux_27659(input [0:0] sel);
    case (sel) 0: mux_27659 = 8'h0; 1: mux_27659 = v_27660;
    endcase
  endfunction
  reg [7:0] v_27660 = 8'h0;
  wire [7:0] v_27661;
  wire [7:0] v_27662;
  function [7:0] mux_27662(input [0:0] sel);
    case (sel) 0: mux_27662 = 8'h0; 1: mux_27662 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27663;
  wire [7:0] v_27664;
  wire [7:0] v_27665;
  function [7:0] mux_27665(input [0:0] sel);
    case (sel) 0: mux_27665 = 8'h0; 1: mux_27665 = v_27666;
    endcase
  endfunction
  reg [7:0] v_27666 = 8'h0;
  wire [7:0] v_27667;
  wire [7:0] v_27668;
  function [7:0] mux_27668(input [0:0] sel);
    case (sel) 0: mux_27668 = 8'h0; 1: mux_27668 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27669;
  wire [7:0] v_27670;
  wire [7:0] v_27671;
  function [7:0] mux_27671(input [0:0] sel);
    case (sel) 0: mux_27671 = 8'h0; 1: mux_27671 = v_27672;
    endcase
  endfunction
  reg [7:0] v_27672 = 8'h0;
  wire [7:0] v_27673;
  wire [7:0] v_27674;
  function [7:0] mux_27674(input [0:0] sel);
    case (sel) 0: mux_27674 = 8'h0; 1: mux_27674 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27675;
  wire [7:0] v_27676;
  wire [7:0] v_27677;
  function [7:0] mux_27677(input [0:0] sel);
    case (sel) 0: mux_27677 = 8'h0; 1: mux_27677 = vout_peek_5668;
    endcase
  endfunction
  wire [7:0] v_27678;
  function [7:0] mux_27678(input [0:0] sel);
    case (sel) 0: mux_27678 = 8'h0; 1: mux_27678 = vout_peek_5659;
    endcase
  endfunction
  wire [7:0] v_27679;
  function [7:0] mux_27679(input [0:0] sel);
    case (sel) 0: mux_27679 = 8'h0; 1: mux_27679 = v_27680;
    endcase
  endfunction
  reg [7:0] v_27680 = 8'h0;
  wire [7:0] v_27681;
  wire [7:0] v_27682;
  function [7:0] mux_27682(input [0:0] sel);
    case (sel) 0: mux_27682 = 8'h0; 1: mux_27682 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27683;
  wire [7:0] v_27684;
  wire [7:0] v_27685;
  function [7:0] mux_27685(input [0:0] sel);
    case (sel) 0: mux_27685 = 8'h0; 1: mux_27685 = vout_peek_5631;
    endcase
  endfunction
  wire [7:0] v_27686;
  function [7:0] mux_27686(input [0:0] sel);
    case (sel) 0: mux_27686 = 8'h0; 1: mux_27686 = vout_peek_5622;
    endcase
  endfunction
  wire [7:0] v_27687;
  function [7:0] mux_27687(input [0:0] sel);
    case (sel) 0: mux_27687 = 8'h0; 1: mux_27687 = v_27688;
    endcase
  endfunction
  reg [7:0] v_27688 = 8'h0;
  wire [7:0] v_27689;
  wire [7:0] v_27690;
  function [7:0] mux_27690(input [0:0] sel);
    case (sel) 0: mux_27690 = 8'h0; 1: mux_27690 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27691;
  wire [7:0] v_27692;
  wire [7:0] v_27693;
  function [7:0] mux_27693(input [0:0] sel);
    case (sel) 0: mux_27693 = 8'h0; 1: mux_27693 = v_27694;
    endcase
  endfunction
  reg [7:0] v_27694 = 8'h0;
  wire [7:0] v_27695;
  wire [7:0] v_27696;
  function [7:0] mux_27696(input [0:0] sel);
    case (sel) 0: mux_27696 = 8'h0; 1: mux_27696 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27697;
  wire [7:0] v_27698;
  wire [7:0] v_27699;
  function [7:0] mux_27699(input [0:0] sel);
    case (sel) 0: mux_27699 = 8'h0; 1: mux_27699 = vout_peek_5575;
    endcase
  endfunction
  wire [7:0] v_27700;
  function [7:0] mux_27700(input [0:0] sel);
    case (sel) 0: mux_27700 = 8'h0; 1: mux_27700 = vout_peek_5566;
    endcase
  endfunction
  wire [7:0] v_27701;
  function [7:0] mux_27701(input [0:0] sel);
    case (sel) 0: mux_27701 = 8'h0; 1: mux_27701 = v_27702;
    endcase
  endfunction
  reg [7:0] v_27702 = 8'h0;
  wire [7:0] v_27703;
  wire [7:0] v_27704;
  function [7:0] mux_27704(input [0:0] sel);
    case (sel) 0: mux_27704 = 8'h0; 1: mux_27704 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27705;
  wire [7:0] v_27706;
  wire [7:0] v_27707;
  function [7:0] mux_27707(input [0:0] sel);
    case (sel) 0: mux_27707 = 8'h0; 1: mux_27707 = vout_peek_5538;
    endcase
  endfunction
  wire [7:0] v_27708;
  function [7:0] mux_27708(input [0:0] sel);
    case (sel) 0: mux_27708 = 8'h0; 1: mux_27708 = vout_peek_5529;
    endcase
  endfunction
  wire [7:0] v_27709;
  function [7:0] mux_27709(input [0:0] sel);
    case (sel) 0: mux_27709 = 8'h0; 1: mux_27709 = v_27710;
    endcase
  endfunction
  reg [7:0] v_27710 = 8'h0;
  wire [7:0] v_27711;
  wire [7:0] v_27712;
  function [7:0] mux_27712(input [0:0] sel);
    case (sel) 0: mux_27712 = 8'h0; 1: mux_27712 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27713;
  wire [7:0] v_27714;
  wire [7:0] v_27715;
  function [7:0] mux_27715(input [0:0] sel);
    case (sel) 0: mux_27715 = 8'h0; 1: mux_27715 = v_27716;
    endcase
  endfunction
  reg [7:0] v_27716 = 8'h0;
  wire [7:0] v_27717;
  wire [7:0] v_27718;
  function [7:0] mux_27718(input [0:0] sel);
    case (sel) 0: mux_27718 = 8'h0; 1: mux_27718 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27719;
  wire [7:0] v_27720;
  wire [7:0] v_27721;
  function [7:0] mux_27721(input [0:0] sel);
    case (sel) 0: mux_27721 = 8'h0; 1: mux_27721 = v_27722;
    endcase
  endfunction
  reg [7:0] v_27722 = 8'h0;
  wire [7:0] v_27723;
  wire [7:0] v_27724;
  function [7:0] mux_27724(input [0:0] sel);
    case (sel) 0: mux_27724 = 8'h0; 1: mux_27724 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27725;
  wire [7:0] v_27726;
  wire [7:0] v_27727;
  function [7:0] mux_27727(input [0:0] sel);
    case (sel) 0: mux_27727 = 8'h0; 1: mux_27727 = vout_peek_5463;
    endcase
  endfunction
  wire [7:0] v_27728;
  function [7:0] mux_27728(input [0:0] sel);
    case (sel) 0: mux_27728 = 8'h0; 1: mux_27728 = vout_peek_5454;
    endcase
  endfunction
  wire [7:0] v_27729;
  function [7:0] mux_27729(input [0:0] sel);
    case (sel) 0: mux_27729 = 8'h0; 1: mux_27729 = v_27730;
    endcase
  endfunction
  reg [7:0] v_27730 = 8'h0;
  wire [7:0] v_27731;
  wire [7:0] v_27732;
  function [7:0] mux_27732(input [0:0] sel);
    case (sel) 0: mux_27732 = 8'h0; 1: mux_27732 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27733;
  wire [7:0] v_27734;
  wire [7:0] v_27735;
  function [7:0] mux_27735(input [0:0] sel);
    case (sel) 0: mux_27735 = 8'h0; 1: mux_27735 = vout_peek_5426;
    endcase
  endfunction
  wire [7:0] v_27736;
  function [7:0] mux_27736(input [0:0] sel);
    case (sel) 0: mux_27736 = 8'h0; 1: mux_27736 = vout_peek_5417;
    endcase
  endfunction
  wire [7:0] v_27737;
  function [7:0] mux_27737(input [0:0] sel);
    case (sel) 0: mux_27737 = 8'h0; 1: mux_27737 = v_27738;
    endcase
  endfunction
  reg [7:0] v_27738 = 8'h0;
  wire [7:0] v_27739;
  wire [7:0] v_27740;
  function [7:0] mux_27740(input [0:0] sel);
    case (sel) 0: mux_27740 = 8'h0; 1: mux_27740 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27741;
  wire [7:0] v_27742;
  wire [7:0] v_27743;
  function [7:0] mux_27743(input [0:0] sel);
    case (sel) 0: mux_27743 = 8'h0; 1: mux_27743 = v_27744;
    endcase
  endfunction
  reg [7:0] v_27744 = 8'h0;
  wire [7:0] v_27745;
  wire [7:0] v_27746;
  function [7:0] mux_27746(input [0:0] sel);
    case (sel) 0: mux_27746 = 8'h0; 1: mux_27746 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27747;
  wire [7:0] v_27748;
  wire [7:0] v_27749;
  function [7:0] mux_27749(input [0:0] sel);
    case (sel) 0: mux_27749 = 8'h0; 1: mux_27749 = vout_peek_5370;
    endcase
  endfunction
  wire [7:0] v_27750;
  function [7:0] mux_27750(input [0:0] sel);
    case (sel) 0: mux_27750 = 8'h0; 1: mux_27750 = vout_peek_5361;
    endcase
  endfunction
  wire [7:0] v_27751;
  function [7:0] mux_27751(input [0:0] sel);
    case (sel) 0: mux_27751 = 8'h0; 1: mux_27751 = v_27752;
    endcase
  endfunction
  reg [7:0] v_27752 = 8'h0;
  wire [7:0] v_27753;
  wire [7:0] v_27754;
  function [7:0] mux_27754(input [0:0] sel);
    case (sel) 0: mux_27754 = 8'h0; 1: mux_27754 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27755;
  wire [7:0] v_27756;
  wire [7:0] v_27757;
  function [7:0] mux_27757(input [0:0] sel);
    case (sel) 0: mux_27757 = 8'h0; 1: mux_27757 = vout_peek_5333;
    endcase
  endfunction
  wire [7:0] v_27758;
  function [7:0] mux_27758(input [0:0] sel);
    case (sel) 0: mux_27758 = 8'h0; 1: mux_27758 = vout_peek_5324;
    endcase
  endfunction
  wire [7:0] v_27759;
  function [7:0] mux_27759(input [0:0] sel);
    case (sel) 0: mux_27759 = 8'h0; 1: mux_27759 = v_27760;
    endcase
  endfunction
  reg [7:0] v_27760 = 8'h0;
  wire [7:0] v_27761;
  wire [7:0] v_27762;
  function [7:0] mux_27762(input [0:0] sel);
    case (sel) 0: mux_27762 = 8'h0; 1: mux_27762 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27763;
  wire [7:0] v_27764;
  wire [7:0] v_27765;
  function [7:0] mux_27765(input [0:0] sel);
    case (sel) 0: mux_27765 = 8'h0; 1: mux_27765 = v_27766;
    endcase
  endfunction
  reg [7:0] v_27766 = 8'h0;
  wire [7:0] v_27767;
  wire [7:0] v_27768;
  function [7:0] mux_27768(input [0:0] sel);
    case (sel) 0: mux_27768 = 8'h0; 1: mux_27768 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27769;
  wire [7:0] v_27770;
  wire [7:0] v_27771;
  function [7:0] mux_27771(input [0:0] sel);
    case (sel) 0: mux_27771 = 8'h0; 1: mux_27771 = v_27772;
    endcase
  endfunction
  reg [7:0] v_27772 = 8'h0;
  wire [7:0] v_27773;
  wire [7:0] v_27774;
  function [7:0] mux_27774(input [0:0] sel);
    case (sel) 0: mux_27774 = 8'h0; 1: mux_27774 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27775;
  wire [7:0] v_27776;
  wire [7:0] v_27777;
  function [7:0] mux_27777(input [0:0] sel);
    case (sel) 0: mux_27777 = 8'h0; 1: mux_27777 = v_27778;
    endcase
  endfunction
  reg [7:0] v_27778 = 8'h0;
  wire [7:0] v_27779;
  wire [7:0] v_27780;
  function [7:0] mux_27780(input [0:0] sel);
    case (sel) 0: mux_27780 = 8'h0; 1: mux_27780 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27781;
  wire [7:0] v_27782;
  wire [7:0] v_27783;
  function [7:0] mux_27783(input [0:0] sel);
    case (sel) 0: mux_27783 = 8'h0; 1: mux_27783 = v_27784;
    endcase
  endfunction
  reg [7:0] v_27784 = 8'h0;
  wire [7:0] v_27785;
  wire [7:0] v_27786;
  function [7:0] mux_27786(input [0:0] sel);
    case (sel) 0: mux_27786 = 8'h0; 1: mux_27786 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27787;
  wire [7:0] v_27788;
  wire [7:0] v_27789;
  function [7:0] mux_27789(input [0:0] sel);
    case (sel) 0: mux_27789 = 8'h0; 1: mux_27789 = vout_peek_5220;
    endcase
  endfunction
  wire [7:0] v_27790;
  function [7:0] mux_27790(input [0:0] sel);
    case (sel) 0: mux_27790 = 8'h0; 1: mux_27790 = vout_peek_5211;
    endcase
  endfunction
  wire [7:0] v_27791;
  function [7:0] mux_27791(input [0:0] sel);
    case (sel) 0: mux_27791 = 8'h0; 1: mux_27791 = v_27792;
    endcase
  endfunction
  reg [7:0] v_27792 = 8'h0;
  wire [7:0] v_27793;
  wire [7:0] v_27794;
  function [7:0] mux_27794(input [0:0] sel);
    case (sel) 0: mux_27794 = 8'h0; 1: mux_27794 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27795;
  wire [7:0] v_27796;
  wire [7:0] v_27797;
  function [7:0] mux_27797(input [0:0] sel);
    case (sel) 0: mux_27797 = 8'h0; 1: mux_27797 = vout_peek_5183;
    endcase
  endfunction
  wire [7:0] v_27798;
  function [7:0] mux_27798(input [0:0] sel);
    case (sel) 0: mux_27798 = 8'h0; 1: mux_27798 = vout_peek_5174;
    endcase
  endfunction
  wire [7:0] v_27799;
  function [7:0] mux_27799(input [0:0] sel);
    case (sel) 0: mux_27799 = 8'h0; 1: mux_27799 = v_27800;
    endcase
  endfunction
  reg [7:0] v_27800 = 8'h0;
  wire [7:0] v_27801;
  wire [7:0] v_27802;
  function [7:0] mux_27802(input [0:0] sel);
    case (sel) 0: mux_27802 = 8'h0; 1: mux_27802 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27803;
  wire [7:0] v_27804;
  wire [7:0] v_27805;
  function [7:0] mux_27805(input [0:0] sel);
    case (sel) 0: mux_27805 = 8'h0; 1: mux_27805 = v_27806;
    endcase
  endfunction
  reg [7:0] v_27806 = 8'h0;
  wire [7:0] v_27807;
  wire [7:0] v_27808;
  function [7:0] mux_27808(input [0:0] sel);
    case (sel) 0: mux_27808 = 8'h0; 1: mux_27808 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27809;
  wire [7:0] v_27810;
  wire [7:0] v_27811;
  function [7:0] mux_27811(input [0:0] sel);
    case (sel) 0: mux_27811 = 8'h0; 1: mux_27811 = vout_peek_5127;
    endcase
  endfunction
  wire [7:0] v_27812;
  function [7:0] mux_27812(input [0:0] sel);
    case (sel) 0: mux_27812 = 8'h0; 1: mux_27812 = vout_peek_5118;
    endcase
  endfunction
  wire [7:0] v_27813;
  function [7:0] mux_27813(input [0:0] sel);
    case (sel) 0: mux_27813 = 8'h0; 1: mux_27813 = v_27814;
    endcase
  endfunction
  reg [7:0] v_27814 = 8'h0;
  wire [7:0] v_27815;
  wire [7:0] v_27816;
  function [7:0] mux_27816(input [0:0] sel);
    case (sel) 0: mux_27816 = 8'h0; 1: mux_27816 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27817;
  wire [7:0] v_27818;
  wire [7:0] v_27819;
  function [7:0] mux_27819(input [0:0] sel);
    case (sel) 0: mux_27819 = 8'h0; 1: mux_27819 = vout_peek_5090;
    endcase
  endfunction
  wire [7:0] v_27820;
  function [7:0] mux_27820(input [0:0] sel);
    case (sel) 0: mux_27820 = 8'h0; 1: mux_27820 = vout_peek_5081;
    endcase
  endfunction
  wire [7:0] v_27821;
  function [7:0] mux_27821(input [0:0] sel);
    case (sel) 0: mux_27821 = 8'h0; 1: mux_27821 = v_27822;
    endcase
  endfunction
  reg [7:0] v_27822 = 8'h0;
  wire [7:0] v_27823;
  wire [7:0] v_27824;
  function [7:0] mux_27824(input [0:0] sel);
    case (sel) 0: mux_27824 = 8'h0; 1: mux_27824 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27825;
  wire [7:0] v_27826;
  wire [7:0] v_27827;
  function [7:0] mux_27827(input [0:0] sel);
    case (sel) 0: mux_27827 = 8'h0; 1: mux_27827 = v_27828;
    endcase
  endfunction
  reg [7:0] v_27828 = 8'h0;
  wire [7:0] v_27829;
  wire [7:0] v_27830;
  function [7:0] mux_27830(input [0:0] sel);
    case (sel) 0: mux_27830 = 8'h0; 1: mux_27830 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27831;
  wire [7:0] v_27832;
  wire [7:0] v_27833;
  function [7:0] mux_27833(input [0:0] sel);
    case (sel) 0: mux_27833 = 8'h0; 1: mux_27833 = v_27834;
    endcase
  endfunction
  reg [7:0] v_27834 = 8'h0;
  wire [7:0] v_27835;
  wire [7:0] v_27836;
  function [7:0] mux_27836(input [0:0] sel);
    case (sel) 0: mux_27836 = 8'h0; 1: mux_27836 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27837;
  wire [7:0] v_27838;
  wire [7:0] v_27839;
  function [7:0] mux_27839(input [0:0] sel);
    case (sel) 0: mux_27839 = 8'h0; 1: mux_27839 = vout_peek_5015;
    endcase
  endfunction
  wire [7:0] v_27840;
  function [7:0] mux_27840(input [0:0] sel);
    case (sel) 0: mux_27840 = 8'h0; 1: mux_27840 = vout_peek_5006;
    endcase
  endfunction
  wire [7:0] v_27841;
  function [7:0] mux_27841(input [0:0] sel);
    case (sel) 0: mux_27841 = 8'h0; 1: mux_27841 = v_27842;
    endcase
  endfunction
  reg [7:0] v_27842 = 8'h0;
  wire [7:0] v_27843;
  wire [7:0] v_27844;
  function [7:0] mux_27844(input [0:0] sel);
    case (sel) 0: mux_27844 = 8'h0; 1: mux_27844 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27845;
  wire [7:0] v_27846;
  wire [7:0] v_27847;
  function [7:0] mux_27847(input [0:0] sel);
    case (sel) 0: mux_27847 = 8'h0; 1: mux_27847 = vout_peek_4978;
    endcase
  endfunction
  wire [7:0] v_27848;
  function [7:0] mux_27848(input [0:0] sel);
    case (sel) 0: mux_27848 = 8'h0; 1: mux_27848 = vout_peek_4969;
    endcase
  endfunction
  wire [7:0] v_27849;
  function [7:0] mux_27849(input [0:0] sel);
    case (sel) 0: mux_27849 = 8'h0; 1: mux_27849 = v_27850;
    endcase
  endfunction
  reg [7:0] v_27850 = 8'h0;
  wire [7:0] v_27851;
  wire [7:0] v_27852;
  function [7:0] mux_27852(input [0:0] sel);
    case (sel) 0: mux_27852 = 8'h0; 1: mux_27852 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27853;
  wire [7:0] v_27854;
  wire [7:0] v_27855;
  function [7:0] mux_27855(input [0:0] sel);
    case (sel) 0: mux_27855 = 8'h0; 1: mux_27855 = v_27856;
    endcase
  endfunction
  reg [7:0] v_27856 = 8'h0;
  wire [7:0] v_27857;
  wire [7:0] v_27858;
  function [7:0] mux_27858(input [0:0] sel);
    case (sel) 0: mux_27858 = 8'h0; 1: mux_27858 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27859;
  wire [7:0] v_27860;
  wire [7:0] v_27861;
  function [7:0] mux_27861(input [0:0] sel);
    case (sel) 0: mux_27861 = 8'h0; 1: mux_27861 = vout_peek_4922;
    endcase
  endfunction
  wire [7:0] v_27862;
  function [7:0] mux_27862(input [0:0] sel);
    case (sel) 0: mux_27862 = 8'h0; 1: mux_27862 = vout_peek_4913;
    endcase
  endfunction
  wire [7:0] v_27863;
  function [7:0] mux_27863(input [0:0] sel);
    case (sel) 0: mux_27863 = 8'h0; 1: mux_27863 = v_27864;
    endcase
  endfunction
  reg [7:0] v_27864 = 8'h0;
  wire [7:0] v_27865;
  wire [7:0] v_27866;
  function [7:0] mux_27866(input [0:0] sel);
    case (sel) 0: mux_27866 = 8'h0; 1: mux_27866 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27867;
  wire [7:0] v_27868;
  wire [7:0] v_27869;
  function [7:0] mux_27869(input [0:0] sel);
    case (sel) 0: mux_27869 = 8'h0; 1: mux_27869 = vout_peek_4885;
    endcase
  endfunction
  wire [7:0] v_27870;
  function [7:0] mux_27870(input [0:0] sel);
    case (sel) 0: mux_27870 = 8'h0; 1: mux_27870 = vout_peek_4876;
    endcase
  endfunction
  wire [7:0] v_27871;
  function [7:0] mux_27871(input [0:0] sel);
    case (sel) 0: mux_27871 = 8'h0; 1: mux_27871 = v_27872;
    endcase
  endfunction
  reg [7:0] v_27872 = 8'h0;
  wire [7:0] v_27873;
  wire [7:0] v_27874;
  function [7:0] mux_27874(input [0:0] sel);
    case (sel) 0: mux_27874 = 8'h0; 1: mux_27874 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27875;
  wire [7:0] v_27876;
  wire [7:0] v_27877;
  function [7:0] mux_27877(input [0:0] sel);
    case (sel) 0: mux_27877 = 8'h0; 1: mux_27877 = v_27878;
    endcase
  endfunction
  reg [7:0] v_27878 = 8'h0;
  wire [7:0] v_27879;
  wire [7:0] v_27880;
  function [7:0] mux_27880(input [0:0] sel);
    case (sel) 0: mux_27880 = 8'h0; 1: mux_27880 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27881;
  wire [7:0] v_27882;
  wire [7:0] v_27883;
  function [7:0] mux_27883(input [0:0] sel);
    case (sel) 0: mux_27883 = 8'h0; 1: mux_27883 = v_27884;
    endcase
  endfunction
  reg [7:0] v_27884 = 8'h0;
  wire [7:0] v_27885;
  wire [7:0] v_27886;
  function [7:0] mux_27886(input [0:0] sel);
    case (sel) 0: mux_27886 = 8'h0; 1: mux_27886 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27887;
  wire [7:0] v_27888;
  wire [7:0] v_27889;
  function [7:0] mux_27889(input [0:0] sel);
    case (sel) 0: mux_27889 = 8'h0; 1: mux_27889 = v_27890;
    endcase
  endfunction
  reg [7:0] v_27890 = 8'h0;
  wire [7:0] v_27891;
  wire [7:0] v_27892;
  function [7:0] mux_27892(input [0:0] sel);
    case (sel) 0: mux_27892 = 8'h0; 1: mux_27892 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27893;
  wire [7:0] v_27894;
  wire [7:0] v_27895;
  function [7:0] mux_27895(input [0:0] sel);
    case (sel) 0: mux_27895 = 8'h0; 1: mux_27895 = vout_peek_4791;
    endcase
  endfunction
  wire [7:0] v_27896;
  function [7:0] mux_27896(input [0:0] sel);
    case (sel) 0: mux_27896 = 8'h0; 1: mux_27896 = vout_peek_4782;
    endcase
  endfunction
  wire [7:0] v_27897;
  function [7:0] mux_27897(input [0:0] sel);
    case (sel) 0: mux_27897 = 8'h0; 1: mux_27897 = v_27898;
    endcase
  endfunction
  reg [7:0] v_27898 = 8'h0;
  wire [7:0] v_27899;
  wire [7:0] v_27900;
  function [7:0] mux_27900(input [0:0] sel);
    case (sel) 0: mux_27900 = 8'h0; 1: mux_27900 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27901;
  wire [7:0] v_27902;
  wire [7:0] v_27903;
  function [7:0] mux_27903(input [0:0] sel);
    case (sel) 0: mux_27903 = 8'h0; 1: mux_27903 = vout_peek_4754;
    endcase
  endfunction
  wire [7:0] v_27904;
  function [7:0] mux_27904(input [0:0] sel);
    case (sel) 0: mux_27904 = 8'h0; 1: mux_27904 = vout_peek_4745;
    endcase
  endfunction
  wire [7:0] v_27905;
  function [7:0] mux_27905(input [0:0] sel);
    case (sel) 0: mux_27905 = 8'h0; 1: mux_27905 = v_27906;
    endcase
  endfunction
  reg [7:0] v_27906 = 8'h0;
  wire [7:0] v_27907;
  wire [7:0] v_27908;
  function [7:0] mux_27908(input [0:0] sel);
    case (sel) 0: mux_27908 = 8'h0; 1: mux_27908 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27909;
  wire [7:0] v_27910;
  wire [7:0] v_27911;
  function [7:0] mux_27911(input [0:0] sel);
    case (sel) 0: mux_27911 = 8'h0; 1: mux_27911 = v_27912;
    endcase
  endfunction
  reg [7:0] v_27912 = 8'h0;
  wire [7:0] v_27913;
  wire [7:0] v_27914;
  function [7:0] mux_27914(input [0:0] sel);
    case (sel) 0: mux_27914 = 8'h0; 1: mux_27914 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27915;
  wire [7:0] v_27916;
  wire [7:0] v_27917;
  function [7:0] mux_27917(input [0:0] sel);
    case (sel) 0: mux_27917 = 8'h0; 1: mux_27917 = vout_peek_4698;
    endcase
  endfunction
  wire [7:0] v_27918;
  function [7:0] mux_27918(input [0:0] sel);
    case (sel) 0: mux_27918 = 8'h0; 1: mux_27918 = vout_peek_4689;
    endcase
  endfunction
  wire [7:0] v_27919;
  function [7:0] mux_27919(input [0:0] sel);
    case (sel) 0: mux_27919 = 8'h0; 1: mux_27919 = v_27920;
    endcase
  endfunction
  reg [7:0] v_27920 = 8'h0;
  wire [7:0] v_27921;
  wire [7:0] v_27922;
  function [7:0] mux_27922(input [0:0] sel);
    case (sel) 0: mux_27922 = 8'h0; 1: mux_27922 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27923;
  wire [7:0] v_27924;
  wire [7:0] v_27925;
  function [7:0] mux_27925(input [0:0] sel);
    case (sel) 0: mux_27925 = 8'h0; 1: mux_27925 = vout_peek_4661;
    endcase
  endfunction
  wire [7:0] v_27926;
  function [7:0] mux_27926(input [0:0] sel);
    case (sel) 0: mux_27926 = 8'h0; 1: mux_27926 = vout_peek_4652;
    endcase
  endfunction
  wire [7:0] v_27927;
  function [7:0] mux_27927(input [0:0] sel);
    case (sel) 0: mux_27927 = 8'h0; 1: mux_27927 = v_27928;
    endcase
  endfunction
  reg [7:0] v_27928 = 8'h0;
  wire [7:0] v_27929;
  wire [7:0] v_27930;
  function [7:0] mux_27930(input [0:0] sel);
    case (sel) 0: mux_27930 = 8'h0; 1: mux_27930 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27931;
  wire [7:0] v_27932;
  wire [7:0] v_27933;
  function [7:0] mux_27933(input [0:0] sel);
    case (sel) 0: mux_27933 = 8'h0; 1: mux_27933 = v_27934;
    endcase
  endfunction
  reg [7:0] v_27934 = 8'h0;
  wire [7:0] v_27935;
  wire [7:0] v_27936;
  function [7:0] mux_27936(input [0:0] sel);
    case (sel) 0: mux_27936 = 8'h0; 1: mux_27936 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27937;
  wire [7:0] v_27938;
  wire [7:0] v_27939;
  function [7:0] mux_27939(input [0:0] sel);
    case (sel) 0: mux_27939 = 8'h0; 1: mux_27939 = v_27940;
    endcase
  endfunction
  reg [7:0] v_27940 = 8'h0;
  wire [7:0] v_27941;
  wire [7:0] v_27942;
  function [7:0] mux_27942(input [0:0] sel);
    case (sel) 0: mux_27942 = 8'h0; 1: mux_27942 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27943;
  wire [7:0] v_27944;
  wire [7:0] v_27945;
  function [7:0] mux_27945(input [0:0] sel);
    case (sel) 0: mux_27945 = 8'h0; 1: mux_27945 = vout_peek_4586;
    endcase
  endfunction
  wire [7:0] v_27946;
  function [7:0] mux_27946(input [0:0] sel);
    case (sel) 0: mux_27946 = 8'h0; 1: mux_27946 = vout_peek_4577;
    endcase
  endfunction
  wire [7:0] v_27947;
  function [7:0] mux_27947(input [0:0] sel);
    case (sel) 0: mux_27947 = 8'h0; 1: mux_27947 = v_27948;
    endcase
  endfunction
  reg [7:0] v_27948 = 8'h0;
  wire [7:0] v_27949;
  wire [7:0] v_27950;
  function [7:0] mux_27950(input [0:0] sel);
    case (sel) 0: mux_27950 = 8'h0; 1: mux_27950 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27951;
  wire [7:0] v_27952;
  wire [7:0] v_27953;
  function [7:0] mux_27953(input [0:0] sel);
    case (sel) 0: mux_27953 = 8'h0; 1: mux_27953 = vout_peek_4549;
    endcase
  endfunction
  wire [7:0] v_27954;
  function [7:0] mux_27954(input [0:0] sel);
    case (sel) 0: mux_27954 = 8'h0; 1: mux_27954 = vout_peek_4540;
    endcase
  endfunction
  wire [7:0] v_27955;
  function [7:0] mux_27955(input [0:0] sel);
    case (sel) 0: mux_27955 = 8'h0; 1: mux_27955 = v_27956;
    endcase
  endfunction
  reg [7:0] v_27956 = 8'h0;
  wire [7:0] v_27957;
  wire [7:0] v_27958;
  function [7:0] mux_27958(input [0:0] sel);
    case (sel) 0: mux_27958 = 8'h0; 1: mux_27958 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27959;
  wire [7:0] v_27960;
  wire [7:0] v_27961;
  function [7:0] mux_27961(input [0:0] sel);
    case (sel) 0: mux_27961 = 8'h0; 1: mux_27961 = v_27962;
    endcase
  endfunction
  reg [7:0] v_27962 = 8'h0;
  wire [7:0] v_27963;
  wire [7:0] v_27964;
  function [7:0] mux_27964(input [0:0] sel);
    case (sel) 0: mux_27964 = 8'h0; 1: mux_27964 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27965;
  wire [7:0] v_27966;
  wire [7:0] v_27967;
  function [7:0] mux_27967(input [0:0] sel);
    case (sel) 0: mux_27967 = 8'h0; 1: mux_27967 = vout_peek_4493;
    endcase
  endfunction
  wire [7:0] v_27968;
  function [7:0] mux_27968(input [0:0] sel);
    case (sel) 0: mux_27968 = 8'h0; 1: mux_27968 = vout_peek_4484;
    endcase
  endfunction
  wire [7:0] v_27969;
  function [7:0] mux_27969(input [0:0] sel);
    case (sel) 0: mux_27969 = 8'h0; 1: mux_27969 = v_27970;
    endcase
  endfunction
  reg [7:0] v_27970 = 8'h0;
  wire [7:0] v_27971;
  wire [7:0] v_27972;
  function [7:0] mux_27972(input [0:0] sel);
    case (sel) 0: mux_27972 = 8'h0; 1: mux_27972 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_27973;
  wire [7:0] v_27974;
  wire [7:0] v_27975;
  function [7:0] mux_27975(input [0:0] sel);
    case (sel) 0: mux_27975 = 8'h0; 1: mux_27975 = vout_peek_4456;
    endcase
  endfunction
  wire [7:0] v_27976;
  function [7:0] mux_27976(input [0:0] sel);
    case (sel) 0: mux_27976 = 8'h0; 1: mux_27976 = vout_peek_4447;
    endcase
  endfunction
  wire [0:0] v_27977;
  wire [7:0] v_27978;
  // Instances
  //////////////////////////////////////////////////////////////////////////////
  assign v_0 = v_1 | v_22377;
  assign v_1 = mux_1(v_2);
  assign v_2 = vout_canPeek_3 & v_4;
  pebbles_core
    pebbles_core_3
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_0),
       .in0_consume_en(vin0_consume_en_3),
       .out_canPeek(vout_canPeek_3),
       .out_peek(vout_peek_3));
  assign v_4 = v_5 & 1'h1;
  assign v_5 = v_6 | 1'h0;
  assign v_6 = ~v_7;
  assign v_8 = v_9 | v_19;
  assign v_9 = act_10 & 1'h1;
  assign act_10 = v_11 | v_2;
  assign v_11 = v_12 & v_4;
  assign v_12 = v_13 & vout_canPeek_14;
  assign v_13 = ~vout_canPeek_3;
  pebbles_core
    pebbles_core_14
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15),
       .in0_consume_en(vin0_consume_en_14),
       .out_canPeek(vout_canPeek_14),
       .out_peek(vout_peek_14));
  assign v_15 = v_16 | v_17;
  assign v_16 = mux_16(v_11);
  assign v_17 = mux_17(v_18);
  assign v_18 = ~v_11;
  assign v_19 = v_20 & 1'h1;
  assign v_20 = v_21 & v_22;
  assign v_21 = ~act_10;
  assign v_22 = v_23 | v_22373;
  assign v_23 = v_24 | v_22371;
  assign v_24 = mux_24(v_25);
  assign v_25 = v_7 & v_26;
  assign v_26 = v_27 & 1'h1;
  assign v_27 = v_28 | 1'h0;
  assign v_28 = ~v_29;
  assign v_30 = v_31 | v_69;
  assign v_31 = act_32 & 1'h1;
  assign act_32 = v_33 | v_25;
  assign v_33 = v_34 & v_26;
  assign v_34 = v_35 & v_36;
  assign v_35 = ~v_7;
  assign v_37 = v_38 | v_57;
  assign v_38 = act_39 & 1'h1;
  assign act_39 = v_40 | v_46;
  assign v_40 = v_41 & v_47;
  assign v_41 = v_42 & vout_canPeek_52;
  assign v_42 = ~vout_canPeek_43;
  pebbles_core
    pebbles_core_43
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_44),
       .in0_consume_en(vin0_consume_en_43),
       .out_canPeek(vout_canPeek_43),
       .out_peek(vout_peek_43));
  assign v_44 = v_45 | v_50;
  assign v_45 = mux_45(v_46);
  assign v_46 = vout_canPeek_43 & v_47;
  assign v_47 = v_48 & 1'h1;
  assign v_48 = v_49 | 1'h0;
  assign v_49 = ~v_36;
  assign v_50 = mux_50(v_51);
  assign v_51 = ~v_46;
  pebbles_core
    pebbles_core_52
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_53),
       .in0_consume_en(vin0_consume_en_52),
       .out_canPeek(vout_canPeek_52),
       .out_peek(vout_peek_52));
  assign v_53 = v_54 | v_55;
  assign v_54 = mux_54(v_40);
  assign v_55 = mux_55(v_56);
  assign v_56 = ~v_40;
  assign v_57 = v_58 & 1'h1;
  assign v_58 = v_59 & v_60;
  assign v_59 = ~act_39;
  assign v_60 = v_61 | v_65;
  assign v_61 = v_62 | v_63;
  assign v_62 = mux_62(v_33);
  assign v_63 = mux_63(v_64);
  assign v_64 = ~v_33;
  assign v_65 = ~v_36;
  assign v_66 = v_67 | v_68;
  assign v_67 = mux_67(v_38);
  assign v_68 = mux_68(v_57);
  assign v_69 = v_70 & 1'h1;
  assign v_70 = v_71 & v_72;
  assign v_71 = ~act_32;
  assign v_72 = v_73 | v_22367;
  assign v_73 = v_74 | v_22365;
  assign v_74 = mux_74(v_75);
  assign v_75 = v_29 & v_76;
  assign v_76 = v_77 & 1'h1;
  assign v_77 = v_78 | 1'h0;
  assign v_78 = ~v_79;
  assign v_80 = v_81 | v_175;
  assign v_81 = act_82 & 1'h1;
  assign act_82 = v_83 | v_75;
  assign v_83 = v_84 & v_76;
  assign v_84 = v_85 & v_86;
  assign v_85 = ~v_29;
  assign v_87 = v_88 | v_163;
  assign v_88 = act_89 & 1'h1;
  assign act_89 = v_90 | v_120;
  assign v_90 = v_91 & v_121;
  assign v_91 = v_92 & v_130;
  assign v_92 = ~v_93;
  assign v_94 = v_95 | v_114;
  assign v_95 = act_96 & 1'h1;
  assign act_96 = v_97 | v_103;
  assign v_97 = v_98 & v_104;
  assign v_98 = v_99 & vout_canPeek_109;
  assign v_99 = ~vout_canPeek_100;
  pebbles_core
    pebbles_core_100
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_101),
       .in0_consume_en(vin0_consume_en_100),
       .out_canPeek(vout_canPeek_100),
       .out_peek(vout_peek_100));
  assign v_101 = v_102 | v_107;
  assign v_102 = mux_102(v_103);
  assign v_103 = vout_canPeek_100 & v_104;
  assign v_104 = v_105 & 1'h1;
  assign v_105 = v_106 | 1'h0;
  assign v_106 = ~v_93;
  assign v_107 = mux_107(v_108);
  assign v_108 = ~v_103;
  pebbles_core
    pebbles_core_109
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_110),
       .in0_consume_en(vin0_consume_en_109),
       .out_canPeek(vout_canPeek_109),
       .out_peek(vout_peek_109));
  assign v_110 = v_111 | v_112;
  assign v_111 = mux_111(v_97);
  assign v_112 = mux_112(v_113);
  assign v_113 = ~v_97;
  assign v_114 = v_115 & 1'h1;
  assign v_115 = v_116 & v_117;
  assign v_116 = ~act_96;
  assign v_117 = v_118 | v_126;
  assign v_118 = v_119 | v_124;
  assign v_119 = mux_119(v_120);
  assign v_120 = v_93 & v_121;
  assign v_121 = v_122 & 1'h1;
  assign v_122 = v_123 | 1'h0;
  assign v_123 = ~v_86;
  assign v_124 = mux_124(v_125);
  assign v_125 = ~v_120;
  assign v_126 = ~v_93;
  assign v_127 = v_128 | v_129;
  assign v_128 = mux_128(v_95);
  assign v_129 = mux_129(v_114);
  assign v_131 = v_132 | v_151;
  assign v_132 = act_133 & 1'h1;
  assign act_133 = v_134 | v_140;
  assign v_134 = v_135 & v_141;
  assign v_135 = v_136 & vout_canPeek_146;
  assign v_136 = ~vout_canPeek_137;
  pebbles_core
    pebbles_core_137
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_138),
       .in0_consume_en(vin0_consume_en_137),
       .out_canPeek(vout_canPeek_137),
       .out_peek(vout_peek_137));
  assign v_138 = v_139 | v_144;
  assign v_139 = mux_139(v_140);
  assign v_140 = vout_canPeek_137 & v_141;
  assign v_141 = v_142 & 1'h1;
  assign v_142 = v_143 | 1'h0;
  assign v_143 = ~v_130;
  assign v_144 = mux_144(v_145);
  assign v_145 = ~v_140;
  pebbles_core
    pebbles_core_146
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_147),
       .in0_consume_en(vin0_consume_en_146),
       .out_canPeek(vout_canPeek_146),
       .out_peek(vout_peek_146));
  assign v_147 = v_148 | v_149;
  assign v_148 = mux_148(v_134);
  assign v_149 = mux_149(v_150);
  assign v_150 = ~v_134;
  assign v_151 = v_152 & 1'h1;
  assign v_152 = v_153 & v_154;
  assign v_153 = ~act_133;
  assign v_154 = v_155 | v_159;
  assign v_155 = v_156 | v_157;
  assign v_156 = mux_156(v_90);
  assign v_157 = mux_157(v_158);
  assign v_158 = ~v_90;
  assign v_159 = ~v_130;
  assign v_160 = v_161 | v_162;
  assign v_161 = mux_161(v_132);
  assign v_162 = mux_162(v_151);
  assign v_163 = v_164 & 1'h1;
  assign v_164 = v_165 & v_166;
  assign v_165 = ~act_89;
  assign v_166 = v_167 | v_171;
  assign v_167 = v_168 | v_169;
  assign v_168 = mux_168(v_83);
  assign v_169 = mux_169(v_170);
  assign v_170 = ~v_83;
  assign v_171 = ~v_86;
  assign v_172 = v_173 | v_174;
  assign v_173 = mux_173(v_88);
  assign v_174 = mux_174(v_163);
  assign v_175 = v_176 & 1'h1;
  assign v_176 = v_177 & v_178;
  assign v_177 = ~act_82;
  assign v_178 = v_179 | v_22361;
  assign v_179 = v_180 | v_22359;
  assign v_180 = mux_180(v_181);
  assign v_181 = v_79 & v_182;
  assign v_182 = v_183 & 1'h1;
  assign v_183 = v_184 | 1'h0;
  assign v_184 = ~v_185;
  assign v_186 = v_187 | v_393;
  assign v_187 = act_188 & 1'h1;
  assign act_188 = v_189 | v_181;
  assign v_189 = v_190 & v_182;
  assign v_190 = v_191 & v_192;
  assign v_191 = ~v_79;
  assign v_193 = v_194 | v_381;
  assign v_194 = act_195 & 1'h1;
  assign act_195 = v_196 | v_282;
  assign v_196 = v_197 & v_283;
  assign v_197 = v_198 & v_292;
  assign v_198 = ~v_199;
  assign v_200 = v_201 | v_276;
  assign v_201 = act_202 & 1'h1;
  assign act_202 = v_203 | v_233;
  assign v_203 = v_204 & v_234;
  assign v_204 = v_205 & v_243;
  assign v_205 = ~v_206;
  assign v_207 = v_208 | v_227;
  assign v_208 = act_209 & 1'h1;
  assign act_209 = v_210 | v_216;
  assign v_210 = v_211 & v_217;
  assign v_211 = v_212 & vout_canPeek_222;
  assign v_212 = ~vout_canPeek_213;
  pebbles_core
    pebbles_core_213
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_214),
       .in0_consume_en(vin0_consume_en_213),
       .out_canPeek(vout_canPeek_213),
       .out_peek(vout_peek_213));
  assign v_214 = v_215 | v_220;
  assign v_215 = mux_215(v_216);
  assign v_216 = vout_canPeek_213 & v_217;
  assign v_217 = v_218 & 1'h1;
  assign v_218 = v_219 | 1'h0;
  assign v_219 = ~v_206;
  assign v_220 = mux_220(v_221);
  assign v_221 = ~v_216;
  pebbles_core
    pebbles_core_222
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_223),
       .in0_consume_en(vin0_consume_en_222),
       .out_canPeek(vout_canPeek_222),
       .out_peek(vout_peek_222));
  assign v_223 = v_224 | v_225;
  assign v_224 = mux_224(v_210);
  assign v_225 = mux_225(v_226);
  assign v_226 = ~v_210;
  assign v_227 = v_228 & 1'h1;
  assign v_228 = v_229 & v_230;
  assign v_229 = ~act_209;
  assign v_230 = v_231 | v_239;
  assign v_231 = v_232 | v_237;
  assign v_232 = mux_232(v_233);
  assign v_233 = v_206 & v_234;
  assign v_234 = v_235 & 1'h1;
  assign v_235 = v_236 | 1'h0;
  assign v_236 = ~v_199;
  assign v_237 = mux_237(v_238);
  assign v_238 = ~v_233;
  assign v_239 = ~v_206;
  assign v_240 = v_241 | v_242;
  assign v_241 = mux_241(v_208);
  assign v_242 = mux_242(v_227);
  assign v_244 = v_245 | v_264;
  assign v_245 = act_246 & 1'h1;
  assign act_246 = v_247 | v_253;
  assign v_247 = v_248 & v_254;
  assign v_248 = v_249 & vout_canPeek_259;
  assign v_249 = ~vout_canPeek_250;
  pebbles_core
    pebbles_core_250
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_251),
       .in0_consume_en(vin0_consume_en_250),
       .out_canPeek(vout_canPeek_250),
       .out_peek(vout_peek_250));
  assign v_251 = v_252 | v_257;
  assign v_252 = mux_252(v_253);
  assign v_253 = vout_canPeek_250 & v_254;
  assign v_254 = v_255 & 1'h1;
  assign v_255 = v_256 | 1'h0;
  assign v_256 = ~v_243;
  assign v_257 = mux_257(v_258);
  assign v_258 = ~v_253;
  pebbles_core
    pebbles_core_259
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_260),
       .in0_consume_en(vin0_consume_en_259),
       .out_canPeek(vout_canPeek_259),
       .out_peek(vout_peek_259));
  assign v_260 = v_261 | v_262;
  assign v_261 = mux_261(v_247);
  assign v_262 = mux_262(v_263);
  assign v_263 = ~v_247;
  assign v_264 = v_265 & 1'h1;
  assign v_265 = v_266 & v_267;
  assign v_266 = ~act_246;
  assign v_267 = v_268 | v_272;
  assign v_268 = v_269 | v_270;
  assign v_269 = mux_269(v_203);
  assign v_270 = mux_270(v_271);
  assign v_271 = ~v_203;
  assign v_272 = ~v_243;
  assign v_273 = v_274 | v_275;
  assign v_274 = mux_274(v_245);
  assign v_275 = mux_275(v_264);
  assign v_276 = v_277 & 1'h1;
  assign v_277 = v_278 & v_279;
  assign v_278 = ~act_202;
  assign v_279 = v_280 | v_288;
  assign v_280 = v_281 | v_286;
  assign v_281 = mux_281(v_282);
  assign v_282 = v_199 & v_283;
  assign v_283 = v_284 & 1'h1;
  assign v_284 = v_285 | 1'h0;
  assign v_285 = ~v_192;
  assign v_286 = mux_286(v_287);
  assign v_287 = ~v_282;
  assign v_288 = ~v_199;
  assign v_289 = v_290 | v_291;
  assign v_290 = mux_290(v_201);
  assign v_291 = mux_291(v_276);
  assign v_293 = v_294 | v_369;
  assign v_294 = act_295 & 1'h1;
  assign act_295 = v_296 | v_326;
  assign v_296 = v_297 & v_327;
  assign v_297 = v_298 & v_336;
  assign v_298 = ~v_299;
  assign v_300 = v_301 | v_320;
  assign v_301 = act_302 & 1'h1;
  assign act_302 = v_303 | v_309;
  assign v_303 = v_304 & v_310;
  assign v_304 = v_305 & vout_canPeek_315;
  assign v_305 = ~vout_canPeek_306;
  pebbles_core
    pebbles_core_306
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_307),
       .in0_consume_en(vin0_consume_en_306),
       .out_canPeek(vout_canPeek_306),
       .out_peek(vout_peek_306));
  assign v_307 = v_308 | v_313;
  assign v_308 = mux_308(v_309);
  assign v_309 = vout_canPeek_306 & v_310;
  assign v_310 = v_311 & 1'h1;
  assign v_311 = v_312 | 1'h0;
  assign v_312 = ~v_299;
  assign v_313 = mux_313(v_314);
  assign v_314 = ~v_309;
  pebbles_core
    pebbles_core_315
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_316),
       .in0_consume_en(vin0_consume_en_315),
       .out_canPeek(vout_canPeek_315),
       .out_peek(vout_peek_315));
  assign v_316 = v_317 | v_318;
  assign v_317 = mux_317(v_303);
  assign v_318 = mux_318(v_319);
  assign v_319 = ~v_303;
  assign v_320 = v_321 & 1'h1;
  assign v_321 = v_322 & v_323;
  assign v_322 = ~act_302;
  assign v_323 = v_324 | v_332;
  assign v_324 = v_325 | v_330;
  assign v_325 = mux_325(v_326);
  assign v_326 = v_299 & v_327;
  assign v_327 = v_328 & 1'h1;
  assign v_328 = v_329 | 1'h0;
  assign v_329 = ~v_292;
  assign v_330 = mux_330(v_331);
  assign v_331 = ~v_326;
  assign v_332 = ~v_299;
  assign v_333 = v_334 | v_335;
  assign v_334 = mux_334(v_301);
  assign v_335 = mux_335(v_320);
  assign v_337 = v_338 | v_357;
  assign v_338 = act_339 & 1'h1;
  assign act_339 = v_340 | v_346;
  assign v_340 = v_341 & v_347;
  assign v_341 = v_342 & vout_canPeek_352;
  assign v_342 = ~vout_canPeek_343;
  pebbles_core
    pebbles_core_343
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_344),
       .in0_consume_en(vin0_consume_en_343),
       .out_canPeek(vout_canPeek_343),
       .out_peek(vout_peek_343));
  assign v_344 = v_345 | v_350;
  assign v_345 = mux_345(v_346);
  assign v_346 = vout_canPeek_343 & v_347;
  assign v_347 = v_348 & 1'h1;
  assign v_348 = v_349 | 1'h0;
  assign v_349 = ~v_336;
  assign v_350 = mux_350(v_351);
  assign v_351 = ~v_346;
  pebbles_core
    pebbles_core_352
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_353),
       .in0_consume_en(vin0_consume_en_352),
       .out_canPeek(vout_canPeek_352),
       .out_peek(vout_peek_352));
  assign v_353 = v_354 | v_355;
  assign v_354 = mux_354(v_340);
  assign v_355 = mux_355(v_356);
  assign v_356 = ~v_340;
  assign v_357 = v_358 & 1'h1;
  assign v_358 = v_359 & v_360;
  assign v_359 = ~act_339;
  assign v_360 = v_361 | v_365;
  assign v_361 = v_362 | v_363;
  assign v_362 = mux_362(v_296);
  assign v_363 = mux_363(v_364);
  assign v_364 = ~v_296;
  assign v_365 = ~v_336;
  assign v_366 = v_367 | v_368;
  assign v_367 = mux_367(v_338);
  assign v_368 = mux_368(v_357);
  assign v_369 = v_370 & 1'h1;
  assign v_370 = v_371 & v_372;
  assign v_371 = ~act_295;
  assign v_372 = v_373 | v_377;
  assign v_373 = v_374 | v_375;
  assign v_374 = mux_374(v_196);
  assign v_375 = mux_375(v_376);
  assign v_376 = ~v_196;
  assign v_377 = ~v_292;
  assign v_378 = v_379 | v_380;
  assign v_379 = mux_379(v_294);
  assign v_380 = mux_380(v_369);
  assign v_381 = v_382 & 1'h1;
  assign v_382 = v_383 & v_384;
  assign v_383 = ~act_195;
  assign v_384 = v_385 | v_389;
  assign v_385 = v_386 | v_387;
  assign v_386 = mux_386(v_189);
  assign v_387 = mux_387(v_388);
  assign v_388 = ~v_189;
  assign v_389 = ~v_192;
  assign v_390 = v_391 | v_392;
  assign v_391 = mux_391(v_194);
  assign v_392 = mux_392(v_381);
  assign v_393 = v_394 & 1'h1;
  assign v_394 = v_395 & v_396;
  assign v_395 = ~act_188;
  assign v_396 = v_397 | v_22355;
  assign v_397 = v_398 | v_22353;
  assign v_398 = mux_398(v_399);
  assign v_399 = v_185 & v_400;
  assign v_400 = v_401 & 1'h1;
  assign v_401 = v_402 | 1'h0;
  assign v_402 = ~v_403;
  assign v_404 = v_405 | v_835;
  assign v_405 = act_406 & 1'h1;
  assign act_406 = v_407 | v_399;
  assign v_407 = v_408 & v_400;
  assign v_408 = v_409 & v_410;
  assign v_409 = ~v_185;
  assign v_411 = v_412 | v_823;
  assign v_412 = act_413 & 1'h1;
  assign act_413 = v_414 | v_612;
  assign v_414 = v_415 & v_613;
  assign v_415 = v_416 & v_622;
  assign v_416 = ~v_417;
  assign v_418 = v_419 | v_606;
  assign v_419 = act_420 & 1'h1;
  assign act_420 = v_421 | v_507;
  assign v_421 = v_422 & v_508;
  assign v_422 = v_423 & v_517;
  assign v_423 = ~v_424;
  assign v_425 = v_426 | v_501;
  assign v_426 = act_427 & 1'h1;
  assign act_427 = v_428 | v_458;
  assign v_428 = v_429 & v_459;
  assign v_429 = v_430 & v_468;
  assign v_430 = ~v_431;
  assign v_432 = v_433 | v_452;
  assign v_433 = act_434 & 1'h1;
  assign act_434 = v_435 | v_441;
  assign v_435 = v_436 & v_442;
  assign v_436 = v_437 & vout_canPeek_447;
  assign v_437 = ~vout_canPeek_438;
  pebbles_core
    pebbles_core_438
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_439),
       .in0_consume_en(vin0_consume_en_438),
       .out_canPeek(vout_canPeek_438),
       .out_peek(vout_peek_438));
  assign v_439 = v_440 | v_445;
  assign v_440 = mux_440(v_441);
  assign v_441 = vout_canPeek_438 & v_442;
  assign v_442 = v_443 & 1'h1;
  assign v_443 = v_444 | 1'h0;
  assign v_444 = ~v_431;
  assign v_445 = mux_445(v_446);
  assign v_446 = ~v_441;
  pebbles_core
    pebbles_core_447
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_448),
       .in0_consume_en(vin0_consume_en_447),
       .out_canPeek(vout_canPeek_447),
       .out_peek(vout_peek_447));
  assign v_448 = v_449 | v_450;
  assign v_449 = mux_449(v_435);
  assign v_450 = mux_450(v_451);
  assign v_451 = ~v_435;
  assign v_452 = v_453 & 1'h1;
  assign v_453 = v_454 & v_455;
  assign v_454 = ~act_434;
  assign v_455 = v_456 | v_464;
  assign v_456 = v_457 | v_462;
  assign v_457 = mux_457(v_458);
  assign v_458 = v_431 & v_459;
  assign v_459 = v_460 & 1'h1;
  assign v_460 = v_461 | 1'h0;
  assign v_461 = ~v_424;
  assign v_462 = mux_462(v_463);
  assign v_463 = ~v_458;
  assign v_464 = ~v_431;
  assign v_465 = v_466 | v_467;
  assign v_466 = mux_466(v_433);
  assign v_467 = mux_467(v_452);
  assign v_469 = v_470 | v_489;
  assign v_470 = act_471 & 1'h1;
  assign act_471 = v_472 | v_478;
  assign v_472 = v_473 & v_479;
  assign v_473 = v_474 & vout_canPeek_484;
  assign v_474 = ~vout_canPeek_475;
  pebbles_core
    pebbles_core_475
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_476),
       .in0_consume_en(vin0_consume_en_475),
       .out_canPeek(vout_canPeek_475),
       .out_peek(vout_peek_475));
  assign v_476 = v_477 | v_482;
  assign v_477 = mux_477(v_478);
  assign v_478 = vout_canPeek_475 & v_479;
  assign v_479 = v_480 & 1'h1;
  assign v_480 = v_481 | 1'h0;
  assign v_481 = ~v_468;
  assign v_482 = mux_482(v_483);
  assign v_483 = ~v_478;
  pebbles_core
    pebbles_core_484
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_485),
       .in0_consume_en(vin0_consume_en_484),
       .out_canPeek(vout_canPeek_484),
       .out_peek(vout_peek_484));
  assign v_485 = v_486 | v_487;
  assign v_486 = mux_486(v_472);
  assign v_487 = mux_487(v_488);
  assign v_488 = ~v_472;
  assign v_489 = v_490 & 1'h1;
  assign v_490 = v_491 & v_492;
  assign v_491 = ~act_471;
  assign v_492 = v_493 | v_497;
  assign v_493 = v_494 | v_495;
  assign v_494 = mux_494(v_428);
  assign v_495 = mux_495(v_496);
  assign v_496 = ~v_428;
  assign v_497 = ~v_468;
  assign v_498 = v_499 | v_500;
  assign v_499 = mux_499(v_470);
  assign v_500 = mux_500(v_489);
  assign v_501 = v_502 & 1'h1;
  assign v_502 = v_503 & v_504;
  assign v_503 = ~act_427;
  assign v_504 = v_505 | v_513;
  assign v_505 = v_506 | v_511;
  assign v_506 = mux_506(v_507);
  assign v_507 = v_424 & v_508;
  assign v_508 = v_509 & 1'h1;
  assign v_509 = v_510 | 1'h0;
  assign v_510 = ~v_417;
  assign v_511 = mux_511(v_512);
  assign v_512 = ~v_507;
  assign v_513 = ~v_424;
  assign v_514 = v_515 | v_516;
  assign v_515 = mux_515(v_426);
  assign v_516 = mux_516(v_501);
  assign v_518 = v_519 | v_594;
  assign v_519 = act_520 & 1'h1;
  assign act_520 = v_521 | v_551;
  assign v_521 = v_522 & v_552;
  assign v_522 = v_523 & v_561;
  assign v_523 = ~v_524;
  assign v_525 = v_526 | v_545;
  assign v_526 = act_527 & 1'h1;
  assign act_527 = v_528 | v_534;
  assign v_528 = v_529 & v_535;
  assign v_529 = v_530 & vout_canPeek_540;
  assign v_530 = ~vout_canPeek_531;
  pebbles_core
    pebbles_core_531
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_532),
       .in0_consume_en(vin0_consume_en_531),
       .out_canPeek(vout_canPeek_531),
       .out_peek(vout_peek_531));
  assign v_532 = v_533 | v_538;
  assign v_533 = mux_533(v_534);
  assign v_534 = vout_canPeek_531 & v_535;
  assign v_535 = v_536 & 1'h1;
  assign v_536 = v_537 | 1'h0;
  assign v_537 = ~v_524;
  assign v_538 = mux_538(v_539);
  assign v_539 = ~v_534;
  pebbles_core
    pebbles_core_540
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_541),
       .in0_consume_en(vin0_consume_en_540),
       .out_canPeek(vout_canPeek_540),
       .out_peek(vout_peek_540));
  assign v_541 = v_542 | v_543;
  assign v_542 = mux_542(v_528);
  assign v_543 = mux_543(v_544);
  assign v_544 = ~v_528;
  assign v_545 = v_546 & 1'h1;
  assign v_546 = v_547 & v_548;
  assign v_547 = ~act_527;
  assign v_548 = v_549 | v_557;
  assign v_549 = v_550 | v_555;
  assign v_550 = mux_550(v_551);
  assign v_551 = v_524 & v_552;
  assign v_552 = v_553 & 1'h1;
  assign v_553 = v_554 | 1'h0;
  assign v_554 = ~v_517;
  assign v_555 = mux_555(v_556);
  assign v_556 = ~v_551;
  assign v_557 = ~v_524;
  assign v_558 = v_559 | v_560;
  assign v_559 = mux_559(v_526);
  assign v_560 = mux_560(v_545);
  assign v_562 = v_563 | v_582;
  assign v_563 = act_564 & 1'h1;
  assign act_564 = v_565 | v_571;
  assign v_565 = v_566 & v_572;
  assign v_566 = v_567 & vout_canPeek_577;
  assign v_567 = ~vout_canPeek_568;
  pebbles_core
    pebbles_core_568
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_569),
       .in0_consume_en(vin0_consume_en_568),
       .out_canPeek(vout_canPeek_568),
       .out_peek(vout_peek_568));
  assign v_569 = v_570 | v_575;
  assign v_570 = mux_570(v_571);
  assign v_571 = vout_canPeek_568 & v_572;
  assign v_572 = v_573 & 1'h1;
  assign v_573 = v_574 | 1'h0;
  assign v_574 = ~v_561;
  assign v_575 = mux_575(v_576);
  assign v_576 = ~v_571;
  pebbles_core
    pebbles_core_577
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_578),
       .in0_consume_en(vin0_consume_en_577),
       .out_canPeek(vout_canPeek_577),
       .out_peek(vout_peek_577));
  assign v_578 = v_579 | v_580;
  assign v_579 = mux_579(v_565);
  assign v_580 = mux_580(v_581);
  assign v_581 = ~v_565;
  assign v_582 = v_583 & 1'h1;
  assign v_583 = v_584 & v_585;
  assign v_584 = ~act_564;
  assign v_585 = v_586 | v_590;
  assign v_586 = v_587 | v_588;
  assign v_587 = mux_587(v_521);
  assign v_588 = mux_588(v_589);
  assign v_589 = ~v_521;
  assign v_590 = ~v_561;
  assign v_591 = v_592 | v_593;
  assign v_592 = mux_592(v_563);
  assign v_593 = mux_593(v_582);
  assign v_594 = v_595 & 1'h1;
  assign v_595 = v_596 & v_597;
  assign v_596 = ~act_520;
  assign v_597 = v_598 | v_602;
  assign v_598 = v_599 | v_600;
  assign v_599 = mux_599(v_421);
  assign v_600 = mux_600(v_601);
  assign v_601 = ~v_421;
  assign v_602 = ~v_517;
  assign v_603 = v_604 | v_605;
  assign v_604 = mux_604(v_519);
  assign v_605 = mux_605(v_594);
  assign v_606 = v_607 & 1'h1;
  assign v_607 = v_608 & v_609;
  assign v_608 = ~act_420;
  assign v_609 = v_610 | v_618;
  assign v_610 = v_611 | v_616;
  assign v_611 = mux_611(v_612);
  assign v_612 = v_417 & v_613;
  assign v_613 = v_614 & 1'h1;
  assign v_614 = v_615 | 1'h0;
  assign v_615 = ~v_410;
  assign v_616 = mux_616(v_617);
  assign v_617 = ~v_612;
  assign v_618 = ~v_417;
  assign v_619 = v_620 | v_621;
  assign v_620 = mux_620(v_419);
  assign v_621 = mux_621(v_606);
  assign v_623 = v_624 | v_811;
  assign v_624 = act_625 & 1'h1;
  assign act_625 = v_626 | v_712;
  assign v_626 = v_627 & v_713;
  assign v_627 = v_628 & v_722;
  assign v_628 = ~v_629;
  assign v_630 = v_631 | v_706;
  assign v_631 = act_632 & 1'h1;
  assign act_632 = v_633 | v_663;
  assign v_633 = v_634 & v_664;
  assign v_634 = v_635 & v_673;
  assign v_635 = ~v_636;
  assign v_637 = v_638 | v_657;
  assign v_638 = act_639 & 1'h1;
  assign act_639 = v_640 | v_646;
  assign v_640 = v_641 & v_647;
  assign v_641 = v_642 & vout_canPeek_652;
  assign v_642 = ~vout_canPeek_643;
  pebbles_core
    pebbles_core_643
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_644),
       .in0_consume_en(vin0_consume_en_643),
       .out_canPeek(vout_canPeek_643),
       .out_peek(vout_peek_643));
  assign v_644 = v_645 | v_650;
  assign v_645 = mux_645(v_646);
  assign v_646 = vout_canPeek_643 & v_647;
  assign v_647 = v_648 & 1'h1;
  assign v_648 = v_649 | 1'h0;
  assign v_649 = ~v_636;
  assign v_650 = mux_650(v_651);
  assign v_651 = ~v_646;
  pebbles_core
    pebbles_core_652
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_653),
       .in0_consume_en(vin0_consume_en_652),
       .out_canPeek(vout_canPeek_652),
       .out_peek(vout_peek_652));
  assign v_653 = v_654 | v_655;
  assign v_654 = mux_654(v_640);
  assign v_655 = mux_655(v_656);
  assign v_656 = ~v_640;
  assign v_657 = v_658 & 1'h1;
  assign v_658 = v_659 & v_660;
  assign v_659 = ~act_639;
  assign v_660 = v_661 | v_669;
  assign v_661 = v_662 | v_667;
  assign v_662 = mux_662(v_663);
  assign v_663 = v_636 & v_664;
  assign v_664 = v_665 & 1'h1;
  assign v_665 = v_666 | 1'h0;
  assign v_666 = ~v_629;
  assign v_667 = mux_667(v_668);
  assign v_668 = ~v_663;
  assign v_669 = ~v_636;
  assign v_670 = v_671 | v_672;
  assign v_671 = mux_671(v_638);
  assign v_672 = mux_672(v_657);
  assign v_674 = v_675 | v_694;
  assign v_675 = act_676 & 1'h1;
  assign act_676 = v_677 | v_683;
  assign v_677 = v_678 & v_684;
  assign v_678 = v_679 & vout_canPeek_689;
  assign v_679 = ~vout_canPeek_680;
  pebbles_core
    pebbles_core_680
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_681),
       .in0_consume_en(vin0_consume_en_680),
       .out_canPeek(vout_canPeek_680),
       .out_peek(vout_peek_680));
  assign v_681 = v_682 | v_687;
  assign v_682 = mux_682(v_683);
  assign v_683 = vout_canPeek_680 & v_684;
  assign v_684 = v_685 & 1'h1;
  assign v_685 = v_686 | 1'h0;
  assign v_686 = ~v_673;
  assign v_687 = mux_687(v_688);
  assign v_688 = ~v_683;
  pebbles_core
    pebbles_core_689
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_690),
       .in0_consume_en(vin0_consume_en_689),
       .out_canPeek(vout_canPeek_689),
       .out_peek(vout_peek_689));
  assign v_690 = v_691 | v_692;
  assign v_691 = mux_691(v_677);
  assign v_692 = mux_692(v_693);
  assign v_693 = ~v_677;
  assign v_694 = v_695 & 1'h1;
  assign v_695 = v_696 & v_697;
  assign v_696 = ~act_676;
  assign v_697 = v_698 | v_702;
  assign v_698 = v_699 | v_700;
  assign v_699 = mux_699(v_633);
  assign v_700 = mux_700(v_701);
  assign v_701 = ~v_633;
  assign v_702 = ~v_673;
  assign v_703 = v_704 | v_705;
  assign v_704 = mux_704(v_675);
  assign v_705 = mux_705(v_694);
  assign v_706 = v_707 & 1'h1;
  assign v_707 = v_708 & v_709;
  assign v_708 = ~act_632;
  assign v_709 = v_710 | v_718;
  assign v_710 = v_711 | v_716;
  assign v_711 = mux_711(v_712);
  assign v_712 = v_629 & v_713;
  assign v_713 = v_714 & 1'h1;
  assign v_714 = v_715 | 1'h0;
  assign v_715 = ~v_622;
  assign v_716 = mux_716(v_717);
  assign v_717 = ~v_712;
  assign v_718 = ~v_629;
  assign v_719 = v_720 | v_721;
  assign v_720 = mux_720(v_631);
  assign v_721 = mux_721(v_706);
  assign v_723 = v_724 | v_799;
  assign v_724 = act_725 & 1'h1;
  assign act_725 = v_726 | v_756;
  assign v_726 = v_727 & v_757;
  assign v_727 = v_728 & v_766;
  assign v_728 = ~v_729;
  assign v_730 = v_731 | v_750;
  assign v_731 = act_732 & 1'h1;
  assign act_732 = v_733 | v_739;
  assign v_733 = v_734 & v_740;
  assign v_734 = v_735 & vout_canPeek_745;
  assign v_735 = ~vout_canPeek_736;
  pebbles_core
    pebbles_core_736
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_737),
       .in0_consume_en(vin0_consume_en_736),
       .out_canPeek(vout_canPeek_736),
       .out_peek(vout_peek_736));
  assign v_737 = v_738 | v_743;
  assign v_738 = mux_738(v_739);
  assign v_739 = vout_canPeek_736 & v_740;
  assign v_740 = v_741 & 1'h1;
  assign v_741 = v_742 | 1'h0;
  assign v_742 = ~v_729;
  assign v_743 = mux_743(v_744);
  assign v_744 = ~v_739;
  pebbles_core
    pebbles_core_745
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_746),
       .in0_consume_en(vin0_consume_en_745),
       .out_canPeek(vout_canPeek_745),
       .out_peek(vout_peek_745));
  assign v_746 = v_747 | v_748;
  assign v_747 = mux_747(v_733);
  assign v_748 = mux_748(v_749);
  assign v_749 = ~v_733;
  assign v_750 = v_751 & 1'h1;
  assign v_751 = v_752 & v_753;
  assign v_752 = ~act_732;
  assign v_753 = v_754 | v_762;
  assign v_754 = v_755 | v_760;
  assign v_755 = mux_755(v_756);
  assign v_756 = v_729 & v_757;
  assign v_757 = v_758 & 1'h1;
  assign v_758 = v_759 | 1'h0;
  assign v_759 = ~v_722;
  assign v_760 = mux_760(v_761);
  assign v_761 = ~v_756;
  assign v_762 = ~v_729;
  assign v_763 = v_764 | v_765;
  assign v_764 = mux_764(v_731);
  assign v_765 = mux_765(v_750);
  assign v_767 = v_768 | v_787;
  assign v_768 = act_769 & 1'h1;
  assign act_769 = v_770 | v_776;
  assign v_770 = v_771 & v_777;
  assign v_771 = v_772 & vout_canPeek_782;
  assign v_772 = ~vout_canPeek_773;
  pebbles_core
    pebbles_core_773
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_774),
       .in0_consume_en(vin0_consume_en_773),
       .out_canPeek(vout_canPeek_773),
       .out_peek(vout_peek_773));
  assign v_774 = v_775 | v_780;
  assign v_775 = mux_775(v_776);
  assign v_776 = vout_canPeek_773 & v_777;
  assign v_777 = v_778 & 1'h1;
  assign v_778 = v_779 | 1'h0;
  assign v_779 = ~v_766;
  assign v_780 = mux_780(v_781);
  assign v_781 = ~v_776;
  pebbles_core
    pebbles_core_782
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_783),
       .in0_consume_en(vin0_consume_en_782),
       .out_canPeek(vout_canPeek_782),
       .out_peek(vout_peek_782));
  assign v_783 = v_784 | v_785;
  assign v_784 = mux_784(v_770);
  assign v_785 = mux_785(v_786);
  assign v_786 = ~v_770;
  assign v_787 = v_788 & 1'h1;
  assign v_788 = v_789 & v_790;
  assign v_789 = ~act_769;
  assign v_790 = v_791 | v_795;
  assign v_791 = v_792 | v_793;
  assign v_792 = mux_792(v_726);
  assign v_793 = mux_793(v_794);
  assign v_794 = ~v_726;
  assign v_795 = ~v_766;
  assign v_796 = v_797 | v_798;
  assign v_797 = mux_797(v_768);
  assign v_798 = mux_798(v_787);
  assign v_799 = v_800 & 1'h1;
  assign v_800 = v_801 & v_802;
  assign v_801 = ~act_725;
  assign v_802 = v_803 | v_807;
  assign v_803 = v_804 | v_805;
  assign v_804 = mux_804(v_626);
  assign v_805 = mux_805(v_806);
  assign v_806 = ~v_626;
  assign v_807 = ~v_722;
  assign v_808 = v_809 | v_810;
  assign v_809 = mux_809(v_724);
  assign v_810 = mux_810(v_799);
  assign v_811 = v_812 & 1'h1;
  assign v_812 = v_813 & v_814;
  assign v_813 = ~act_625;
  assign v_814 = v_815 | v_819;
  assign v_815 = v_816 | v_817;
  assign v_816 = mux_816(v_414);
  assign v_817 = mux_817(v_818);
  assign v_818 = ~v_414;
  assign v_819 = ~v_622;
  assign v_820 = v_821 | v_822;
  assign v_821 = mux_821(v_624);
  assign v_822 = mux_822(v_811);
  assign v_823 = v_824 & 1'h1;
  assign v_824 = v_825 & v_826;
  assign v_825 = ~act_413;
  assign v_826 = v_827 | v_831;
  assign v_827 = v_828 | v_829;
  assign v_828 = mux_828(v_407);
  assign v_829 = mux_829(v_830);
  assign v_830 = ~v_407;
  assign v_831 = ~v_410;
  assign v_832 = v_833 | v_834;
  assign v_833 = mux_833(v_412);
  assign v_834 = mux_834(v_823);
  assign v_835 = v_836 & 1'h1;
  assign v_836 = v_837 & v_838;
  assign v_837 = ~act_406;
  assign v_838 = v_839 | v_22349;
  assign v_839 = v_840 | v_22347;
  assign v_840 = mux_840(v_841);
  assign v_841 = v_403 & v_842;
  assign v_842 = v_843 & 1'h1;
  assign v_843 = v_844 | 1'h0;
  assign v_844 = ~v_845;
  assign v_846 = v_847 | v_1725;
  assign v_847 = act_848 & 1'h1;
  assign act_848 = v_849 | v_841;
  assign v_849 = v_850 & v_842;
  assign v_850 = v_851 & v_852;
  assign v_851 = ~v_403;
  assign v_853 = v_854 | v_1713;
  assign v_854 = act_855 & 1'h1;
  assign act_855 = v_856 | v_1278;
  assign v_856 = v_857 & v_1279;
  assign v_857 = v_858 & v_1288;
  assign v_858 = ~v_859;
  assign v_860 = v_861 | v_1272;
  assign v_861 = act_862 & 1'h1;
  assign act_862 = v_863 | v_1061;
  assign v_863 = v_864 & v_1062;
  assign v_864 = v_865 & v_1071;
  assign v_865 = ~v_866;
  assign v_867 = v_868 | v_1055;
  assign v_868 = act_869 & 1'h1;
  assign act_869 = v_870 | v_956;
  assign v_870 = v_871 & v_957;
  assign v_871 = v_872 & v_966;
  assign v_872 = ~v_873;
  assign v_874 = v_875 | v_950;
  assign v_875 = act_876 & 1'h1;
  assign act_876 = v_877 | v_907;
  assign v_877 = v_878 & v_908;
  assign v_878 = v_879 & v_917;
  assign v_879 = ~v_880;
  assign v_881 = v_882 | v_901;
  assign v_882 = act_883 & 1'h1;
  assign act_883 = v_884 | v_890;
  assign v_884 = v_885 & v_891;
  assign v_885 = v_886 & vout_canPeek_896;
  assign v_886 = ~vout_canPeek_887;
  pebbles_core
    pebbles_core_887
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_888),
       .in0_consume_en(vin0_consume_en_887),
       .out_canPeek(vout_canPeek_887),
       .out_peek(vout_peek_887));
  assign v_888 = v_889 | v_894;
  assign v_889 = mux_889(v_890);
  assign v_890 = vout_canPeek_887 & v_891;
  assign v_891 = v_892 & 1'h1;
  assign v_892 = v_893 | 1'h0;
  assign v_893 = ~v_880;
  assign v_894 = mux_894(v_895);
  assign v_895 = ~v_890;
  pebbles_core
    pebbles_core_896
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_897),
       .in0_consume_en(vin0_consume_en_896),
       .out_canPeek(vout_canPeek_896),
       .out_peek(vout_peek_896));
  assign v_897 = v_898 | v_899;
  assign v_898 = mux_898(v_884);
  assign v_899 = mux_899(v_900);
  assign v_900 = ~v_884;
  assign v_901 = v_902 & 1'h1;
  assign v_902 = v_903 & v_904;
  assign v_903 = ~act_883;
  assign v_904 = v_905 | v_913;
  assign v_905 = v_906 | v_911;
  assign v_906 = mux_906(v_907);
  assign v_907 = v_880 & v_908;
  assign v_908 = v_909 & 1'h1;
  assign v_909 = v_910 | 1'h0;
  assign v_910 = ~v_873;
  assign v_911 = mux_911(v_912);
  assign v_912 = ~v_907;
  assign v_913 = ~v_880;
  assign v_914 = v_915 | v_916;
  assign v_915 = mux_915(v_882);
  assign v_916 = mux_916(v_901);
  assign v_918 = v_919 | v_938;
  assign v_919 = act_920 & 1'h1;
  assign act_920 = v_921 | v_927;
  assign v_921 = v_922 & v_928;
  assign v_922 = v_923 & vout_canPeek_933;
  assign v_923 = ~vout_canPeek_924;
  pebbles_core
    pebbles_core_924
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_925),
       .in0_consume_en(vin0_consume_en_924),
       .out_canPeek(vout_canPeek_924),
       .out_peek(vout_peek_924));
  assign v_925 = v_926 | v_931;
  assign v_926 = mux_926(v_927);
  assign v_927 = vout_canPeek_924 & v_928;
  assign v_928 = v_929 & 1'h1;
  assign v_929 = v_930 | 1'h0;
  assign v_930 = ~v_917;
  assign v_931 = mux_931(v_932);
  assign v_932 = ~v_927;
  pebbles_core
    pebbles_core_933
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_934),
       .in0_consume_en(vin0_consume_en_933),
       .out_canPeek(vout_canPeek_933),
       .out_peek(vout_peek_933));
  assign v_934 = v_935 | v_936;
  assign v_935 = mux_935(v_921);
  assign v_936 = mux_936(v_937);
  assign v_937 = ~v_921;
  assign v_938 = v_939 & 1'h1;
  assign v_939 = v_940 & v_941;
  assign v_940 = ~act_920;
  assign v_941 = v_942 | v_946;
  assign v_942 = v_943 | v_944;
  assign v_943 = mux_943(v_877);
  assign v_944 = mux_944(v_945);
  assign v_945 = ~v_877;
  assign v_946 = ~v_917;
  assign v_947 = v_948 | v_949;
  assign v_948 = mux_948(v_919);
  assign v_949 = mux_949(v_938);
  assign v_950 = v_951 & 1'h1;
  assign v_951 = v_952 & v_953;
  assign v_952 = ~act_876;
  assign v_953 = v_954 | v_962;
  assign v_954 = v_955 | v_960;
  assign v_955 = mux_955(v_956);
  assign v_956 = v_873 & v_957;
  assign v_957 = v_958 & 1'h1;
  assign v_958 = v_959 | 1'h0;
  assign v_959 = ~v_866;
  assign v_960 = mux_960(v_961);
  assign v_961 = ~v_956;
  assign v_962 = ~v_873;
  assign v_963 = v_964 | v_965;
  assign v_964 = mux_964(v_875);
  assign v_965 = mux_965(v_950);
  assign v_967 = v_968 | v_1043;
  assign v_968 = act_969 & 1'h1;
  assign act_969 = v_970 | v_1000;
  assign v_970 = v_971 & v_1001;
  assign v_971 = v_972 & v_1010;
  assign v_972 = ~v_973;
  assign v_974 = v_975 | v_994;
  assign v_975 = act_976 & 1'h1;
  assign act_976 = v_977 | v_983;
  assign v_977 = v_978 & v_984;
  assign v_978 = v_979 & vout_canPeek_989;
  assign v_979 = ~vout_canPeek_980;
  pebbles_core
    pebbles_core_980
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_981),
       .in0_consume_en(vin0_consume_en_980),
       .out_canPeek(vout_canPeek_980),
       .out_peek(vout_peek_980));
  assign v_981 = v_982 | v_987;
  assign v_982 = mux_982(v_983);
  assign v_983 = vout_canPeek_980 & v_984;
  assign v_984 = v_985 & 1'h1;
  assign v_985 = v_986 | 1'h0;
  assign v_986 = ~v_973;
  assign v_987 = mux_987(v_988);
  assign v_988 = ~v_983;
  pebbles_core
    pebbles_core_989
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_990),
       .in0_consume_en(vin0_consume_en_989),
       .out_canPeek(vout_canPeek_989),
       .out_peek(vout_peek_989));
  assign v_990 = v_991 | v_992;
  assign v_991 = mux_991(v_977);
  assign v_992 = mux_992(v_993);
  assign v_993 = ~v_977;
  assign v_994 = v_995 & 1'h1;
  assign v_995 = v_996 & v_997;
  assign v_996 = ~act_976;
  assign v_997 = v_998 | v_1006;
  assign v_998 = v_999 | v_1004;
  assign v_999 = mux_999(v_1000);
  assign v_1000 = v_973 & v_1001;
  assign v_1001 = v_1002 & 1'h1;
  assign v_1002 = v_1003 | 1'h0;
  assign v_1003 = ~v_966;
  assign v_1004 = mux_1004(v_1005);
  assign v_1005 = ~v_1000;
  assign v_1006 = ~v_973;
  assign v_1007 = v_1008 | v_1009;
  assign v_1008 = mux_1008(v_975);
  assign v_1009 = mux_1009(v_994);
  assign v_1011 = v_1012 | v_1031;
  assign v_1012 = act_1013 & 1'h1;
  assign act_1013 = v_1014 | v_1020;
  assign v_1014 = v_1015 & v_1021;
  assign v_1015 = v_1016 & vout_canPeek_1026;
  assign v_1016 = ~vout_canPeek_1017;
  pebbles_core
    pebbles_core_1017
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1018),
       .in0_consume_en(vin0_consume_en_1017),
       .out_canPeek(vout_canPeek_1017),
       .out_peek(vout_peek_1017));
  assign v_1018 = v_1019 | v_1024;
  assign v_1019 = mux_1019(v_1020);
  assign v_1020 = vout_canPeek_1017 & v_1021;
  assign v_1021 = v_1022 & 1'h1;
  assign v_1022 = v_1023 | 1'h0;
  assign v_1023 = ~v_1010;
  assign v_1024 = mux_1024(v_1025);
  assign v_1025 = ~v_1020;
  pebbles_core
    pebbles_core_1026
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1027),
       .in0_consume_en(vin0_consume_en_1026),
       .out_canPeek(vout_canPeek_1026),
       .out_peek(vout_peek_1026));
  assign v_1027 = v_1028 | v_1029;
  assign v_1028 = mux_1028(v_1014);
  assign v_1029 = mux_1029(v_1030);
  assign v_1030 = ~v_1014;
  assign v_1031 = v_1032 & 1'h1;
  assign v_1032 = v_1033 & v_1034;
  assign v_1033 = ~act_1013;
  assign v_1034 = v_1035 | v_1039;
  assign v_1035 = v_1036 | v_1037;
  assign v_1036 = mux_1036(v_970);
  assign v_1037 = mux_1037(v_1038);
  assign v_1038 = ~v_970;
  assign v_1039 = ~v_1010;
  assign v_1040 = v_1041 | v_1042;
  assign v_1041 = mux_1041(v_1012);
  assign v_1042 = mux_1042(v_1031);
  assign v_1043 = v_1044 & 1'h1;
  assign v_1044 = v_1045 & v_1046;
  assign v_1045 = ~act_969;
  assign v_1046 = v_1047 | v_1051;
  assign v_1047 = v_1048 | v_1049;
  assign v_1048 = mux_1048(v_870);
  assign v_1049 = mux_1049(v_1050);
  assign v_1050 = ~v_870;
  assign v_1051 = ~v_966;
  assign v_1052 = v_1053 | v_1054;
  assign v_1053 = mux_1053(v_968);
  assign v_1054 = mux_1054(v_1043);
  assign v_1055 = v_1056 & 1'h1;
  assign v_1056 = v_1057 & v_1058;
  assign v_1057 = ~act_869;
  assign v_1058 = v_1059 | v_1067;
  assign v_1059 = v_1060 | v_1065;
  assign v_1060 = mux_1060(v_1061);
  assign v_1061 = v_866 & v_1062;
  assign v_1062 = v_1063 & 1'h1;
  assign v_1063 = v_1064 | 1'h0;
  assign v_1064 = ~v_859;
  assign v_1065 = mux_1065(v_1066);
  assign v_1066 = ~v_1061;
  assign v_1067 = ~v_866;
  assign v_1068 = v_1069 | v_1070;
  assign v_1069 = mux_1069(v_868);
  assign v_1070 = mux_1070(v_1055);
  assign v_1072 = v_1073 | v_1260;
  assign v_1073 = act_1074 & 1'h1;
  assign act_1074 = v_1075 | v_1161;
  assign v_1075 = v_1076 & v_1162;
  assign v_1076 = v_1077 & v_1171;
  assign v_1077 = ~v_1078;
  assign v_1079 = v_1080 | v_1155;
  assign v_1080 = act_1081 & 1'h1;
  assign act_1081 = v_1082 | v_1112;
  assign v_1082 = v_1083 & v_1113;
  assign v_1083 = v_1084 & v_1122;
  assign v_1084 = ~v_1085;
  assign v_1086 = v_1087 | v_1106;
  assign v_1087 = act_1088 & 1'h1;
  assign act_1088 = v_1089 | v_1095;
  assign v_1089 = v_1090 & v_1096;
  assign v_1090 = v_1091 & vout_canPeek_1101;
  assign v_1091 = ~vout_canPeek_1092;
  pebbles_core
    pebbles_core_1092
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1093),
       .in0_consume_en(vin0_consume_en_1092),
       .out_canPeek(vout_canPeek_1092),
       .out_peek(vout_peek_1092));
  assign v_1093 = v_1094 | v_1099;
  assign v_1094 = mux_1094(v_1095);
  assign v_1095 = vout_canPeek_1092 & v_1096;
  assign v_1096 = v_1097 & 1'h1;
  assign v_1097 = v_1098 | 1'h0;
  assign v_1098 = ~v_1085;
  assign v_1099 = mux_1099(v_1100);
  assign v_1100 = ~v_1095;
  pebbles_core
    pebbles_core_1101
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1102),
       .in0_consume_en(vin0_consume_en_1101),
       .out_canPeek(vout_canPeek_1101),
       .out_peek(vout_peek_1101));
  assign v_1102 = v_1103 | v_1104;
  assign v_1103 = mux_1103(v_1089);
  assign v_1104 = mux_1104(v_1105);
  assign v_1105 = ~v_1089;
  assign v_1106 = v_1107 & 1'h1;
  assign v_1107 = v_1108 & v_1109;
  assign v_1108 = ~act_1088;
  assign v_1109 = v_1110 | v_1118;
  assign v_1110 = v_1111 | v_1116;
  assign v_1111 = mux_1111(v_1112);
  assign v_1112 = v_1085 & v_1113;
  assign v_1113 = v_1114 & 1'h1;
  assign v_1114 = v_1115 | 1'h0;
  assign v_1115 = ~v_1078;
  assign v_1116 = mux_1116(v_1117);
  assign v_1117 = ~v_1112;
  assign v_1118 = ~v_1085;
  assign v_1119 = v_1120 | v_1121;
  assign v_1120 = mux_1120(v_1087);
  assign v_1121 = mux_1121(v_1106);
  assign v_1123 = v_1124 | v_1143;
  assign v_1124 = act_1125 & 1'h1;
  assign act_1125 = v_1126 | v_1132;
  assign v_1126 = v_1127 & v_1133;
  assign v_1127 = v_1128 & vout_canPeek_1138;
  assign v_1128 = ~vout_canPeek_1129;
  pebbles_core
    pebbles_core_1129
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1130),
       .in0_consume_en(vin0_consume_en_1129),
       .out_canPeek(vout_canPeek_1129),
       .out_peek(vout_peek_1129));
  assign v_1130 = v_1131 | v_1136;
  assign v_1131 = mux_1131(v_1132);
  assign v_1132 = vout_canPeek_1129 & v_1133;
  assign v_1133 = v_1134 & 1'h1;
  assign v_1134 = v_1135 | 1'h0;
  assign v_1135 = ~v_1122;
  assign v_1136 = mux_1136(v_1137);
  assign v_1137 = ~v_1132;
  pebbles_core
    pebbles_core_1138
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1139),
       .in0_consume_en(vin0_consume_en_1138),
       .out_canPeek(vout_canPeek_1138),
       .out_peek(vout_peek_1138));
  assign v_1139 = v_1140 | v_1141;
  assign v_1140 = mux_1140(v_1126);
  assign v_1141 = mux_1141(v_1142);
  assign v_1142 = ~v_1126;
  assign v_1143 = v_1144 & 1'h1;
  assign v_1144 = v_1145 & v_1146;
  assign v_1145 = ~act_1125;
  assign v_1146 = v_1147 | v_1151;
  assign v_1147 = v_1148 | v_1149;
  assign v_1148 = mux_1148(v_1082);
  assign v_1149 = mux_1149(v_1150);
  assign v_1150 = ~v_1082;
  assign v_1151 = ~v_1122;
  assign v_1152 = v_1153 | v_1154;
  assign v_1153 = mux_1153(v_1124);
  assign v_1154 = mux_1154(v_1143);
  assign v_1155 = v_1156 & 1'h1;
  assign v_1156 = v_1157 & v_1158;
  assign v_1157 = ~act_1081;
  assign v_1158 = v_1159 | v_1167;
  assign v_1159 = v_1160 | v_1165;
  assign v_1160 = mux_1160(v_1161);
  assign v_1161 = v_1078 & v_1162;
  assign v_1162 = v_1163 & 1'h1;
  assign v_1163 = v_1164 | 1'h0;
  assign v_1164 = ~v_1071;
  assign v_1165 = mux_1165(v_1166);
  assign v_1166 = ~v_1161;
  assign v_1167 = ~v_1078;
  assign v_1168 = v_1169 | v_1170;
  assign v_1169 = mux_1169(v_1080);
  assign v_1170 = mux_1170(v_1155);
  assign v_1172 = v_1173 | v_1248;
  assign v_1173 = act_1174 & 1'h1;
  assign act_1174 = v_1175 | v_1205;
  assign v_1175 = v_1176 & v_1206;
  assign v_1176 = v_1177 & v_1215;
  assign v_1177 = ~v_1178;
  assign v_1179 = v_1180 | v_1199;
  assign v_1180 = act_1181 & 1'h1;
  assign act_1181 = v_1182 | v_1188;
  assign v_1182 = v_1183 & v_1189;
  assign v_1183 = v_1184 & vout_canPeek_1194;
  assign v_1184 = ~vout_canPeek_1185;
  pebbles_core
    pebbles_core_1185
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1186),
       .in0_consume_en(vin0_consume_en_1185),
       .out_canPeek(vout_canPeek_1185),
       .out_peek(vout_peek_1185));
  assign v_1186 = v_1187 | v_1192;
  assign v_1187 = mux_1187(v_1188);
  assign v_1188 = vout_canPeek_1185 & v_1189;
  assign v_1189 = v_1190 & 1'h1;
  assign v_1190 = v_1191 | 1'h0;
  assign v_1191 = ~v_1178;
  assign v_1192 = mux_1192(v_1193);
  assign v_1193 = ~v_1188;
  pebbles_core
    pebbles_core_1194
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1195),
       .in0_consume_en(vin0_consume_en_1194),
       .out_canPeek(vout_canPeek_1194),
       .out_peek(vout_peek_1194));
  assign v_1195 = v_1196 | v_1197;
  assign v_1196 = mux_1196(v_1182);
  assign v_1197 = mux_1197(v_1198);
  assign v_1198 = ~v_1182;
  assign v_1199 = v_1200 & 1'h1;
  assign v_1200 = v_1201 & v_1202;
  assign v_1201 = ~act_1181;
  assign v_1202 = v_1203 | v_1211;
  assign v_1203 = v_1204 | v_1209;
  assign v_1204 = mux_1204(v_1205);
  assign v_1205 = v_1178 & v_1206;
  assign v_1206 = v_1207 & 1'h1;
  assign v_1207 = v_1208 | 1'h0;
  assign v_1208 = ~v_1171;
  assign v_1209 = mux_1209(v_1210);
  assign v_1210 = ~v_1205;
  assign v_1211 = ~v_1178;
  assign v_1212 = v_1213 | v_1214;
  assign v_1213 = mux_1213(v_1180);
  assign v_1214 = mux_1214(v_1199);
  assign v_1216 = v_1217 | v_1236;
  assign v_1217 = act_1218 & 1'h1;
  assign act_1218 = v_1219 | v_1225;
  assign v_1219 = v_1220 & v_1226;
  assign v_1220 = v_1221 & vout_canPeek_1231;
  assign v_1221 = ~vout_canPeek_1222;
  pebbles_core
    pebbles_core_1222
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1223),
       .in0_consume_en(vin0_consume_en_1222),
       .out_canPeek(vout_canPeek_1222),
       .out_peek(vout_peek_1222));
  assign v_1223 = v_1224 | v_1229;
  assign v_1224 = mux_1224(v_1225);
  assign v_1225 = vout_canPeek_1222 & v_1226;
  assign v_1226 = v_1227 & 1'h1;
  assign v_1227 = v_1228 | 1'h0;
  assign v_1228 = ~v_1215;
  assign v_1229 = mux_1229(v_1230);
  assign v_1230 = ~v_1225;
  pebbles_core
    pebbles_core_1231
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1232),
       .in0_consume_en(vin0_consume_en_1231),
       .out_canPeek(vout_canPeek_1231),
       .out_peek(vout_peek_1231));
  assign v_1232 = v_1233 | v_1234;
  assign v_1233 = mux_1233(v_1219);
  assign v_1234 = mux_1234(v_1235);
  assign v_1235 = ~v_1219;
  assign v_1236 = v_1237 & 1'h1;
  assign v_1237 = v_1238 & v_1239;
  assign v_1238 = ~act_1218;
  assign v_1239 = v_1240 | v_1244;
  assign v_1240 = v_1241 | v_1242;
  assign v_1241 = mux_1241(v_1175);
  assign v_1242 = mux_1242(v_1243);
  assign v_1243 = ~v_1175;
  assign v_1244 = ~v_1215;
  assign v_1245 = v_1246 | v_1247;
  assign v_1246 = mux_1246(v_1217);
  assign v_1247 = mux_1247(v_1236);
  assign v_1248 = v_1249 & 1'h1;
  assign v_1249 = v_1250 & v_1251;
  assign v_1250 = ~act_1174;
  assign v_1251 = v_1252 | v_1256;
  assign v_1252 = v_1253 | v_1254;
  assign v_1253 = mux_1253(v_1075);
  assign v_1254 = mux_1254(v_1255);
  assign v_1255 = ~v_1075;
  assign v_1256 = ~v_1171;
  assign v_1257 = v_1258 | v_1259;
  assign v_1258 = mux_1258(v_1173);
  assign v_1259 = mux_1259(v_1248);
  assign v_1260 = v_1261 & 1'h1;
  assign v_1261 = v_1262 & v_1263;
  assign v_1262 = ~act_1074;
  assign v_1263 = v_1264 | v_1268;
  assign v_1264 = v_1265 | v_1266;
  assign v_1265 = mux_1265(v_863);
  assign v_1266 = mux_1266(v_1267);
  assign v_1267 = ~v_863;
  assign v_1268 = ~v_1071;
  assign v_1269 = v_1270 | v_1271;
  assign v_1270 = mux_1270(v_1073);
  assign v_1271 = mux_1271(v_1260);
  assign v_1272 = v_1273 & 1'h1;
  assign v_1273 = v_1274 & v_1275;
  assign v_1274 = ~act_862;
  assign v_1275 = v_1276 | v_1284;
  assign v_1276 = v_1277 | v_1282;
  assign v_1277 = mux_1277(v_1278);
  assign v_1278 = v_859 & v_1279;
  assign v_1279 = v_1280 & 1'h1;
  assign v_1280 = v_1281 | 1'h0;
  assign v_1281 = ~v_852;
  assign v_1282 = mux_1282(v_1283);
  assign v_1283 = ~v_1278;
  assign v_1284 = ~v_859;
  assign v_1285 = v_1286 | v_1287;
  assign v_1286 = mux_1286(v_861);
  assign v_1287 = mux_1287(v_1272);
  assign v_1289 = v_1290 | v_1701;
  assign v_1290 = act_1291 & 1'h1;
  assign act_1291 = v_1292 | v_1490;
  assign v_1292 = v_1293 & v_1491;
  assign v_1293 = v_1294 & v_1500;
  assign v_1294 = ~v_1295;
  assign v_1296 = v_1297 | v_1484;
  assign v_1297 = act_1298 & 1'h1;
  assign act_1298 = v_1299 | v_1385;
  assign v_1299 = v_1300 & v_1386;
  assign v_1300 = v_1301 & v_1395;
  assign v_1301 = ~v_1302;
  assign v_1303 = v_1304 | v_1379;
  assign v_1304 = act_1305 & 1'h1;
  assign act_1305 = v_1306 | v_1336;
  assign v_1306 = v_1307 & v_1337;
  assign v_1307 = v_1308 & v_1346;
  assign v_1308 = ~v_1309;
  assign v_1310 = v_1311 | v_1330;
  assign v_1311 = act_1312 & 1'h1;
  assign act_1312 = v_1313 | v_1319;
  assign v_1313 = v_1314 & v_1320;
  assign v_1314 = v_1315 & vout_canPeek_1325;
  assign v_1315 = ~vout_canPeek_1316;
  pebbles_core
    pebbles_core_1316
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1317),
       .in0_consume_en(vin0_consume_en_1316),
       .out_canPeek(vout_canPeek_1316),
       .out_peek(vout_peek_1316));
  assign v_1317 = v_1318 | v_1323;
  assign v_1318 = mux_1318(v_1319);
  assign v_1319 = vout_canPeek_1316 & v_1320;
  assign v_1320 = v_1321 & 1'h1;
  assign v_1321 = v_1322 | 1'h0;
  assign v_1322 = ~v_1309;
  assign v_1323 = mux_1323(v_1324);
  assign v_1324 = ~v_1319;
  pebbles_core
    pebbles_core_1325
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1326),
       .in0_consume_en(vin0_consume_en_1325),
       .out_canPeek(vout_canPeek_1325),
       .out_peek(vout_peek_1325));
  assign v_1326 = v_1327 | v_1328;
  assign v_1327 = mux_1327(v_1313);
  assign v_1328 = mux_1328(v_1329);
  assign v_1329 = ~v_1313;
  assign v_1330 = v_1331 & 1'h1;
  assign v_1331 = v_1332 & v_1333;
  assign v_1332 = ~act_1312;
  assign v_1333 = v_1334 | v_1342;
  assign v_1334 = v_1335 | v_1340;
  assign v_1335 = mux_1335(v_1336);
  assign v_1336 = v_1309 & v_1337;
  assign v_1337 = v_1338 & 1'h1;
  assign v_1338 = v_1339 | 1'h0;
  assign v_1339 = ~v_1302;
  assign v_1340 = mux_1340(v_1341);
  assign v_1341 = ~v_1336;
  assign v_1342 = ~v_1309;
  assign v_1343 = v_1344 | v_1345;
  assign v_1344 = mux_1344(v_1311);
  assign v_1345 = mux_1345(v_1330);
  assign v_1347 = v_1348 | v_1367;
  assign v_1348 = act_1349 & 1'h1;
  assign act_1349 = v_1350 | v_1356;
  assign v_1350 = v_1351 & v_1357;
  assign v_1351 = v_1352 & vout_canPeek_1362;
  assign v_1352 = ~vout_canPeek_1353;
  pebbles_core
    pebbles_core_1353
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1354),
       .in0_consume_en(vin0_consume_en_1353),
       .out_canPeek(vout_canPeek_1353),
       .out_peek(vout_peek_1353));
  assign v_1354 = v_1355 | v_1360;
  assign v_1355 = mux_1355(v_1356);
  assign v_1356 = vout_canPeek_1353 & v_1357;
  assign v_1357 = v_1358 & 1'h1;
  assign v_1358 = v_1359 | 1'h0;
  assign v_1359 = ~v_1346;
  assign v_1360 = mux_1360(v_1361);
  assign v_1361 = ~v_1356;
  pebbles_core
    pebbles_core_1362
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1363),
       .in0_consume_en(vin0_consume_en_1362),
       .out_canPeek(vout_canPeek_1362),
       .out_peek(vout_peek_1362));
  assign v_1363 = v_1364 | v_1365;
  assign v_1364 = mux_1364(v_1350);
  assign v_1365 = mux_1365(v_1366);
  assign v_1366 = ~v_1350;
  assign v_1367 = v_1368 & 1'h1;
  assign v_1368 = v_1369 & v_1370;
  assign v_1369 = ~act_1349;
  assign v_1370 = v_1371 | v_1375;
  assign v_1371 = v_1372 | v_1373;
  assign v_1372 = mux_1372(v_1306);
  assign v_1373 = mux_1373(v_1374);
  assign v_1374 = ~v_1306;
  assign v_1375 = ~v_1346;
  assign v_1376 = v_1377 | v_1378;
  assign v_1377 = mux_1377(v_1348);
  assign v_1378 = mux_1378(v_1367);
  assign v_1379 = v_1380 & 1'h1;
  assign v_1380 = v_1381 & v_1382;
  assign v_1381 = ~act_1305;
  assign v_1382 = v_1383 | v_1391;
  assign v_1383 = v_1384 | v_1389;
  assign v_1384 = mux_1384(v_1385);
  assign v_1385 = v_1302 & v_1386;
  assign v_1386 = v_1387 & 1'h1;
  assign v_1387 = v_1388 | 1'h0;
  assign v_1388 = ~v_1295;
  assign v_1389 = mux_1389(v_1390);
  assign v_1390 = ~v_1385;
  assign v_1391 = ~v_1302;
  assign v_1392 = v_1393 | v_1394;
  assign v_1393 = mux_1393(v_1304);
  assign v_1394 = mux_1394(v_1379);
  assign v_1396 = v_1397 | v_1472;
  assign v_1397 = act_1398 & 1'h1;
  assign act_1398 = v_1399 | v_1429;
  assign v_1399 = v_1400 & v_1430;
  assign v_1400 = v_1401 & v_1439;
  assign v_1401 = ~v_1402;
  assign v_1403 = v_1404 | v_1423;
  assign v_1404 = act_1405 & 1'h1;
  assign act_1405 = v_1406 | v_1412;
  assign v_1406 = v_1407 & v_1413;
  assign v_1407 = v_1408 & vout_canPeek_1418;
  assign v_1408 = ~vout_canPeek_1409;
  pebbles_core
    pebbles_core_1409
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1410),
       .in0_consume_en(vin0_consume_en_1409),
       .out_canPeek(vout_canPeek_1409),
       .out_peek(vout_peek_1409));
  assign v_1410 = v_1411 | v_1416;
  assign v_1411 = mux_1411(v_1412);
  assign v_1412 = vout_canPeek_1409 & v_1413;
  assign v_1413 = v_1414 & 1'h1;
  assign v_1414 = v_1415 | 1'h0;
  assign v_1415 = ~v_1402;
  assign v_1416 = mux_1416(v_1417);
  assign v_1417 = ~v_1412;
  pebbles_core
    pebbles_core_1418
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1419),
       .in0_consume_en(vin0_consume_en_1418),
       .out_canPeek(vout_canPeek_1418),
       .out_peek(vout_peek_1418));
  assign v_1419 = v_1420 | v_1421;
  assign v_1420 = mux_1420(v_1406);
  assign v_1421 = mux_1421(v_1422);
  assign v_1422 = ~v_1406;
  assign v_1423 = v_1424 & 1'h1;
  assign v_1424 = v_1425 & v_1426;
  assign v_1425 = ~act_1405;
  assign v_1426 = v_1427 | v_1435;
  assign v_1427 = v_1428 | v_1433;
  assign v_1428 = mux_1428(v_1429);
  assign v_1429 = v_1402 & v_1430;
  assign v_1430 = v_1431 & 1'h1;
  assign v_1431 = v_1432 | 1'h0;
  assign v_1432 = ~v_1395;
  assign v_1433 = mux_1433(v_1434);
  assign v_1434 = ~v_1429;
  assign v_1435 = ~v_1402;
  assign v_1436 = v_1437 | v_1438;
  assign v_1437 = mux_1437(v_1404);
  assign v_1438 = mux_1438(v_1423);
  assign v_1440 = v_1441 | v_1460;
  assign v_1441 = act_1442 & 1'h1;
  assign act_1442 = v_1443 | v_1449;
  assign v_1443 = v_1444 & v_1450;
  assign v_1444 = v_1445 & vout_canPeek_1455;
  assign v_1445 = ~vout_canPeek_1446;
  pebbles_core
    pebbles_core_1446
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1447),
       .in0_consume_en(vin0_consume_en_1446),
       .out_canPeek(vout_canPeek_1446),
       .out_peek(vout_peek_1446));
  assign v_1447 = v_1448 | v_1453;
  assign v_1448 = mux_1448(v_1449);
  assign v_1449 = vout_canPeek_1446 & v_1450;
  assign v_1450 = v_1451 & 1'h1;
  assign v_1451 = v_1452 | 1'h0;
  assign v_1452 = ~v_1439;
  assign v_1453 = mux_1453(v_1454);
  assign v_1454 = ~v_1449;
  pebbles_core
    pebbles_core_1455
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1456),
       .in0_consume_en(vin0_consume_en_1455),
       .out_canPeek(vout_canPeek_1455),
       .out_peek(vout_peek_1455));
  assign v_1456 = v_1457 | v_1458;
  assign v_1457 = mux_1457(v_1443);
  assign v_1458 = mux_1458(v_1459);
  assign v_1459 = ~v_1443;
  assign v_1460 = v_1461 & 1'h1;
  assign v_1461 = v_1462 & v_1463;
  assign v_1462 = ~act_1442;
  assign v_1463 = v_1464 | v_1468;
  assign v_1464 = v_1465 | v_1466;
  assign v_1465 = mux_1465(v_1399);
  assign v_1466 = mux_1466(v_1467);
  assign v_1467 = ~v_1399;
  assign v_1468 = ~v_1439;
  assign v_1469 = v_1470 | v_1471;
  assign v_1470 = mux_1470(v_1441);
  assign v_1471 = mux_1471(v_1460);
  assign v_1472 = v_1473 & 1'h1;
  assign v_1473 = v_1474 & v_1475;
  assign v_1474 = ~act_1398;
  assign v_1475 = v_1476 | v_1480;
  assign v_1476 = v_1477 | v_1478;
  assign v_1477 = mux_1477(v_1299);
  assign v_1478 = mux_1478(v_1479);
  assign v_1479 = ~v_1299;
  assign v_1480 = ~v_1395;
  assign v_1481 = v_1482 | v_1483;
  assign v_1482 = mux_1482(v_1397);
  assign v_1483 = mux_1483(v_1472);
  assign v_1484 = v_1485 & 1'h1;
  assign v_1485 = v_1486 & v_1487;
  assign v_1486 = ~act_1298;
  assign v_1487 = v_1488 | v_1496;
  assign v_1488 = v_1489 | v_1494;
  assign v_1489 = mux_1489(v_1490);
  assign v_1490 = v_1295 & v_1491;
  assign v_1491 = v_1492 & 1'h1;
  assign v_1492 = v_1493 | 1'h0;
  assign v_1493 = ~v_1288;
  assign v_1494 = mux_1494(v_1495);
  assign v_1495 = ~v_1490;
  assign v_1496 = ~v_1295;
  assign v_1497 = v_1498 | v_1499;
  assign v_1498 = mux_1498(v_1297);
  assign v_1499 = mux_1499(v_1484);
  assign v_1501 = v_1502 | v_1689;
  assign v_1502 = act_1503 & 1'h1;
  assign act_1503 = v_1504 | v_1590;
  assign v_1504 = v_1505 & v_1591;
  assign v_1505 = v_1506 & v_1600;
  assign v_1506 = ~v_1507;
  assign v_1508 = v_1509 | v_1584;
  assign v_1509 = act_1510 & 1'h1;
  assign act_1510 = v_1511 | v_1541;
  assign v_1511 = v_1512 & v_1542;
  assign v_1512 = v_1513 & v_1551;
  assign v_1513 = ~v_1514;
  assign v_1515 = v_1516 | v_1535;
  assign v_1516 = act_1517 & 1'h1;
  assign act_1517 = v_1518 | v_1524;
  assign v_1518 = v_1519 & v_1525;
  assign v_1519 = v_1520 & vout_canPeek_1530;
  assign v_1520 = ~vout_canPeek_1521;
  pebbles_core
    pebbles_core_1521
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1522),
       .in0_consume_en(vin0_consume_en_1521),
       .out_canPeek(vout_canPeek_1521),
       .out_peek(vout_peek_1521));
  assign v_1522 = v_1523 | v_1528;
  assign v_1523 = mux_1523(v_1524);
  assign v_1524 = vout_canPeek_1521 & v_1525;
  assign v_1525 = v_1526 & 1'h1;
  assign v_1526 = v_1527 | 1'h0;
  assign v_1527 = ~v_1514;
  assign v_1528 = mux_1528(v_1529);
  assign v_1529 = ~v_1524;
  pebbles_core
    pebbles_core_1530
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1531),
       .in0_consume_en(vin0_consume_en_1530),
       .out_canPeek(vout_canPeek_1530),
       .out_peek(vout_peek_1530));
  assign v_1531 = v_1532 | v_1533;
  assign v_1532 = mux_1532(v_1518);
  assign v_1533 = mux_1533(v_1534);
  assign v_1534 = ~v_1518;
  assign v_1535 = v_1536 & 1'h1;
  assign v_1536 = v_1537 & v_1538;
  assign v_1537 = ~act_1517;
  assign v_1538 = v_1539 | v_1547;
  assign v_1539 = v_1540 | v_1545;
  assign v_1540 = mux_1540(v_1541);
  assign v_1541 = v_1514 & v_1542;
  assign v_1542 = v_1543 & 1'h1;
  assign v_1543 = v_1544 | 1'h0;
  assign v_1544 = ~v_1507;
  assign v_1545 = mux_1545(v_1546);
  assign v_1546 = ~v_1541;
  assign v_1547 = ~v_1514;
  assign v_1548 = v_1549 | v_1550;
  assign v_1549 = mux_1549(v_1516);
  assign v_1550 = mux_1550(v_1535);
  assign v_1552 = v_1553 | v_1572;
  assign v_1553 = act_1554 & 1'h1;
  assign act_1554 = v_1555 | v_1561;
  assign v_1555 = v_1556 & v_1562;
  assign v_1556 = v_1557 & vout_canPeek_1567;
  assign v_1557 = ~vout_canPeek_1558;
  pebbles_core
    pebbles_core_1558
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1559),
       .in0_consume_en(vin0_consume_en_1558),
       .out_canPeek(vout_canPeek_1558),
       .out_peek(vout_peek_1558));
  assign v_1559 = v_1560 | v_1565;
  assign v_1560 = mux_1560(v_1561);
  assign v_1561 = vout_canPeek_1558 & v_1562;
  assign v_1562 = v_1563 & 1'h1;
  assign v_1563 = v_1564 | 1'h0;
  assign v_1564 = ~v_1551;
  assign v_1565 = mux_1565(v_1566);
  assign v_1566 = ~v_1561;
  pebbles_core
    pebbles_core_1567
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1568),
       .in0_consume_en(vin0_consume_en_1567),
       .out_canPeek(vout_canPeek_1567),
       .out_peek(vout_peek_1567));
  assign v_1568 = v_1569 | v_1570;
  assign v_1569 = mux_1569(v_1555);
  assign v_1570 = mux_1570(v_1571);
  assign v_1571 = ~v_1555;
  assign v_1572 = v_1573 & 1'h1;
  assign v_1573 = v_1574 & v_1575;
  assign v_1574 = ~act_1554;
  assign v_1575 = v_1576 | v_1580;
  assign v_1576 = v_1577 | v_1578;
  assign v_1577 = mux_1577(v_1511);
  assign v_1578 = mux_1578(v_1579);
  assign v_1579 = ~v_1511;
  assign v_1580 = ~v_1551;
  assign v_1581 = v_1582 | v_1583;
  assign v_1582 = mux_1582(v_1553);
  assign v_1583 = mux_1583(v_1572);
  assign v_1584 = v_1585 & 1'h1;
  assign v_1585 = v_1586 & v_1587;
  assign v_1586 = ~act_1510;
  assign v_1587 = v_1588 | v_1596;
  assign v_1588 = v_1589 | v_1594;
  assign v_1589 = mux_1589(v_1590);
  assign v_1590 = v_1507 & v_1591;
  assign v_1591 = v_1592 & 1'h1;
  assign v_1592 = v_1593 | 1'h0;
  assign v_1593 = ~v_1500;
  assign v_1594 = mux_1594(v_1595);
  assign v_1595 = ~v_1590;
  assign v_1596 = ~v_1507;
  assign v_1597 = v_1598 | v_1599;
  assign v_1598 = mux_1598(v_1509);
  assign v_1599 = mux_1599(v_1584);
  assign v_1601 = v_1602 | v_1677;
  assign v_1602 = act_1603 & 1'h1;
  assign act_1603 = v_1604 | v_1634;
  assign v_1604 = v_1605 & v_1635;
  assign v_1605 = v_1606 & v_1644;
  assign v_1606 = ~v_1607;
  assign v_1608 = v_1609 | v_1628;
  assign v_1609 = act_1610 & 1'h1;
  assign act_1610 = v_1611 | v_1617;
  assign v_1611 = v_1612 & v_1618;
  assign v_1612 = v_1613 & vout_canPeek_1623;
  assign v_1613 = ~vout_canPeek_1614;
  pebbles_core
    pebbles_core_1614
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1615),
       .in0_consume_en(vin0_consume_en_1614),
       .out_canPeek(vout_canPeek_1614),
       .out_peek(vout_peek_1614));
  assign v_1615 = v_1616 | v_1621;
  assign v_1616 = mux_1616(v_1617);
  assign v_1617 = vout_canPeek_1614 & v_1618;
  assign v_1618 = v_1619 & 1'h1;
  assign v_1619 = v_1620 | 1'h0;
  assign v_1620 = ~v_1607;
  assign v_1621 = mux_1621(v_1622);
  assign v_1622 = ~v_1617;
  pebbles_core
    pebbles_core_1623
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1624),
       .in0_consume_en(vin0_consume_en_1623),
       .out_canPeek(vout_canPeek_1623),
       .out_peek(vout_peek_1623));
  assign v_1624 = v_1625 | v_1626;
  assign v_1625 = mux_1625(v_1611);
  assign v_1626 = mux_1626(v_1627);
  assign v_1627 = ~v_1611;
  assign v_1628 = v_1629 & 1'h1;
  assign v_1629 = v_1630 & v_1631;
  assign v_1630 = ~act_1610;
  assign v_1631 = v_1632 | v_1640;
  assign v_1632 = v_1633 | v_1638;
  assign v_1633 = mux_1633(v_1634);
  assign v_1634 = v_1607 & v_1635;
  assign v_1635 = v_1636 & 1'h1;
  assign v_1636 = v_1637 | 1'h0;
  assign v_1637 = ~v_1600;
  assign v_1638 = mux_1638(v_1639);
  assign v_1639 = ~v_1634;
  assign v_1640 = ~v_1607;
  assign v_1641 = v_1642 | v_1643;
  assign v_1642 = mux_1642(v_1609);
  assign v_1643 = mux_1643(v_1628);
  assign v_1645 = v_1646 | v_1665;
  assign v_1646 = act_1647 & 1'h1;
  assign act_1647 = v_1648 | v_1654;
  assign v_1648 = v_1649 & v_1655;
  assign v_1649 = v_1650 & vout_canPeek_1660;
  assign v_1650 = ~vout_canPeek_1651;
  pebbles_core
    pebbles_core_1651
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1652),
       .in0_consume_en(vin0_consume_en_1651),
       .out_canPeek(vout_canPeek_1651),
       .out_peek(vout_peek_1651));
  assign v_1652 = v_1653 | v_1658;
  assign v_1653 = mux_1653(v_1654);
  assign v_1654 = vout_canPeek_1651 & v_1655;
  assign v_1655 = v_1656 & 1'h1;
  assign v_1656 = v_1657 | 1'h0;
  assign v_1657 = ~v_1644;
  assign v_1658 = mux_1658(v_1659);
  assign v_1659 = ~v_1654;
  pebbles_core
    pebbles_core_1660
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1661),
       .in0_consume_en(vin0_consume_en_1660),
       .out_canPeek(vout_canPeek_1660),
       .out_peek(vout_peek_1660));
  assign v_1661 = v_1662 | v_1663;
  assign v_1662 = mux_1662(v_1648);
  assign v_1663 = mux_1663(v_1664);
  assign v_1664 = ~v_1648;
  assign v_1665 = v_1666 & 1'h1;
  assign v_1666 = v_1667 & v_1668;
  assign v_1667 = ~act_1647;
  assign v_1668 = v_1669 | v_1673;
  assign v_1669 = v_1670 | v_1671;
  assign v_1670 = mux_1670(v_1604);
  assign v_1671 = mux_1671(v_1672);
  assign v_1672 = ~v_1604;
  assign v_1673 = ~v_1644;
  assign v_1674 = v_1675 | v_1676;
  assign v_1675 = mux_1675(v_1646);
  assign v_1676 = mux_1676(v_1665);
  assign v_1677 = v_1678 & 1'h1;
  assign v_1678 = v_1679 & v_1680;
  assign v_1679 = ~act_1603;
  assign v_1680 = v_1681 | v_1685;
  assign v_1681 = v_1682 | v_1683;
  assign v_1682 = mux_1682(v_1504);
  assign v_1683 = mux_1683(v_1684);
  assign v_1684 = ~v_1504;
  assign v_1685 = ~v_1600;
  assign v_1686 = v_1687 | v_1688;
  assign v_1687 = mux_1687(v_1602);
  assign v_1688 = mux_1688(v_1677);
  assign v_1689 = v_1690 & 1'h1;
  assign v_1690 = v_1691 & v_1692;
  assign v_1691 = ~act_1503;
  assign v_1692 = v_1693 | v_1697;
  assign v_1693 = v_1694 | v_1695;
  assign v_1694 = mux_1694(v_1292);
  assign v_1695 = mux_1695(v_1696);
  assign v_1696 = ~v_1292;
  assign v_1697 = ~v_1500;
  assign v_1698 = v_1699 | v_1700;
  assign v_1699 = mux_1699(v_1502);
  assign v_1700 = mux_1700(v_1689);
  assign v_1701 = v_1702 & 1'h1;
  assign v_1702 = v_1703 & v_1704;
  assign v_1703 = ~act_1291;
  assign v_1704 = v_1705 | v_1709;
  assign v_1705 = v_1706 | v_1707;
  assign v_1706 = mux_1706(v_856);
  assign v_1707 = mux_1707(v_1708);
  assign v_1708 = ~v_856;
  assign v_1709 = ~v_1288;
  assign v_1710 = v_1711 | v_1712;
  assign v_1711 = mux_1711(v_1290);
  assign v_1712 = mux_1712(v_1701);
  assign v_1713 = v_1714 & 1'h1;
  assign v_1714 = v_1715 & v_1716;
  assign v_1715 = ~act_855;
  assign v_1716 = v_1717 | v_1721;
  assign v_1717 = v_1718 | v_1719;
  assign v_1718 = mux_1718(v_849);
  assign v_1719 = mux_1719(v_1720);
  assign v_1720 = ~v_849;
  assign v_1721 = ~v_852;
  assign v_1722 = v_1723 | v_1724;
  assign v_1723 = mux_1723(v_854);
  assign v_1724 = mux_1724(v_1713);
  assign v_1725 = v_1726 & 1'h1;
  assign v_1726 = v_1727 & v_1728;
  assign v_1727 = ~act_848;
  assign v_1728 = v_1729 | v_22343;
  assign v_1729 = v_1730 | v_22341;
  assign v_1730 = mux_1730(v_1731);
  assign v_1731 = v_1732 & v_2602;
  assign v_1732 = v_1733 & v_845;
  assign v_1733 = ~v_1734;
  assign v_1735 = v_1736 | v_2595;
  assign v_1736 = act_1737 & 1'h1;
  assign act_1737 = v_1738 | v_2160;
  assign v_1738 = v_1739 & v_2161;
  assign v_1739 = v_1740 & v_2170;
  assign v_1740 = ~v_1741;
  assign v_1742 = v_1743 | v_2154;
  assign v_1743 = act_1744 & 1'h1;
  assign act_1744 = v_1745 | v_1943;
  assign v_1745 = v_1746 & v_1944;
  assign v_1746 = v_1747 & v_1953;
  assign v_1747 = ~v_1748;
  assign v_1749 = v_1750 | v_1937;
  assign v_1750 = act_1751 & 1'h1;
  assign act_1751 = v_1752 | v_1838;
  assign v_1752 = v_1753 & v_1839;
  assign v_1753 = v_1754 & v_1848;
  assign v_1754 = ~v_1755;
  assign v_1756 = v_1757 | v_1832;
  assign v_1757 = act_1758 & 1'h1;
  assign act_1758 = v_1759 | v_1789;
  assign v_1759 = v_1760 & v_1790;
  assign v_1760 = v_1761 & v_1799;
  assign v_1761 = ~v_1762;
  assign v_1763 = v_1764 | v_1783;
  assign v_1764 = act_1765 & 1'h1;
  assign act_1765 = v_1766 | v_1772;
  assign v_1766 = v_1767 & v_1773;
  assign v_1767 = v_1768 & vout_canPeek_1778;
  assign v_1768 = ~vout_canPeek_1769;
  pebbles_core
    pebbles_core_1769
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1770),
       .in0_consume_en(vin0_consume_en_1769),
       .out_canPeek(vout_canPeek_1769),
       .out_peek(vout_peek_1769));
  assign v_1770 = v_1771 | v_1776;
  assign v_1771 = mux_1771(v_1772);
  assign v_1772 = vout_canPeek_1769 & v_1773;
  assign v_1773 = v_1774 & 1'h1;
  assign v_1774 = v_1775 | 1'h0;
  assign v_1775 = ~v_1762;
  assign v_1776 = mux_1776(v_1777);
  assign v_1777 = ~v_1772;
  pebbles_core
    pebbles_core_1778
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1779),
       .in0_consume_en(vin0_consume_en_1778),
       .out_canPeek(vout_canPeek_1778),
       .out_peek(vout_peek_1778));
  assign v_1779 = v_1780 | v_1781;
  assign v_1780 = mux_1780(v_1766);
  assign v_1781 = mux_1781(v_1782);
  assign v_1782 = ~v_1766;
  assign v_1783 = v_1784 & 1'h1;
  assign v_1784 = v_1785 & v_1786;
  assign v_1785 = ~act_1765;
  assign v_1786 = v_1787 | v_1795;
  assign v_1787 = v_1788 | v_1793;
  assign v_1788 = mux_1788(v_1789);
  assign v_1789 = v_1762 & v_1790;
  assign v_1790 = v_1791 & 1'h1;
  assign v_1791 = v_1792 | 1'h0;
  assign v_1792 = ~v_1755;
  assign v_1793 = mux_1793(v_1794);
  assign v_1794 = ~v_1789;
  assign v_1795 = ~v_1762;
  assign v_1796 = v_1797 | v_1798;
  assign v_1797 = mux_1797(v_1764);
  assign v_1798 = mux_1798(v_1783);
  assign v_1800 = v_1801 | v_1820;
  assign v_1801 = act_1802 & 1'h1;
  assign act_1802 = v_1803 | v_1809;
  assign v_1803 = v_1804 & v_1810;
  assign v_1804 = v_1805 & vout_canPeek_1815;
  assign v_1805 = ~vout_canPeek_1806;
  pebbles_core
    pebbles_core_1806
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1807),
       .in0_consume_en(vin0_consume_en_1806),
       .out_canPeek(vout_canPeek_1806),
       .out_peek(vout_peek_1806));
  assign v_1807 = v_1808 | v_1813;
  assign v_1808 = mux_1808(v_1809);
  assign v_1809 = vout_canPeek_1806 & v_1810;
  assign v_1810 = v_1811 & 1'h1;
  assign v_1811 = v_1812 | 1'h0;
  assign v_1812 = ~v_1799;
  assign v_1813 = mux_1813(v_1814);
  assign v_1814 = ~v_1809;
  pebbles_core
    pebbles_core_1815
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1816),
       .in0_consume_en(vin0_consume_en_1815),
       .out_canPeek(vout_canPeek_1815),
       .out_peek(vout_peek_1815));
  assign v_1816 = v_1817 | v_1818;
  assign v_1817 = mux_1817(v_1803);
  assign v_1818 = mux_1818(v_1819);
  assign v_1819 = ~v_1803;
  assign v_1820 = v_1821 & 1'h1;
  assign v_1821 = v_1822 & v_1823;
  assign v_1822 = ~act_1802;
  assign v_1823 = v_1824 | v_1828;
  assign v_1824 = v_1825 | v_1826;
  assign v_1825 = mux_1825(v_1759);
  assign v_1826 = mux_1826(v_1827);
  assign v_1827 = ~v_1759;
  assign v_1828 = ~v_1799;
  assign v_1829 = v_1830 | v_1831;
  assign v_1830 = mux_1830(v_1801);
  assign v_1831 = mux_1831(v_1820);
  assign v_1832 = v_1833 & 1'h1;
  assign v_1833 = v_1834 & v_1835;
  assign v_1834 = ~act_1758;
  assign v_1835 = v_1836 | v_1844;
  assign v_1836 = v_1837 | v_1842;
  assign v_1837 = mux_1837(v_1838);
  assign v_1838 = v_1755 & v_1839;
  assign v_1839 = v_1840 & 1'h1;
  assign v_1840 = v_1841 | 1'h0;
  assign v_1841 = ~v_1748;
  assign v_1842 = mux_1842(v_1843);
  assign v_1843 = ~v_1838;
  assign v_1844 = ~v_1755;
  assign v_1845 = v_1846 | v_1847;
  assign v_1846 = mux_1846(v_1757);
  assign v_1847 = mux_1847(v_1832);
  assign v_1849 = v_1850 | v_1925;
  assign v_1850 = act_1851 & 1'h1;
  assign act_1851 = v_1852 | v_1882;
  assign v_1852 = v_1853 & v_1883;
  assign v_1853 = v_1854 & v_1892;
  assign v_1854 = ~v_1855;
  assign v_1856 = v_1857 | v_1876;
  assign v_1857 = act_1858 & 1'h1;
  assign act_1858 = v_1859 | v_1865;
  assign v_1859 = v_1860 & v_1866;
  assign v_1860 = v_1861 & vout_canPeek_1871;
  assign v_1861 = ~vout_canPeek_1862;
  pebbles_core
    pebbles_core_1862
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1863),
       .in0_consume_en(vin0_consume_en_1862),
       .out_canPeek(vout_canPeek_1862),
       .out_peek(vout_peek_1862));
  assign v_1863 = v_1864 | v_1869;
  assign v_1864 = mux_1864(v_1865);
  assign v_1865 = vout_canPeek_1862 & v_1866;
  assign v_1866 = v_1867 & 1'h1;
  assign v_1867 = v_1868 | 1'h0;
  assign v_1868 = ~v_1855;
  assign v_1869 = mux_1869(v_1870);
  assign v_1870 = ~v_1865;
  pebbles_core
    pebbles_core_1871
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1872),
       .in0_consume_en(vin0_consume_en_1871),
       .out_canPeek(vout_canPeek_1871),
       .out_peek(vout_peek_1871));
  assign v_1872 = v_1873 | v_1874;
  assign v_1873 = mux_1873(v_1859);
  assign v_1874 = mux_1874(v_1875);
  assign v_1875 = ~v_1859;
  assign v_1876 = v_1877 & 1'h1;
  assign v_1877 = v_1878 & v_1879;
  assign v_1878 = ~act_1858;
  assign v_1879 = v_1880 | v_1888;
  assign v_1880 = v_1881 | v_1886;
  assign v_1881 = mux_1881(v_1882);
  assign v_1882 = v_1855 & v_1883;
  assign v_1883 = v_1884 & 1'h1;
  assign v_1884 = v_1885 | 1'h0;
  assign v_1885 = ~v_1848;
  assign v_1886 = mux_1886(v_1887);
  assign v_1887 = ~v_1882;
  assign v_1888 = ~v_1855;
  assign v_1889 = v_1890 | v_1891;
  assign v_1890 = mux_1890(v_1857);
  assign v_1891 = mux_1891(v_1876);
  assign v_1893 = v_1894 | v_1913;
  assign v_1894 = act_1895 & 1'h1;
  assign act_1895 = v_1896 | v_1902;
  assign v_1896 = v_1897 & v_1903;
  assign v_1897 = v_1898 & vout_canPeek_1908;
  assign v_1898 = ~vout_canPeek_1899;
  pebbles_core
    pebbles_core_1899
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1900),
       .in0_consume_en(vin0_consume_en_1899),
       .out_canPeek(vout_canPeek_1899),
       .out_peek(vout_peek_1899));
  assign v_1900 = v_1901 | v_1906;
  assign v_1901 = mux_1901(v_1902);
  assign v_1902 = vout_canPeek_1899 & v_1903;
  assign v_1903 = v_1904 & 1'h1;
  assign v_1904 = v_1905 | 1'h0;
  assign v_1905 = ~v_1892;
  assign v_1906 = mux_1906(v_1907);
  assign v_1907 = ~v_1902;
  pebbles_core
    pebbles_core_1908
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1909),
       .in0_consume_en(vin0_consume_en_1908),
       .out_canPeek(vout_canPeek_1908),
       .out_peek(vout_peek_1908));
  assign v_1909 = v_1910 | v_1911;
  assign v_1910 = mux_1910(v_1896);
  assign v_1911 = mux_1911(v_1912);
  assign v_1912 = ~v_1896;
  assign v_1913 = v_1914 & 1'h1;
  assign v_1914 = v_1915 & v_1916;
  assign v_1915 = ~act_1895;
  assign v_1916 = v_1917 | v_1921;
  assign v_1917 = v_1918 | v_1919;
  assign v_1918 = mux_1918(v_1852);
  assign v_1919 = mux_1919(v_1920);
  assign v_1920 = ~v_1852;
  assign v_1921 = ~v_1892;
  assign v_1922 = v_1923 | v_1924;
  assign v_1923 = mux_1923(v_1894);
  assign v_1924 = mux_1924(v_1913);
  assign v_1925 = v_1926 & 1'h1;
  assign v_1926 = v_1927 & v_1928;
  assign v_1927 = ~act_1851;
  assign v_1928 = v_1929 | v_1933;
  assign v_1929 = v_1930 | v_1931;
  assign v_1930 = mux_1930(v_1752);
  assign v_1931 = mux_1931(v_1932);
  assign v_1932 = ~v_1752;
  assign v_1933 = ~v_1848;
  assign v_1934 = v_1935 | v_1936;
  assign v_1935 = mux_1935(v_1850);
  assign v_1936 = mux_1936(v_1925);
  assign v_1937 = v_1938 & 1'h1;
  assign v_1938 = v_1939 & v_1940;
  assign v_1939 = ~act_1751;
  assign v_1940 = v_1941 | v_1949;
  assign v_1941 = v_1942 | v_1947;
  assign v_1942 = mux_1942(v_1943);
  assign v_1943 = v_1748 & v_1944;
  assign v_1944 = v_1945 & 1'h1;
  assign v_1945 = v_1946 | 1'h0;
  assign v_1946 = ~v_1741;
  assign v_1947 = mux_1947(v_1948);
  assign v_1948 = ~v_1943;
  assign v_1949 = ~v_1748;
  assign v_1950 = v_1951 | v_1952;
  assign v_1951 = mux_1951(v_1750);
  assign v_1952 = mux_1952(v_1937);
  assign v_1954 = v_1955 | v_2142;
  assign v_1955 = act_1956 & 1'h1;
  assign act_1956 = v_1957 | v_2043;
  assign v_1957 = v_1958 & v_2044;
  assign v_1958 = v_1959 & v_2053;
  assign v_1959 = ~v_1960;
  assign v_1961 = v_1962 | v_2037;
  assign v_1962 = act_1963 & 1'h1;
  assign act_1963 = v_1964 | v_1994;
  assign v_1964 = v_1965 & v_1995;
  assign v_1965 = v_1966 & v_2004;
  assign v_1966 = ~v_1967;
  assign v_1968 = v_1969 | v_1988;
  assign v_1969 = act_1970 & 1'h1;
  assign act_1970 = v_1971 | v_1977;
  assign v_1971 = v_1972 & v_1978;
  assign v_1972 = v_1973 & vout_canPeek_1983;
  assign v_1973 = ~vout_canPeek_1974;
  pebbles_core
    pebbles_core_1974
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1975),
       .in0_consume_en(vin0_consume_en_1974),
       .out_canPeek(vout_canPeek_1974),
       .out_peek(vout_peek_1974));
  assign v_1975 = v_1976 | v_1981;
  assign v_1976 = mux_1976(v_1977);
  assign v_1977 = vout_canPeek_1974 & v_1978;
  assign v_1978 = v_1979 & 1'h1;
  assign v_1979 = v_1980 | 1'h0;
  assign v_1980 = ~v_1967;
  assign v_1981 = mux_1981(v_1982);
  assign v_1982 = ~v_1977;
  pebbles_core
    pebbles_core_1983
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1984),
       .in0_consume_en(vin0_consume_en_1983),
       .out_canPeek(vout_canPeek_1983),
       .out_peek(vout_peek_1983));
  assign v_1984 = v_1985 | v_1986;
  assign v_1985 = mux_1985(v_1971);
  assign v_1986 = mux_1986(v_1987);
  assign v_1987 = ~v_1971;
  assign v_1988 = v_1989 & 1'h1;
  assign v_1989 = v_1990 & v_1991;
  assign v_1990 = ~act_1970;
  assign v_1991 = v_1992 | v_2000;
  assign v_1992 = v_1993 | v_1998;
  assign v_1993 = mux_1993(v_1994);
  assign v_1994 = v_1967 & v_1995;
  assign v_1995 = v_1996 & 1'h1;
  assign v_1996 = v_1997 | 1'h0;
  assign v_1997 = ~v_1960;
  assign v_1998 = mux_1998(v_1999);
  assign v_1999 = ~v_1994;
  assign v_2000 = ~v_1967;
  assign v_2001 = v_2002 | v_2003;
  assign v_2002 = mux_2002(v_1969);
  assign v_2003 = mux_2003(v_1988);
  assign v_2005 = v_2006 | v_2025;
  assign v_2006 = act_2007 & 1'h1;
  assign act_2007 = v_2008 | v_2014;
  assign v_2008 = v_2009 & v_2015;
  assign v_2009 = v_2010 & vout_canPeek_2020;
  assign v_2010 = ~vout_canPeek_2011;
  pebbles_core
    pebbles_core_2011
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2012),
       .in0_consume_en(vin0_consume_en_2011),
       .out_canPeek(vout_canPeek_2011),
       .out_peek(vout_peek_2011));
  assign v_2012 = v_2013 | v_2018;
  assign v_2013 = mux_2013(v_2014);
  assign v_2014 = vout_canPeek_2011 & v_2015;
  assign v_2015 = v_2016 & 1'h1;
  assign v_2016 = v_2017 | 1'h0;
  assign v_2017 = ~v_2004;
  assign v_2018 = mux_2018(v_2019);
  assign v_2019 = ~v_2014;
  pebbles_core
    pebbles_core_2020
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2021),
       .in0_consume_en(vin0_consume_en_2020),
       .out_canPeek(vout_canPeek_2020),
       .out_peek(vout_peek_2020));
  assign v_2021 = v_2022 | v_2023;
  assign v_2022 = mux_2022(v_2008);
  assign v_2023 = mux_2023(v_2024);
  assign v_2024 = ~v_2008;
  assign v_2025 = v_2026 & 1'h1;
  assign v_2026 = v_2027 & v_2028;
  assign v_2027 = ~act_2007;
  assign v_2028 = v_2029 | v_2033;
  assign v_2029 = v_2030 | v_2031;
  assign v_2030 = mux_2030(v_1964);
  assign v_2031 = mux_2031(v_2032);
  assign v_2032 = ~v_1964;
  assign v_2033 = ~v_2004;
  assign v_2034 = v_2035 | v_2036;
  assign v_2035 = mux_2035(v_2006);
  assign v_2036 = mux_2036(v_2025);
  assign v_2037 = v_2038 & 1'h1;
  assign v_2038 = v_2039 & v_2040;
  assign v_2039 = ~act_1963;
  assign v_2040 = v_2041 | v_2049;
  assign v_2041 = v_2042 | v_2047;
  assign v_2042 = mux_2042(v_2043);
  assign v_2043 = v_1960 & v_2044;
  assign v_2044 = v_2045 & 1'h1;
  assign v_2045 = v_2046 | 1'h0;
  assign v_2046 = ~v_1953;
  assign v_2047 = mux_2047(v_2048);
  assign v_2048 = ~v_2043;
  assign v_2049 = ~v_1960;
  assign v_2050 = v_2051 | v_2052;
  assign v_2051 = mux_2051(v_1962);
  assign v_2052 = mux_2052(v_2037);
  assign v_2054 = v_2055 | v_2130;
  assign v_2055 = act_2056 & 1'h1;
  assign act_2056 = v_2057 | v_2087;
  assign v_2057 = v_2058 & v_2088;
  assign v_2058 = v_2059 & v_2097;
  assign v_2059 = ~v_2060;
  assign v_2061 = v_2062 | v_2081;
  assign v_2062 = act_2063 & 1'h1;
  assign act_2063 = v_2064 | v_2070;
  assign v_2064 = v_2065 & v_2071;
  assign v_2065 = v_2066 & vout_canPeek_2076;
  assign v_2066 = ~vout_canPeek_2067;
  pebbles_core
    pebbles_core_2067
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2068),
       .in0_consume_en(vin0_consume_en_2067),
       .out_canPeek(vout_canPeek_2067),
       .out_peek(vout_peek_2067));
  assign v_2068 = v_2069 | v_2074;
  assign v_2069 = mux_2069(v_2070);
  assign v_2070 = vout_canPeek_2067 & v_2071;
  assign v_2071 = v_2072 & 1'h1;
  assign v_2072 = v_2073 | 1'h0;
  assign v_2073 = ~v_2060;
  assign v_2074 = mux_2074(v_2075);
  assign v_2075 = ~v_2070;
  pebbles_core
    pebbles_core_2076
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2077),
       .in0_consume_en(vin0_consume_en_2076),
       .out_canPeek(vout_canPeek_2076),
       .out_peek(vout_peek_2076));
  assign v_2077 = v_2078 | v_2079;
  assign v_2078 = mux_2078(v_2064);
  assign v_2079 = mux_2079(v_2080);
  assign v_2080 = ~v_2064;
  assign v_2081 = v_2082 & 1'h1;
  assign v_2082 = v_2083 & v_2084;
  assign v_2083 = ~act_2063;
  assign v_2084 = v_2085 | v_2093;
  assign v_2085 = v_2086 | v_2091;
  assign v_2086 = mux_2086(v_2087);
  assign v_2087 = v_2060 & v_2088;
  assign v_2088 = v_2089 & 1'h1;
  assign v_2089 = v_2090 | 1'h0;
  assign v_2090 = ~v_2053;
  assign v_2091 = mux_2091(v_2092);
  assign v_2092 = ~v_2087;
  assign v_2093 = ~v_2060;
  assign v_2094 = v_2095 | v_2096;
  assign v_2095 = mux_2095(v_2062);
  assign v_2096 = mux_2096(v_2081);
  assign v_2098 = v_2099 | v_2118;
  assign v_2099 = act_2100 & 1'h1;
  assign act_2100 = v_2101 | v_2107;
  assign v_2101 = v_2102 & v_2108;
  assign v_2102 = v_2103 & vout_canPeek_2113;
  assign v_2103 = ~vout_canPeek_2104;
  pebbles_core
    pebbles_core_2104
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2105),
       .in0_consume_en(vin0_consume_en_2104),
       .out_canPeek(vout_canPeek_2104),
       .out_peek(vout_peek_2104));
  assign v_2105 = v_2106 | v_2111;
  assign v_2106 = mux_2106(v_2107);
  assign v_2107 = vout_canPeek_2104 & v_2108;
  assign v_2108 = v_2109 & 1'h1;
  assign v_2109 = v_2110 | 1'h0;
  assign v_2110 = ~v_2097;
  assign v_2111 = mux_2111(v_2112);
  assign v_2112 = ~v_2107;
  pebbles_core
    pebbles_core_2113
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2114),
       .in0_consume_en(vin0_consume_en_2113),
       .out_canPeek(vout_canPeek_2113),
       .out_peek(vout_peek_2113));
  assign v_2114 = v_2115 | v_2116;
  assign v_2115 = mux_2115(v_2101);
  assign v_2116 = mux_2116(v_2117);
  assign v_2117 = ~v_2101;
  assign v_2118 = v_2119 & 1'h1;
  assign v_2119 = v_2120 & v_2121;
  assign v_2120 = ~act_2100;
  assign v_2121 = v_2122 | v_2126;
  assign v_2122 = v_2123 | v_2124;
  assign v_2123 = mux_2123(v_2057);
  assign v_2124 = mux_2124(v_2125);
  assign v_2125 = ~v_2057;
  assign v_2126 = ~v_2097;
  assign v_2127 = v_2128 | v_2129;
  assign v_2128 = mux_2128(v_2099);
  assign v_2129 = mux_2129(v_2118);
  assign v_2130 = v_2131 & 1'h1;
  assign v_2131 = v_2132 & v_2133;
  assign v_2132 = ~act_2056;
  assign v_2133 = v_2134 | v_2138;
  assign v_2134 = v_2135 | v_2136;
  assign v_2135 = mux_2135(v_1957);
  assign v_2136 = mux_2136(v_2137);
  assign v_2137 = ~v_1957;
  assign v_2138 = ~v_2053;
  assign v_2139 = v_2140 | v_2141;
  assign v_2140 = mux_2140(v_2055);
  assign v_2141 = mux_2141(v_2130);
  assign v_2142 = v_2143 & 1'h1;
  assign v_2143 = v_2144 & v_2145;
  assign v_2144 = ~act_1956;
  assign v_2145 = v_2146 | v_2150;
  assign v_2146 = v_2147 | v_2148;
  assign v_2147 = mux_2147(v_1745);
  assign v_2148 = mux_2148(v_2149);
  assign v_2149 = ~v_1745;
  assign v_2150 = ~v_1953;
  assign v_2151 = v_2152 | v_2153;
  assign v_2152 = mux_2152(v_1955);
  assign v_2153 = mux_2153(v_2142);
  assign v_2154 = v_2155 & 1'h1;
  assign v_2155 = v_2156 & v_2157;
  assign v_2156 = ~act_1744;
  assign v_2157 = v_2158 | v_2166;
  assign v_2158 = v_2159 | v_2164;
  assign v_2159 = mux_2159(v_2160);
  assign v_2160 = v_1741 & v_2161;
  assign v_2161 = v_2162 & 1'h1;
  assign v_2162 = v_2163 | 1'h0;
  assign v_2163 = ~v_1734;
  assign v_2164 = mux_2164(v_2165);
  assign v_2165 = ~v_2160;
  assign v_2166 = ~v_1741;
  assign v_2167 = v_2168 | v_2169;
  assign v_2168 = mux_2168(v_1743);
  assign v_2169 = mux_2169(v_2154);
  assign v_2171 = v_2172 | v_2583;
  assign v_2172 = act_2173 & 1'h1;
  assign act_2173 = v_2174 | v_2372;
  assign v_2174 = v_2175 & v_2373;
  assign v_2175 = v_2176 & v_2382;
  assign v_2176 = ~v_2177;
  assign v_2178 = v_2179 | v_2366;
  assign v_2179 = act_2180 & 1'h1;
  assign act_2180 = v_2181 | v_2267;
  assign v_2181 = v_2182 & v_2268;
  assign v_2182 = v_2183 & v_2277;
  assign v_2183 = ~v_2184;
  assign v_2185 = v_2186 | v_2261;
  assign v_2186 = act_2187 & 1'h1;
  assign act_2187 = v_2188 | v_2218;
  assign v_2188 = v_2189 & v_2219;
  assign v_2189 = v_2190 & v_2228;
  assign v_2190 = ~v_2191;
  assign v_2192 = v_2193 | v_2212;
  assign v_2193 = act_2194 & 1'h1;
  assign act_2194 = v_2195 | v_2201;
  assign v_2195 = v_2196 & v_2202;
  assign v_2196 = v_2197 & vout_canPeek_2207;
  assign v_2197 = ~vout_canPeek_2198;
  pebbles_core
    pebbles_core_2198
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2199),
       .in0_consume_en(vin0_consume_en_2198),
       .out_canPeek(vout_canPeek_2198),
       .out_peek(vout_peek_2198));
  assign v_2199 = v_2200 | v_2205;
  assign v_2200 = mux_2200(v_2201);
  assign v_2201 = vout_canPeek_2198 & v_2202;
  assign v_2202 = v_2203 & 1'h1;
  assign v_2203 = v_2204 | 1'h0;
  assign v_2204 = ~v_2191;
  assign v_2205 = mux_2205(v_2206);
  assign v_2206 = ~v_2201;
  pebbles_core
    pebbles_core_2207
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2208),
       .in0_consume_en(vin0_consume_en_2207),
       .out_canPeek(vout_canPeek_2207),
       .out_peek(vout_peek_2207));
  assign v_2208 = v_2209 | v_2210;
  assign v_2209 = mux_2209(v_2195);
  assign v_2210 = mux_2210(v_2211);
  assign v_2211 = ~v_2195;
  assign v_2212 = v_2213 & 1'h1;
  assign v_2213 = v_2214 & v_2215;
  assign v_2214 = ~act_2194;
  assign v_2215 = v_2216 | v_2224;
  assign v_2216 = v_2217 | v_2222;
  assign v_2217 = mux_2217(v_2218);
  assign v_2218 = v_2191 & v_2219;
  assign v_2219 = v_2220 & 1'h1;
  assign v_2220 = v_2221 | 1'h0;
  assign v_2221 = ~v_2184;
  assign v_2222 = mux_2222(v_2223);
  assign v_2223 = ~v_2218;
  assign v_2224 = ~v_2191;
  assign v_2225 = v_2226 | v_2227;
  assign v_2226 = mux_2226(v_2193);
  assign v_2227 = mux_2227(v_2212);
  assign v_2229 = v_2230 | v_2249;
  assign v_2230 = act_2231 & 1'h1;
  assign act_2231 = v_2232 | v_2238;
  assign v_2232 = v_2233 & v_2239;
  assign v_2233 = v_2234 & vout_canPeek_2244;
  assign v_2234 = ~vout_canPeek_2235;
  pebbles_core
    pebbles_core_2235
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2236),
       .in0_consume_en(vin0_consume_en_2235),
       .out_canPeek(vout_canPeek_2235),
       .out_peek(vout_peek_2235));
  assign v_2236 = v_2237 | v_2242;
  assign v_2237 = mux_2237(v_2238);
  assign v_2238 = vout_canPeek_2235 & v_2239;
  assign v_2239 = v_2240 & 1'h1;
  assign v_2240 = v_2241 | 1'h0;
  assign v_2241 = ~v_2228;
  assign v_2242 = mux_2242(v_2243);
  assign v_2243 = ~v_2238;
  pebbles_core
    pebbles_core_2244
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2245),
       .in0_consume_en(vin0_consume_en_2244),
       .out_canPeek(vout_canPeek_2244),
       .out_peek(vout_peek_2244));
  assign v_2245 = v_2246 | v_2247;
  assign v_2246 = mux_2246(v_2232);
  assign v_2247 = mux_2247(v_2248);
  assign v_2248 = ~v_2232;
  assign v_2249 = v_2250 & 1'h1;
  assign v_2250 = v_2251 & v_2252;
  assign v_2251 = ~act_2231;
  assign v_2252 = v_2253 | v_2257;
  assign v_2253 = v_2254 | v_2255;
  assign v_2254 = mux_2254(v_2188);
  assign v_2255 = mux_2255(v_2256);
  assign v_2256 = ~v_2188;
  assign v_2257 = ~v_2228;
  assign v_2258 = v_2259 | v_2260;
  assign v_2259 = mux_2259(v_2230);
  assign v_2260 = mux_2260(v_2249);
  assign v_2261 = v_2262 & 1'h1;
  assign v_2262 = v_2263 & v_2264;
  assign v_2263 = ~act_2187;
  assign v_2264 = v_2265 | v_2273;
  assign v_2265 = v_2266 | v_2271;
  assign v_2266 = mux_2266(v_2267);
  assign v_2267 = v_2184 & v_2268;
  assign v_2268 = v_2269 & 1'h1;
  assign v_2269 = v_2270 | 1'h0;
  assign v_2270 = ~v_2177;
  assign v_2271 = mux_2271(v_2272);
  assign v_2272 = ~v_2267;
  assign v_2273 = ~v_2184;
  assign v_2274 = v_2275 | v_2276;
  assign v_2275 = mux_2275(v_2186);
  assign v_2276 = mux_2276(v_2261);
  assign v_2278 = v_2279 | v_2354;
  assign v_2279 = act_2280 & 1'h1;
  assign act_2280 = v_2281 | v_2311;
  assign v_2281 = v_2282 & v_2312;
  assign v_2282 = v_2283 & v_2321;
  assign v_2283 = ~v_2284;
  assign v_2285 = v_2286 | v_2305;
  assign v_2286 = act_2287 & 1'h1;
  assign act_2287 = v_2288 | v_2294;
  assign v_2288 = v_2289 & v_2295;
  assign v_2289 = v_2290 & vout_canPeek_2300;
  assign v_2290 = ~vout_canPeek_2291;
  pebbles_core
    pebbles_core_2291
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2292),
       .in0_consume_en(vin0_consume_en_2291),
       .out_canPeek(vout_canPeek_2291),
       .out_peek(vout_peek_2291));
  assign v_2292 = v_2293 | v_2298;
  assign v_2293 = mux_2293(v_2294);
  assign v_2294 = vout_canPeek_2291 & v_2295;
  assign v_2295 = v_2296 & 1'h1;
  assign v_2296 = v_2297 | 1'h0;
  assign v_2297 = ~v_2284;
  assign v_2298 = mux_2298(v_2299);
  assign v_2299 = ~v_2294;
  pebbles_core
    pebbles_core_2300
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2301),
       .in0_consume_en(vin0_consume_en_2300),
       .out_canPeek(vout_canPeek_2300),
       .out_peek(vout_peek_2300));
  assign v_2301 = v_2302 | v_2303;
  assign v_2302 = mux_2302(v_2288);
  assign v_2303 = mux_2303(v_2304);
  assign v_2304 = ~v_2288;
  assign v_2305 = v_2306 & 1'h1;
  assign v_2306 = v_2307 & v_2308;
  assign v_2307 = ~act_2287;
  assign v_2308 = v_2309 | v_2317;
  assign v_2309 = v_2310 | v_2315;
  assign v_2310 = mux_2310(v_2311);
  assign v_2311 = v_2284 & v_2312;
  assign v_2312 = v_2313 & 1'h1;
  assign v_2313 = v_2314 | 1'h0;
  assign v_2314 = ~v_2277;
  assign v_2315 = mux_2315(v_2316);
  assign v_2316 = ~v_2311;
  assign v_2317 = ~v_2284;
  assign v_2318 = v_2319 | v_2320;
  assign v_2319 = mux_2319(v_2286);
  assign v_2320 = mux_2320(v_2305);
  assign v_2322 = v_2323 | v_2342;
  assign v_2323 = act_2324 & 1'h1;
  assign act_2324 = v_2325 | v_2331;
  assign v_2325 = v_2326 & v_2332;
  assign v_2326 = v_2327 & vout_canPeek_2337;
  assign v_2327 = ~vout_canPeek_2328;
  pebbles_core
    pebbles_core_2328
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2329),
       .in0_consume_en(vin0_consume_en_2328),
       .out_canPeek(vout_canPeek_2328),
       .out_peek(vout_peek_2328));
  assign v_2329 = v_2330 | v_2335;
  assign v_2330 = mux_2330(v_2331);
  assign v_2331 = vout_canPeek_2328 & v_2332;
  assign v_2332 = v_2333 & 1'h1;
  assign v_2333 = v_2334 | 1'h0;
  assign v_2334 = ~v_2321;
  assign v_2335 = mux_2335(v_2336);
  assign v_2336 = ~v_2331;
  pebbles_core
    pebbles_core_2337
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2338),
       .in0_consume_en(vin0_consume_en_2337),
       .out_canPeek(vout_canPeek_2337),
       .out_peek(vout_peek_2337));
  assign v_2338 = v_2339 | v_2340;
  assign v_2339 = mux_2339(v_2325);
  assign v_2340 = mux_2340(v_2341);
  assign v_2341 = ~v_2325;
  assign v_2342 = v_2343 & 1'h1;
  assign v_2343 = v_2344 & v_2345;
  assign v_2344 = ~act_2324;
  assign v_2345 = v_2346 | v_2350;
  assign v_2346 = v_2347 | v_2348;
  assign v_2347 = mux_2347(v_2281);
  assign v_2348 = mux_2348(v_2349);
  assign v_2349 = ~v_2281;
  assign v_2350 = ~v_2321;
  assign v_2351 = v_2352 | v_2353;
  assign v_2352 = mux_2352(v_2323);
  assign v_2353 = mux_2353(v_2342);
  assign v_2354 = v_2355 & 1'h1;
  assign v_2355 = v_2356 & v_2357;
  assign v_2356 = ~act_2280;
  assign v_2357 = v_2358 | v_2362;
  assign v_2358 = v_2359 | v_2360;
  assign v_2359 = mux_2359(v_2181);
  assign v_2360 = mux_2360(v_2361);
  assign v_2361 = ~v_2181;
  assign v_2362 = ~v_2277;
  assign v_2363 = v_2364 | v_2365;
  assign v_2364 = mux_2364(v_2279);
  assign v_2365 = mux_2365(v_2354);
  assign v_2366 = v_2367 & 1'h1;
  assign v_2367 = v_2368 & v_2369;
  assign v_2368 = ~act_2180;
  assign v_2369 = v_2370 | v_2378;
  assign v_2370 = v_2371 | v_2376;
  assign v_2371 = mux_2371(v_2372);
  assign v_2372 = v_2177 & v_2373;
  assign v_2373 = v_2374 & 1'h1;
  assign v_2374 = v_2375 | 1'h0;
  assign v_2375 = ~v_2170;
  assign v_2376 = mux_2376(v_2377);
  assign v_2377 = ~v_2372;
  assign v_2378 = ~v_2177;
  assign v_2379 = v_2380 | v_2381;
  assign v_2380 = mux_2380(v_2179);
  assign v_2381 = mux_2381(v_2366);
  assign v_2383 = v_2384 | v_2571;
  assign v_2384 = act_2385 & 1'h1;
  assign act_2385 = v_2386 | v_2472;
  assign v_2386 = v_2387 & v_2473;
  assign v_2387 = v_2388 & v_2482;
  assign v_2388 = ~v_2389;
  assign v_2390 = v_2391 | v_2466;
  assign v_2391 = act_2392 & 1'h1;
  assign act_2392 = v_2393 | v_2423;
  assign v_2393 = v_2394 & v_2424;
  assign v_2394 = v_2395 & v_2433;
  assign v_2395 = ~v_2396;
  assign v_2397 = v_2398 | v_2417;
  assign v_2398 = act_2399 & 1'h1;
  assign act_2399 = v_2400 | v_2406;
  assign v_2400 = v_2401 & v_2407;
  assign v_2401 = v_2402 & vout_canPeek_2412;
  assign v_2402 = ~vout_canPeek_2403;
  pebbles_core
    pebbles_core_2403
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2404),
       .in0_consume_en(vin0_consume_en_2403),
       .out_canPeek(vout_canPeek_2403),
       .out_peek(vout_peek_2403));
  assign v_2404 = v_2405 | v_2410;
  assign v_2405 = mux_2405(v_2406);
  assign v_2406 = vout_canPeek_2403 & v_2407;
  assign v_2407 = v_2408 & 1'h1;
  assign v_2408 = v_2409 | 1'h0;
  assign v_2409 = ~v_2396;
  assign v_2410 = mux_2410(v_2411);
  assign v_2411 = ~v_2406;
  pebbles_core
    pebbles_core_2412
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2413),
       .in0_consume_en(vin0_consume_en_2412),
       .out_canPeek(vout_canPeek_2412),
       .out_peek(vout_peek_2412));
  assign v_2413 = v_2414 | v_2415;
  assign v_2414 = mux_2414(v_2400);
  assign v_2415 = mux_2415(v_2416);
  assign v_2416 = ~v_2400;
  assign v_2417 = v_2418 & 1'h1;
  assign v_2418 = v_2419 & v_2420;
  assign v_2419 = ~act_2399;
  assign v_2420 = v_2421 | v_2429;
  assign v_2421 = v_2422 | v_2427;
  assign v_2422 = mux_2422(v_2423);
  assign v_2423 = v_2396 & v_2424;
  assign v_2424 = v_2425 & 1'h1;
  assign v_2425 = v_2426 | 1'h0;
  assign v_2426 = ~v_2389;
  assign v_2427 = mux_2427(v_2428);
  assign v_2428 = ~v_2423;
  assign v_2429 = ~v_2396;
  assign v_2430 = v_2431 | v_2432;
  assign v_2431 = mux_2431(v_2398);
  assign v_2432 = mux_2432(v_2417);
  assign v_2434 = v_2435 | v_2454;
  assign v_2435 = act_2436 & 1'h1;
  assign act_2436 = v_2437 | v_2443;
  assign v_2437 = v_2438 & v_2444;
  assign v_2438 = v_2439 & vout_canPeek_2449;
  assign v_2439 = ~vout_canPeek_2440;
  pebbles_core
    pebbles_core_2440
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2441),
       .in0_consume_en(vin0_consume_en_2440),
       .out_canPeek(vout_canPeek_2440),
       .out_peek(vout_peek_2440));
  assign v_2441 = v_2442 | v_2447;
  assign v_2442 = mux_2442(v_2443);
  assign v_2443 = vout_canPeek_2440 & v_2444;
  assign v_2444 = v_2445 & 1'h1;
  assign v_2445 = v_2446 | 1'h0;
  assign v_2446 = ~v_2433;
  assign v_2447 = mux_2447(v_2448);
  assign v_2448 = ~v_2443;
  pebbles_core
    pebbles_core_2449
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2450),
       .in0_consume_en(vin0_consume_en_2449),
       .out_canPeek(vout_canPeek_2449),
       .out_peek(vout_peek_2449));
  assign v_2450 = v_2451 | v_2452;
  assign v_2451 = mux_2451(v_2437);
  assign v_2452 = mux_2452(v_2453);
  assign v_2453 = ~v_2437;
  assign v_2454 = v_2455 & 1'h1;
  assign v_2455 = v_2456 & v_2457;
  assign v_2456 = ~act_2436;
  assign v_2457 = v_2458 | v_2462;
  assign v_2458 = v_2459 | v_2460;
  assign v_2459 = mux_2459(v_2393);
  assign v_2460 = mux_2460(v_2461);
  assign v_2461 = ~v_2393;
  assign v_2462 = ~v_2433;
  assign v_2463 = v_2464 | v_2465;
  assign v_2464 = mux_2464(v_2435);
  assign v_2465 = mux_2465(v_2454);
  assign v_2466 = v_2467 & 1'h1;
  assign v_2467 = v_2468 & v_2469;
  assign v_2468 = ~act_2392;
  assign v_2469 = v_2470 | v_2478;
  assign v_2470 = v_2471 | v_2476;
  assign v_2471 = mux_2471(v_2472);
  assign v_2472 = v_2389 & v_2473;
  assign v_2473 = v_2474 & 1'h1;
  assign v_2474 = v_2475 | 1'h0;
  assign v_2475 = ~v_2382;
  assign v_2476 = mux_2476(v_2477);
  assign v_2477 = ~v_2472;
  assign v_2478 = ~v_2389;
  assign v_2479 = v_2480 | v_2481;
  assign v_2480 = mux_2480(v_2391);
  assign v_2481 = mux_2481(v_2466);
  assign v_2483 = v_2484 | v_2559;
  assign v_2484 = act_2485 & 1'h1;
  assign act_2485 = v_2486 | v_2516;
  assign v_2486 = v_2487 & v_2517;
  assign v_2487 = v_2488 & v_2526;
  assign v_2488 = ~v_2489;
  assign v_2490 = v_2491 | v_2510;
  assign v_2491 = act_2492 & 1'h1;
  assign act_2492 = v_2493 | v_2499;
  assign v_2493 = v_2494 & v_2500;
  assign v_2494 = v_2495 & vout_canPeek_2505;
  assign v_2495 = ~vout_canPeek_2496;
  pebbles_core
    pebbles_core_2496
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2497),
       .in0_consume_en(vin0_consume_en_2496),
       .out_canPeek(vout_canPeek_2496),
       .out_peek(vout_peek_2496));
  assign v_2497 = v_2498 | v_2503;
  assign v_2498 = mux_2498(v_2499);
  assign v_2499 = vout_canPeek_2496 & v_2500;
  assign v_2500 = v_2501 & 1'h1;
  assign v_2501 = v_2502 | 1'h0;
  assign v_2502 = ~v_2489;
  assign v_2503 = mux_2503(v_2504);
  assign v_2504 = ~v_2499;
  pebbles_core
    pebbles_core_2505
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2506),
       .in0_consume_en(vin0_consume_en_2505),
       .out_canPeek(vout_canPeek_2505),
       .out_peek(vout_peek_2505));
  assign v_2506 = v_2507 | v_2508;
  assign v_2507 = mux_2507(v_2493);
  assign v_2508 = mux_2508(v_2509);
  assign v_2509 = ~v_2493;
  assign v_2510 = v_2511 & 1'h1;
  assign v_2511 = v_2512 & v_2513;
  assign v_2512 = ~act_2492;
  assign v_2513 = v_2514 | v_2522;
  assign v_2514 = v_2515 | v_2520;
  assign v_2515 = mux_2515(v_2516);
  assign v_2516 = v_2489 & v_2517;
  assign v_2517 = v_2518 & 1'h1;
  assign v_2518 = v_2519 | 1'h0;
  assign v_2519 = ~v_2482;
  assign v_2520 = mux_2520(v_2521);
  assign v_2521 = ~v_2516;
  assign v_2522 = ~v_2489;
  assign v_2523 = v_2524 | v_2525;
  assign v_2524 = mux_2524(v_2491);
  assign v_2525 = mux_2525(v_2510);
  assign v_2527 = v_2528 | v_2547;
  assign v_2528 = act_2529 & 1'h1;
  assign act_2529 = v_2530 | v_2536;
  assign v_2530 = v_2531 & v_2537;
  assign v_2531 = v_2532 & vout_canPeek_2542;
  assign v_2532 = ~vout_canPeek_2533;
  pebbles_core
    pebbles_core_2533
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2534),
       .in0_consume_en(vin0_consume_en_2533),
       .out_canPeek(vout_canPeek_2533),
       .out_peek(vout_peek_2533));
  assign v_2534 = v_2535 | v_2540;
  assign v_2535 = mux_2535(v_2536);
  assign v_2536 = vout_canPeek_2533 & v_2537;
  assign v_2537 = v_2538 & 1'h1;
  assign v_2538 = v_2539 | 1'h0;
  assign v_2539 = ~v_2526;
  assign v_2540 = mux_2540(v_2541);
  assign v_2541 = ~v_2536;
  pebbles_core
    pebbles_core_2542
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2543),
       .in0_consume_en(vin0_consume_en_2542),
       .out_canPeek(vout_canPeek_2542),
       .out_peek(vout_peek_2542));
  assign v_2543 = v_2544 | v_2545;
  assign v_2544 = mux_2544(v_2530);
  assign v_2545 = mux_2545(v_2546);
  assign v_2546 = ~v_2530;
  assign v_2547 = v_2548 & 1'h1;
  assign v_2548 = v_2549 & v_2550;
  assign v_2549 = ~act_2529;
  assign v_2550 = v_2551 | v_2555;
  assign v_2551 = v_2552 | v_2553;
  assign v_2552 = mux_2552(v_2486);
  assign v_2553 = mux_2553(v_2554);
  assign v_2554 = ~v_2486;
  assign v_2555 = ~v_2526;
  assign v_2556 = v_2557 | v_2558;
  assign v_2557 = mux_2557(v_2528);
  assign v_2558 = mux_2558(v_2547);
  assign v_2559 = v_2560 & 1'h1;
  assign v_2560 = v_2561 & v_2562;
  assign v_2561 = ~act_2485;
  assign v_2562 = v_2563 | v_2567;
  assign v_2563 = v_2564 | v_2565;
  assign v_2564 = mux_2564(v_2386);
  assign v_2565 = mux_2565(v_2566);
  assign v_2566 = ~v_2386;
  assign v_2567 = ~v_2482;
  assign v_2568 = v_2569 | v_2570;
  assign v_2569 = mux_2569(v_2484);
  assign v_2570 = mux_2570(v_2559);
  assign v_2571 = v_2572 & 1'h1;
  assign v_2572 = v_2573 & v_2574;
  assign v_2573 = ~act_2385;
  assign v_2574 = v_2575 | v_2579;
  assign v_2575 = v_2576 | v_2577;
  assign v_2576 = mux_2576(v_2174);
  assign v_2577 = mux_2577(v_2578);
  assign v_2578 = ~v_2174;
  assign v_2579 = ~v_2382;
  assign v_2580 = v_2581 | v_2582;
  assign v_2581 = mux_2581(v_2384);
  assign v_2582 = mux_2582(v_2571);
  assign v_2583 = v_2584 & 1'h1;
  assign v_2584 = v_2585 & v_2586;
  assign v_2585 = ~act_2173;
  assign v_2586 = v_2587 | v_2591;
  assign v_2587 = v_2588 | v_2589;
  assign v_2588 = mux_2588(v_1738);
  assign v_2589 = mux_2589(v_2590);
  assign v_2590 = ~v_1738;
  assign v_2591 = ~v_2170;
  assign v_2592 = v_2593 | v_2594;
  assign v_2593 = mux_2593(v_2172);
  assign v_2594 = mux_2594(v_2583);
  assign v_2595 = v_2596 & 1'h1;
  assign v_2596 = v_2597 & v_2598;
  assign v_2597 = ~act_1737;
  assign v_2598 = v_2599 | v_22337;
  assign v_2599 = v_2600 | v_22335;
  assign v_2600 = mux_2600(v_2601);
  assign v_2601 = v_1734 & v_2602;
  assign v_2602 = v_2603 & 1'h1;
  assign v_2603 = v_2604 | 1'h0;
  assign v_2604 = ~v_2605;
  assign v_2606 = v_2607 | v_2609;
  assign v_2607 = act_2608 & 1'h1;
  assign act_2608 = v_1731 | v_2601;
  assign v_2609 = v_2610 & 1'h1;
  assign v_2610 = v_2611 & v_2612;
  assign v_2611 = ~act_2608;
  assign v_2612 = v_2613 | v_22331;
  assign v_2613 = v_2614 | v_22329;
  assign v_2614 = mux_2614(v_2615);
  assign v_2615 = v_2616 & v_4382;
  assign v_2616 = v_2617 & v_2605;
  assign v_2617 = ~v_2618;
  assign v_2619 = v_2620 | v_4375;
  assign v_2620 = act_2621 & 1'h1;
  assign act_2621 = v_2622 | v_3492;
  assign v_2622 = v_2623 & v_3493;
  assign v_2623 = v_2624 & v_3502;
  assign v_2624 = ~v_2625;
  assign v_2626 = v_2627 | v_3486;
  assign v_2627 = act_2628 & 1'h1;
  assign act_2628 = v_2629 | v_3051;
  assign v_2629 = v_2630 & v_3052;
  assign v_2630 = v_2631 & v_3061;
  assign v_2631 = ~v_2632;
  assign v_2633 = v_2634 | v_3045;
  assign v_2634 = act_2635 & 1'h1;
  assign act_2635 = v_2636 | v_2834;
  assign v_2636 = v_2637 & v_2835;
  assign v_2637 = v_2638 & v_2844;
  assign v_2638 = ~v_2639;
  assign v_2640 = v_2641 | v_2828;
  assign v_2641 = act_2642 & 1'h1;
  assign act_2642 = v_2643 | v_2729;
  assign v_2643 = v_2644 & v_2730;
  assign v_2644 = v_2645 & v_2739;
  assign v_2645 = ~v_2646;
  assign v_2647 = v_2648 | v_2723;
  assign v_2648 = act_2649 & 1'h1;
  assign act_2649 = v_2650 | v_2680;
  assign v_2650 = v_2651 & v_2681;
  assign v_2651 = v_2652 & v_2690;
  assign v_2652 = ~v_2653;
  assign v_2654 = v_2655 | v_2674;
  assign v_2655 = act_2656 & 1'h1;
  assign act_2656 = v_2657 | v_2663;
  assign v_2657 = v_2658 & v_2664;
  assign v_2658 = v_2659 & vout_canPeek_2669;
  assign v_2659 = ~vout_canPeek_2660;
  pebbles_core
    pebbles_core_2660
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2661),
       .in0_consume_en(vin0_consume_en_2660),
       .out_canPeek(vout_canPeek_2660),
       .out_peek(vout_peek_2660));
  assign v_2661 = v_2662 | v_2667;
  assign v_2662 = mux_2662(v_2663);
  assign v_2663 = vout_canPeek_2660 & v_2664;
  assign v_2664 = v_2665 & 1'h1;
  assign v_2665 = v_2666 | 1'h0;
  assign v_2666 = ~v_2653;
  assign v_2667 = mux_2667(v_2668);
  assign v_2668 = ~v_2663;
  pebbles_core
    pebbles_core_2669
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2670),
       .in0_consume_en(vin0_consume_en_2669),
       .out_canPeek(vout_canPeek_2669),
       .out_peek(vout_peek_2669));
  assign v_2670 = v_2671 | v_2672;
  assign v_2671 = mux_2671(v_2657);
  assign v_2672 = mux_2672(v_2673);
  assign v_2673 = ~v_2657;
  assign v_2674 = v_2675 & 1'h1;
  assign v_2675 = v_2676 & v_2677;
  assign v_2676 = ~act_2656;
  assign v_2677 = v_2678 | v_2686;
  assign v_2678 = v_2679 | v_2684;
  assign v_2679 = mux_2679(v_2680);
  assign v_2680 = v_2653 & v_2681;
  assign v_2681 = v_2682 & 1'h1;
  assign v_2682 = v_2683 | 1'h0;
  assign v_2683 = ~v_2646;
  assign v_2684 = mux_2684(v_2685);
  assign v_2685 = ~v_2680;
  assign v_2686 = ~v_2653;
  assign v_2687 = v_2688 | v_2689;
  assign v_2688 = mux_2688(v_2655);
  assign v_2689 = mux_2689(v_2674);
  assign v_2691 = v_2692 | v_2711;
  assign v_2692 = act_2693 & 1'h1;
  assign act_2693 = v_2694 | v_2700;
  assign v_2694 = v_2695 & v_2701;
  assign v_2695 = v_2696 & vout_canPeek_2706;
  assign v_2696 = ~vout_canPeek_2697;
  pebbles_core
    pebbles_core_2697
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2698),
       .in0_consume_en(vin0_consume_en_2697),
       .out_canPeek(vout_canPeek_2697),
       .out_peek(vout_peek_2697));
  assign v_2698 = v_2699 | v_2704;
  assign v_2699 = mux_2699(v_2700);
  assign v_2700 = vout_canPeek_2697 & v_2701;
  assign v_2701 = v_2702 & 1'h1;
  assign v_2702 = v_2703 | 1'h0;
  assign v_2703 = ~v_2690;
  assign v_2704 = mux_2704(v_2705);
  assign v_2705 = ~v_2700;
  pebbles_core
    pebbles_core_2706
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2707),
       .in0_consume_en(vin0_consume_en_2706),
       .out_canPeek(vout_canPeek_2706),
       .out_peek(vout_peek_2706));
  assign v_2707 = v_2708 | v_2709;
  assign v_2708 = mux_2708(v_2694);
  assign v_2709 = mux_2709(v_2710);
  assign v_2710 = ~v_2694;
  assign v_2711 = v_2712 & 1'h1;
  assign v_2712 = v_2713 & v_2714;
  assign v_2713 = ~act_2693;
  assign v_2714 = v_2715 | v_2719;
  assign v_2715 = v_2716 | v_2717;
  assign v_2716 = mux_2716(v_2650);
  assign v_2717 = mux_2717(v_2718);
  assign v_2718 = ~v_2650;
  assign v_2719 = ~v_2690;
  assign v_2720 = v_2721 | v_2722;
  assign v_2721 = mux_2721(v_2692);
  assign v_2722 = mux_2722(v_2711);
  assign v_2723 = v_2724 & 1'h1;
  assign v_2724 = v_2725 & v_2726;
  assign v_2725 = ~act_2649;
  assign v_2726 = v_2727 | v_2735;
  assign v_2727 = v_2728 | v_2733;
  assign v_2728 = mux_2728(v_2729);
  assign v_2729 = v_2646 & v_2730;
  assign v_2730 = v_2731 & 1'h1;
  assign v_2731 = v_2732 | 1'h0;
  assign v_2732 = ~v_2639;
  assign v_2733 = mux_2733(v_2734);
  assign v_2734 = ~v_2729;
  assign v_2735 = ~v_2646;
  assign v_2736 = v_2737 | v_2738;
  assign v_2737 = mux_2737(v_2648);
  assign v_2738 = mux_2738(v_2723);
  assign v_2740 = v_2741 | v_2816;
  assign v_2741 = act_2742 & 1'h1;
  assign act_2742 = v_2743 | v_2773;
  assign v_2743 = v_2744 & v_2774;
  assign v_2744 = v_2745 & v_2783;
  assign v_2745 = ~v_2746;
  assign v_2747 = v_2748 | v_2767;
  assign v_2748 = act_2749 & 1'h1;
  assign act_2749 = v_2750 | v_2756;
  assign v_2750 = v_2751 & v_2757;
  assign v_2751 = v_2752 & vout_canPeek_2762;
  assign v_2752 = ~vout_canPeek_2753;
  pebbles_core
    pebbles_core_2753
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2754),
       .in0_consume_en(vin0_consume_en_2753),
       .out_canPeek(vout_canPeek_2753),
       .out_peek(vout_peek_2753));
  assign v_2754 = v_2755 | v_2760;
  assign v_2755 = mux_2755(v_2756);
  assign v_2756 = vout_canPeek_2753 & v_2757;
  assign v_2757 = v_2758 & 1'h1;
  assign v_2758 = v_2759 | 1'h0;
  assign v_2759 = ~v_2746;
  assign v_2760 = mux_2760(v_2761);
  assign v_2761 = ~v_2756;
  pebbles_core
    pebbles_core_2762
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2763),
       .in0_consume_en(vin0_consume_en_2762),
       .out_canPeek(vout_canPeek_2762),
       .out_peek(vout_peek_2762));
  assign v_2763 = v_2764 | v_2765;
  assign v_2764 = mux_2764(v_2750);
  assign v_2765 = mux_2765(v_2766);
  assign v_2766 = ~v_2750;
  assign v_2767 = v_2768 & 1'h1;
  assign v_2768 = v_2769 & v_2770;
  assign v_2769 = ~act_2749;
  assign v_2770 = v_2771 | v_2779;
  assign v_2771 = v_2772 | v_2777;
  assign v_2772 = mux_2772(v_2773);
  assign v_2773 = v_2746 & v_2774;
  assign v_2774 = v_2775 & 1'h1;
  assign v_2775 = v_2776 | 1'h0;
  assign v_2776 = ~v_2739;
  assign v_2777 = mux_2777(v_2778);
  assign v_2778 = ~v_2773;
  assign v_2779 = ~v_2746;
  assign v_2780 = v_2781 | v_2782;
  assign v_2781 = mux_2781(v_2748);
  assign v_2782 = mux_2782(v_2767);
  assign v_2784 = v_2785 | v_2804;
  assign v_2785 = act_2786 & 1'h1;
  assign act_2786 = v_2787 | v_2793;
  assign v_2787 = v_2788 & v_2794;
  assign v_2788 = v_2789 & vout_canPeek_2799;
  assign v_2789 = ~vout_canPeek_2790;
  pebbles_core
    pebbles_core_2790
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2791),
       .in0_consume_en(vin0_consume_en_2790),
       .out_canPeek(vout_canPeek_2790),
       .out_peek(vout_peek_2790));
  assign v_2791 = v_2792 | v_2797;
  assign v_2792 = mux_2792(v_2793);
  assign v_2793 = vout_canPeek_2790 & v_2794;
  assign v_2794 = v_2795 & 1'h1;
  assign v_2795 = v_2796 | 1'h0;
  assign v_2796 = ~v_2783;
  assign v_2797 = mux_2797(v_2798);
  assign v_2798 = ~v_2793;
  pebbles_core
    pebbles_core_2799
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2800),
       .in0_consume_en(vin0_consume_en_2799),
       .out_canPeek(vout_canPeek_2799),
       .out_peek(vout_peek_2799));
  assign v_2800 = v_2801 | v_2802;
  assign v_2801 = mux_2801(v_2787);
  assign v_2802 = mux_2802(v_2803);
  assign v_2803 = ~v_2787;
  assign v_2804 = v_2805 & 1'h1;
  assign v_2805 = v_2806 & v_2807;
  assign v_2806 = ~act_2786;
  assign v_2807 = v_2808 | v_2812;
  assign v_2808 = v_2809 | v_2810;
  assign v_2809 = mux_2809(v_2743);
  assign v_2810 = mux_2810(v_2811);
  assign v_2811 = ~v_2743;
  assign v_2812 = ~v_2783;
  assign v_2813 = v_2814 | v_2815;
  assign v_2814 = mux_2814(v_2785);
  assign v_2815 = mux_2815(v_2804);
  assign v_2816 = v_2817 & 1'h1;
  assign v_2817 = v_2818 & v_2819;
  assign v_2818 = ~act_2742;
  assign v_2819 = v_2820 | v_2824;
  assign v_2820 = v_2821 | v_2822;
  assign v_2821 = mux_2821(v_2643);
  assign v_2822 = mux_2822(v_2823);
  assign v_2823 = ~v_2643;
  assign v_2824 = ~v_2739;
  assign v_2825 = v_2826 | v_2827;
  assign v_2826 = mux_2826(v_2741);
  assign v_2827 = mux_2827(v_2816);
  assign v_2828 = v_2829 & 1'h1;
  assign v_2829 = v_2830 & v_2831;
  assign v_2830 = ~act_2642;
  assign v_2831 = v_2832 | v_2840;
  assign v_2832 = v_2833 | v_2838;
  assign v_2833 = mux_2833(v_2834);
  assign v_2834 = v_2639 & v_2835;
  assign v_2835 = v_2836 & 1'h1;
  assign v_2836 = v_2837 | 1'h0;
  assign v_2837 = ~v_2632;
  assign v_2838 = mux_2838(v_2839);
  assign v_2839 = ~v_2834;
  assign v_2840 = ~v_2639;
  assign v_2841 = v_2842 | v_2843;
  assign v_2842 = mux_2842(v_2641);
  assign v_2843 = mux_2843(v_2828);
  assign v_2845 = v_2846 | v_3033;
  assign v_2846 = act_2847 & 1'h1;
  assign act_2847 = v_2848 | v_2934;
  assign v_2848 = v_2849 & v_2935;
  assign v_2849 = v_2850 & v_2944;
  assign v_2850 = ~v_2851;
  assign v_2852 = v_2853 | v_2928;
  assign v_2853 = act_2854 & 1'h1;
  assign act_2854 = v_2855 | v_2885;
  assign v_2855 = v_2856 & v_2886;
  assign v_2856 = v_2857 & v_2895;
  assign v_2857 = ~v_2858;
  assign v_2859 = v_2860 | v_2879;
  assign v_2860 = act_2861 & 1'h1;
  assign act_2861 = v_2862 | v_2868;
  assign v_2862 = v_2863 & v_2869;
  assign v_2863 = v_2864 & vout_canPeek_2874;
  assign v_2864 = ~vout_canPeek_2865;
  pebbles_core
    pebbles_core_2865
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2866),
       .in0_consume_en(vin0_consume_en_2865),
       .out_canPeek(vout_canPeek_2865),
       .out_peek(vout_peek_2865));
  assign v_2866 = v_2867 | v_2872;
  assign v_2867 = mux_2867(v_2868);
  assign v_2868 = vout_canPeek_2865 & v_2869;
  assign v_2869 = v_2870 & 1'h1;
  assign v_2870 = v_2871 | 1'h0;
  assign v_2871 = ~v_2858;
  assign v_2872 = mux_2872(v_2873);
  assign v_2873 = ~v_2868;
  pebbles_core
    pebbles_core_2874
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2875),
       .in0_consume_en(vin0_consume_en_2874),
       .out_canPeek(vout_canPeek_2874),
       .out_peek(vout_peek_2874));
  assign v_2875 = v_2876 | v_2877;
  assign v_2876 = mux_2876(v_2862);
  assign v_2877 = mux_2877(v_2878);
  assign v_2878 = ~v_2862;
  assign v_2879 = v_2880 & 1'h1;
  assign v_2880 = v_2881 & v_2882;
  assign v_2881 = ~act_2861;
  assign v_2882 = v_2883 | v_2891;
  assign v_2883 = v_2884 | v_2889;
  assign v_2884 = mux_2884(v_2885);
  assign v_2885 = v_2858 & v_2886;
  assign v_2886 = v_2887 & 1'h1;
  assign v_2887 = v_2888 | 1'h0;
  assign v_2888 = ~v_2851;
  assign v_2889 = mux_2889(v_2890);
  assign v_2890 = ~v_2885;
  assign v_2891 = ~v_2858;
  assign v_2892 = v_2893 | v_2894;
  assign v_2893 = mux_2893(v_2860);
  assign v_2894 = mux_2894(v_2879);
  assign v_2896 = v_2897 | v_2916;
  assign v_2897 = act_2898 & 1'h1;
  assign act_2898 = v_2899 | v_2905;
  assign v_2899 = v_2900 & v_2906;
  assign v_2900 = v_2901 & vout_canPeek_2911;
  assign v_2901 = ~vout_canPeek_2902;
  pebbles_core
    pebbles_core_2902
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2903),
       .in0_consume_en(vin0_consume_en_2902),
       .out_canPeek(vout_canPeek_2902),
       .out_peek(vout_peek_2902));
  assign v_2903 = v_2904 | v_2909;
  assign v_2904 = mux_2904(v_2905);
  assign v_2905 = vout_canPeek_2902 & v_2906;
  assign v_2906 = v_2907 & 1'h1;
  assign v_2907 = v_2908 | 1'h0;
  assign v_2908 = ~v_2895;
  assign v_2909 = mux_2909(v_2910);
  assign v_2910 = ~v_2905;
  pebbles_core
    pebbles_core_2911
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2912),
       .in0_consume_en(vin0_consume_en_2911),
       .out_canPeek(vout_canPeek_2911),
       .out_peek(vout_peek_2911));
  assign v_2912 = v_2913 | v_2914;
  assign v_2913 = mux_2913(v_2899);
  assign v_2914 = mux_2914(v_2915);
  assign v_2915 = ~v_2899;
  assign v_2916 = v_2917 & 1'h1;
  assign v_2917 = v_2918 & v_2919;
  assign v_2918 = ~act_2898;
  assign v_2919 = v_2920 | v_2924;
  assign v_2920 = v_2921 | v_2922;
  assign v_2921 = mux_2921(v_2855);
  assign v_2922 = mux_2922(v_2923);
  assign v_2923 = ~v_2855;
  assign v_2924 = ~v_2895;
  assign v_2925 = v_2926 | v_2927;
  assign v_2926 = mux_2926(v_2897);
  assign v_2927 = mux_2927(v_2916);
  assign v_2928 = v_2929 & 1'h1;
  assign v_2929 = v_2930 & v_2931;
  assign v_2930 = ~act_2854;
  assign v_2931 = v_2932 | v_2940;
  assign v_2932 = v_2933 | v_2938;
  assign v_2933 = mux_2933(v_2934);
  assign v_2934 = v_2851 & v_2935;
  assign v_2935 = v_2936 & 1'h1;
  assign v_2936 = v_2937 | 1'h0;
  assign v_2937 = ~v_2844;
  assign v_2938 = mux_2938(v_2939);
  assign v_2939 = ~v_2934;
  assign v_2940 = ~v_2851;
  assign v_2941 = v_2942 | v_2943;
  assign v_2942 = mux_2942(v_2853);
  assign v_2943 = mux_2943(v_2928);
  assign v_2945 = v_2946 | v_3021;
  assign v_2946 = act_2947 & 1'h1;
  assign act_2947 = v_2948 | v_2978;
  assign v_2948 = v_2949 & v_2979;
  assign v_2949 = v_2950 & v_2988;
  assign v_2950 = ~v_2951;
  assign v_2952 = v_2953 | v_2972;
  assign v_2953 = act_2954 & 1'h1;
  assign act_2954 = v_2955 | v_2961;
  assign v_2955 = v_2956 & v_2962;
  assign v_2956 = v_2957 & vout_canPeek_2967;
  assign v_2957 = ~vout_canPeek_2958;
  pebbles_core
    pebbles_core_2958
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2959),
       .in0_consume_en(vin0_consume_en_2958),
       .out_canPeek(vout_canPeek_2958),
       .out_peek(vout_peek_2958));
  assign v_2959 = v_2960 | v_2965;
  assign v_2960 = mux_2960(v_2961);
  assign v_2961 = vout_canPeek_2958 & v_2962;
  assign v_2962 = v_2963 & 1'h1;
  assign v_2963 = v_2964 | 1'h0;
  assign v_2964 = ~v_2951;
  assign v_2965 = mux_2965(v_2966);
  assign v_2966 = ~v_2961;
  pebbles_core
    pebbles_core_2967
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2968),
       .in0_consume_en(vin0_consume_en_2967),
       .out_canPeek(vout_canPeek_2967),
       .out_peek(vout_peek_2967));
  assign v_2968 = v_2969 | v_2970;
  assign v_2969 = mux_2969(v_2955);
  assign v_2970 = mux_2970(v_2971);
  assign v_2971 = ~v_2955;
  assign v_2972 = v_2973 & 1'h1;
  assign v_2973 = v_2974 & v_2975;
  assign v_2974 = ~act_2954;
  assign v_2975 = v_2976 | v_2984;
  assign v_2976 = v_2977 | v_2982;
  assign v_2977 = mux_2977(v_2978);
  assign v_2978 = v_2951 & v_2979;
  assign v_2979 = v_2980 & 1'h1;
  assign v_2980 = v_2981 | 1'h0;
  assign v_2981 = ~v_2944;
  assign v_2982 = mux_2982(v_2983);
  assign v_2983 = ~v_2978;
  assign v_2984 = ~v_2951;
  assign v_2985 = v_2986 | v_2987;
  assign v_2986 = mux_2986(v_2953);
  assign v_2987 = mux_2987(v_2972);
  assign v_2989 = v_2990 | v_3009;
  assign v_2990 = act_2991 & 1'h1;
  assign act_2991 = v_2992 | v_2998;
  assign v_2992 = v_2993 & v_2999;
  assign v_2993 = v_2994 & vout_canPeek_3004;
  assign v_2994 = ~vout_canPeek_2995;
  pebbles_core
    pebbles_core_2995
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2996),
       .in0_consume_en(vin0_consume_en_2995),
       .out_canPeek(vout_canPeek_2995),
       .out_peek(vout_peek_2995));
  assign v_2996 = v_2997 | v_3002;
  assign v_2997 = mux_2997(v_2998);
  assign v_2998 = vout_canPeek_2995 & v_2999;
  assign v_2999 = v_3000 & 1'h1;
  assign v_3000 = v_3001 | 1'h0;
  assign v_3001 = ~v_2988;
  assign v_3002 = mux_3002(v_3003);
  assign v_3003 = ~v_2998;
  pebbles_core
    pebbles_core_3004
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3005),
       .in0_consume_en(vin0_consume_en_3004),
       .out_canPeek(vout_canPeek_3004),
       .out_peek(vout_peek_3004));
  assign v_3005 = v_3006 | v_3007;
  assign v_3006 = mux_3006(v_2992);
  assign v_3007 = mux_3007(v_3008);
  assign v_3008 = ~v_2992;
  assign v_3009 = v_3010 & 1'h1;
  assign v_3010 = v_3011 & v_3012;
  assign v_3011 = ~act_2991;
  assign v_3012 = v_3013 | v_3017;
  assign v_3013 = v_3014 | v_3015;
  assign v_3014 = mux_3014(v_2948);
  assign v_3015 = mux_3015(v_3016);
  assign v_3016 = ~v_2948;
  assign v_3017 = ~v_2988;
  assign v_3018 = v_3019 | v_3020;
  assign v_3019 = mux_3019(v_2990);
  assign v_3020 = mux_3020(v_3009);
  assign v_3021 = v_3022 & 1'h1;
  assign v_3022 = v_3023 & v_3024;
  assign v_3023 = ~act_2947;
  assign v_3024 = v_3025 | v_3029;
  assign v_3025 = v_3026 | v_3027;
  assign v_3026 = mux_3026(v_2848);
  assign v_3027 = mux_3027(v_3028);
  assign v_3028 = ~v_2848;
  assign v_3029 = ~v_2944;
  assign v_3030 = v_3031 | v_3032;
  assign v_3031 = mux_3031(v_2946);
  assign v_3032 = mux_3032(v_3021);
  assign v_3033 = v_3034 & 1'h1;
  assign v_3034 = v_3035 & v_3036;
  assign v_3035 = ~act_2847;
  assign v_3036 = v_3037 | v_3041;
  assign v_3037 = v_3038 | v_3039;
  assign v_3038 = mux_3038(v_2636);
  assign v_3039 = mux_3039(v_3040);
  assign v_3040 = ~v_2636;
  assign v_3041 = ~v_2844;
  assign v_3042 = v_3043 | v_3044;
  assign v_3043 = mux_3043(v_2846);
  assign v_3044 = mux_3044(v_3033);
  assign v_3045 = v_3046 & 1'h1;
  assign v_3046 = v_3047 & v_3048;
  assign v_3047 = ~act_2635;
  assign v_3048 = v_3049 | v_3057;
  assign v_3049 = v_3050 | v_3055;
  assign v_3050 = mux_3050(v_3051);
  assign v_3051 = v_2632 & v_3052;
  assign v_3052 = v_3053 & 1'h1;
  assign v_3053 = v_3054 | 1'h0;
  assign v_3054 = ~v_2625;
  assign v_3055 = mux_3055(v_3056);
  assign v_3056 = ~v_3051;
  assign v_3057 = ~v_2632;
  assign v_3058 = v_3059 | v_3060;
  assign v_3059 = mux_3059(v_2634);
  assign v_3060 = mux_3060(v_3045);
  assign v_3062 = v_3063 | v_3474;
  assign v_3063 = act_3064 & 1'h1;
  assign act_3064 = v_3065 | v_3263;
  assign v_3065 = v_3066 & v_3264;
  assign v_3066 = v_3067 & v_3273;
  assign v_3067 = ~v_3068;
  assign v_3069 = v_3070 | v_3257;
  assign v_3070 = act_3071 & 1'h1;
  assign act_3071 = v_3072 | v_3158;
  assign v_3072 = v_3073 & v_3159;
  assign v_3073 = v_3074 & v_3168;
  assign v_3074 = ~v_3075;
  assign v_3076 = v_3077 | v_3152;
  assign v_3077 = act_3078 & 1'h1;
  assign act_3078 = v_3079 | v_3109;
  assign v_3079 = v_3080 & v_3110;
  assign v_3080 = v_3081 & v_3119;
  assign v_3081 = ~v_3082;
  assign v_3083 = v_3084 | v_3103;
  assign v_3084 = act_3085 & 1'h1;
  assign act_3085 = v_3086 | v_3092;
  assign v_3086 = v_3087 & v_3093;
  assign v_3087 = v_3088 & vout_canPeek_3098;
  assign v_3088 = ~vout_canPeek_3089;
  pebbles_core
    pebbles_core_3089
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3090),
       .in0_consume_en(vin0_consume_en_3089),
       .out_canPeek(vout_canPeek_3089),
       .out_peek(vout_peek_3089));
  assign v_3090 = v_3091 | v_3096;
  assign v_3091 = mux_3091(v_3092);
  assign v_3092 = vout_canPeek_3089 & v_3093;
  assign v_3093 = v_3094 & 1'h1;
  assign v_3094 = v_3095 | 1'h0;
  assign v_3095 = ~v_3082;
  assign v_3096 = mux_3096(v_3097);
  assign v_3097 = ~v_3092;
  pebbles_core
    pebbles_core_3098
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3099),
       .in0_consume_en(vin0_consume_en_3098),
       .out_canPeek(vout_canPeek_3098),
       .out_peek(vout_peek_3098));
  assign v_3099 = v_3100 | v_3101;
  assign v_3100 = mux_3100(v_3086);
  assign v_3101 = mux_3101(v_3102);
  assign v_3102 = ~v_3086;
  assign v_3103 = v_3104 & 1'h1;
  assign v_3104 = v_3105 & v_3106;
  assign v_3105 = ~act_3085;
  assign v_3106 = v_3107 | v_3115;
  assign v_3107 = v_3108 | v_3113;
  assign v_3108 = mux_3108(v_3109);
  assign v_3109 = v_3082 & v_3110;
  assign v_3110 = v_3111 & 1'h1;
  assign v_3111 = v_3112 | 1'h0;
  assign v_3112 = ~v_3075;
  assign v_3113 = mux_3113(v_3114);
  assign v_3114 = ~v_3109;
  assign v_3115 = ~v_3082;
  assign v_3116 = v_3117 | v_3118;
  assign v_3117 = mux_3117(v_3084);
  assign v_3118 = mux_3118(v_3103);
  assign v_3120 = v_3121 | v_3140;
  assign v_3121 = act_3122 & 1'h1;
  assign act_3122 = v_3123 | v_3129;
  assign v_3123 = v_3124 & v_3130;
  assign v_3124 = v_3125 & vout_canPeek_3135;
  assign v_3125 = ~vout_canPeek_3126;
  pebbles_core
    pebbles_core_3126
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3127),
       .in0_consume_en(vin0_consume_en_3126),
       .out_canPeek(vout_canPeek_3126),
       .out_peek(vout_peek_3126));
  assign v_3127 = v_3128 | v_3133;
  assign v_3128 = mux_3128(v_3129);
  assign v_3129 = vout_canPeek_3126 & v_3130;
  assign v_3130 = v_3131 & 1'h1;
  assign v_3131 = v_3132 | 1'h0;
  assign v_3132 = ~v_3119;
  assign v_3133 = mux_3133(v_3134);
  assign v_3134 = ~v_3129;
  pebbles_core
    pebbles_core_3135
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3136),
       .in0_consume_en(vin0_consume_en_3135),
       .out_canPeek(vout_canPeek_3135),
       .out_peek(vout_peek_3135));
  assign v_3136 = v_3137 | v_3138;
  assign v_3137 = mux_3137(v_3123);
  assign v_3138 = mux_3138(v_3139);
  assign v_3139 = ~v_3123;
  assign v_3140 = v_3141 & 1'h1;
  assign v_3141 = v_3142 & v_3143;
  assign v_3142 = ~act_3122;
  assign v_3143 = v_3144 | v_3148;
  assign v_3144 = v_3145 | v_3146;
  assign v_3145 = mux_3145(v_3079);
  assign v_3146 = mux_3146(v_3147);
  assign v_3147 = ~v_3079;
  assign v_3148 = ~v_3119;
  assign v_3149 = v_3150 | v_3151;
  assign v_3150 = mux_3150(v_3121);
  assign v_3151 = mux_3151(v_3140);
  assign v_3152 = v_3153 & 1'h1;
  assign v_3153 = v_3154 & v_3155;
  assign v_3154 = ~act_3078;
  assign v_3155 = v_3156 | v_3164;
  assign v_3156 = v_3157 | v_3162;
  assign v_3157 = mux_3157(v_3158);
  assign v_3158 = v_3075 & v_3159;
  assign v_3159 = v_3160 & 1'h1;
  assign v_3160 = v_3161 | 1'h0;
  assign v_3161 = ~v_3068;
  assign v_3162 = mux_3162(v_3163);
  assign v_3163 = ~v_3158;
  assign v_3164 = ~v_3075;
  assign v_3165 = v_3166 | v_3167;
  assign v_3166 = mux_3166(v_3077);
  assign v_3167 = mux_3167(v_3152);
  assign v_3169 = v_3170 | v_3245;
  assign v_3170 = act_3171 & 1'h1;
  assign act_3171 = v_3172 | v_3202;
  assign v_3172 = v_3173 & v_3203;
  assign v_3173 = v_3174 & v_3212;
  assign v_3174 = ~v_3175;
  assign v_3176 = v_3177 | v_3196;
  assign v_3177 = act_3178 & 1'h1;
  assign act_3178 = v_3179 | v_3185;
  assign v_3179 = v_3180 & v_3186;
  assign v_3180 = v_3181 & vout_canPeek_3191;
  assign v_3181 = ~vout_canPeek_3182;
  pebbles_core
    pebbles_core_3182
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3183),
       .in0_consume_en(vin0_consume_en_3182),
       .out_canPeek(vout_canPeek_3182),
       .out_peek(vout_peek_3182));
  assign v_3183 = v_3184 | v_3189;
  assign v_3184 = mux_3184(v_3185);
  assign v_3185 = vout_canPeek_3182 & v_3186;
  assign v_3186 = v_3187 & 1'h1;
  assign v_3187 = v_3188 | 1'h0;
  assign v_3188 = ~v_3175;
  assign v_3189 = mux_3189(v_3190);
  assign v_3190 = ~v_3185;
  pebbles_core
    pebbles_core_3191
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3192),
       .in0_consume_en(vin0_consume_en_3191),
       .out_canPeek(vout_canPeek_3191),
       .out_peek(vout_peek_3191));
  assign v_3192 = v_3193 | v_3194;
  assign v_3193 = mux_3193(v_3179);
  assign v_3194 = mux_3194(v_3195);
  assign v_3195 = ~v_3179;
  assign v_3196 = v_3197 & 1'h1;
  assign v_3197 = v_3198 & v_3199;
  assign v_3198 = ~act_3178;
  assign v_3199 = v_3200 | v_3208;
  assign v_3200 = v_3201 | v_3206;
  assign v_3201 = mux_3201(v_3202);
  assign v_3202 = v_3175 & v_3203;
  assign v_3203 = v_3204 & 1'h1;
  assign v_3204 = v_3205 | 1'h0;
  assign v_3205 = ~v_3168;
  assign v_3206 = mux_3206(v_3207);
  assign v_3207 = ~v_3202;
  assign v_3208 = ~v_3175;
  assign v_3209 = v_3210 | v_3211;
  assign v_3210 = mux_3210(v_3177);
  assign v_3211 = mux_3211(v_3196);
  assign v_3213 = v_3214 | v_3233;
  assign v_3214 = act_3215 & 1'h1;
  assign act_3215 = v_3216 | v_3222;
  assign v_3216 = v_3217 & v_3223;
  assign v_3217 = v_3218 & vout_canPeek_3228;
  assign v_3218 = ~vout_canPeek_3219;
  pebbles_core
    pebbles_core_3219
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3220),
       .in0_consume_en(vin0_consume_en_3219),
       .out_canPeek(vout_canPeek_3219),
       .out_peek(vout_peek_3219));
  assign v_3220 = v_3221 | v_3226;
  assign v_3221 = mux_3221(v_3222);
  assign v_3222 = vout_canPeek_3219 & v_3223;
  assign v_3223 = v_3224 & 1'h1;
  assign v_3224 = v_3225 | 1'h0;
  assign v_3225 = ~v_3212;
  assign v_3226 = mux_3226(v_3227);
  assign v_3227 = ~v_3222;
  pebbles_core
    pebbles_core_3228
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3229),
       .in0_consume_en(vin0_consume_en_3228),
       .out_canPeek(vout_canPeek_3228),
       .out_peek(vout_peek_3228));
  assign v_3229 = v_3230 | v_3231;
  assign v_3230 = mux_3230(v_3216);
  assign v_3231 = mux_3231(v_3232);
  assign v_3232 = ~v_3216;
  assign v_3233 = v_3234 & 1'h1;
  assign v_3234 = v_3235 & v_3236;
  assign v_3235 = ~act_3215;
  assign v_3236 = v_3237 | v_3241;
  assign v_3237 = v_3238 | v_3239;
  assign v_3238 = mux_3238(v_3172);
  assign v_3239 = mux_3239(v_3240);
  assign v_3240 = ~v_3172;
  assign v_3241 = ~v_3212;
  assign v_3242 = v_3243 | v_3244;
  assign v_3243 = mux_3243(v_3214);
  assign v_3244 = mux_3244(v_3233);
  assign v_3245 = v_3246 & 1'h1;
  assign v_3246 = v_3247 & v_3248;
  assign v_3247 = ~act_3171;
  assign v_3248 = v_3249 | v_3253;
  assign v_3249 = v_3250 | v_3251;
  assign v_3250 = mux_3250(v_3072);
  assign v_3251 = mux_3251(v_3252);
  assign v_3252 = ~v_3072;
  assign v_3253 = ~v_3168;
  assign v_3254 = v_3255 | v_3256;
  assign v_3255 = mux_3255(v_3170);
  assign v_3256 = mux_3256(v_3245);
  assign v_3257 = v_3258 & 1'h1;
  assign v_3258 = v_3259 & v_3260;
  assign v_3259 = ~act_3071;
  assign v_3260 = v_3261 | v_3269;
  assign v_3261 = v_3262 | v_3267;
  assign v_3262 = mux_3262(v_3263);
  assign v_3263 = v_3068 & v_3264;
  assign v_3264 = v_3265 & 1'h1;
  assign v_3265 = v_3266 | 1'h0;
  assign v_3266 = ~v_3061;
  assign v_3267 = mux_3267(v_3268);
  assign v_3268 = ~v_3263;
  assign v_3269 = ~v_3068;
  assign v_3270 = v_3271 | v_3272;
  assign v_3271 = mux_3271(v_3070);
  assign v_3272 = mux_3272(v_3257);
  assign v_3274 = v_3275 | v_3462;
  assign v_3275 = act_3276 & 1'h1;
  assign act_3276 = v_3277 | v_3363;
  assign v_3277 = v_3278 & v_3364;
  assign v_3278 = v_3279 & v_3373;
  assign v_3279 = ~v_3280;
  assign v_3281 = v_3282 | v_3357;
  assign v_3282 = act_3283 & 1'h1;
  assign act_3283 = v_3284 | v_3314;
  assign v_3284 = v_3285 & v_3315;
  assign v_3285 = v_3286 & v_3324;
  assign v_3286 = ~v_3287;
  assign v_3288 = v_3289 | v_3308;
  assign v_3289 = act_3290 & 1'h1;
  assign act_3290 = v_3291 | v_3297;
  assign v_3291 = v_3292 & v_3298;
  assign v_3292 = v_3293 & vout_canPeek_3303;
  assign v_3293 = ~vout_canPeek_3294;
  pebbles_core
    pebbles_core_3294
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3295),
       .in0_consume_en(vin0_consume_en_3294),
       .out_canPeek(vout_canPeek_3294),
       .out_peek(vout_peek_3294));
  assign v_3295 = v_3296 | v_3301;
  assign v_3296 = mux_3296(v_3297);
  assign v_3297 = vout_canPeek_3294 & v_3298;
  assign v_3298 = v_3299 & 1'h1;
  assign v_3299 = v_3300 | 1'h0;
  assign v_3300 = ~v_3287;
  assign v_3301 = mux_3301(v_3302);
  assign v_3302 = ~v_3297;
  pebbles_core
    pebbles_core_3303
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3304),
       .in0_consume_en(vin0_consume_en_3303),
       .out_canPeek(vout_canPeek_3303),
       .out_peek(vout_peek_3303));
  assign v_3304 = v_3305 | v_3306;
  assign v_3305 = mux_3305(v_3291);
  assign v_3306 = mux_3306(v_3307);
  assign v_3307 = ~v_3291;
  assign v_3308 = v_3309 & 1'h1;
  assign v_3309 = v_3310 & v_3311;
  assign v_3310 = ~act_3290;
  assign v_3311 = v_3312 | v_3320;
  assign v_3312 = v_3313 | v_3318;
  assign v_3313 = mux_3313(v_3314);
  assign v_3314 = v_3287 & v_3315;
  assign v_3315 = v_3316 & 1'h1;
  assign v_3316 = v_3317 | 1'h0;
  assign v_3317 = ~v_3280;
  assign v_3318 = mux_3318(v_3319);
  assign v_3319 = ~v_3314;
  assign v_3320 = ~v_3287;
  assign v_3321 = v_3322 | v_3323;
  assign v_3322 = mux_3322(v_3289);
  assign v_3323 = mux_3323(v_3308);
  assign v_3325 = v_3326 | v_3345;
  assign v_3326 = act_3327 & 1'h1;
  assign act_3327 = v_3328 | v_3334;
  assign v_3328 = v_3329 & v_3335;
  assign v_3329 = v_3330 & vout_canPeek_3340;
  assign v_3330 = ~vout_canPeek_3331;
  pebbles_core
    pebbles_core_3331
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3332),
       .in0_consume_en(vin0_consume_en_3331),
       .out_canPeek(vout_canPeek_3331),
       .out_peek(vout_peek_3331));
  assign v_3332 = v_3333 | v_3338;
  assign v_3333 = mux_3333(v_3334);
  assign v_3334 = vout_canPeek_3331 & v_3335;
  assign v_3335 = v_3336 & 1'h1;
  assign v_3336 = v_3337 | 1'h0;
  assign v_3337 = ~v_3324;
  assign v_3338 = mux_3338(v_3339);
  assign v_3339 = ~v_3334;
  pebbles_core
    pebbles_core_3340
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3341),
       .in0_consume_en(vin0_consume_en_3340),
       .out_canPeek(vout_canPeek_3340),
       .out_peek(vout_peek_3340));
  assign v_3341 = v_3342 | v_3343;
  assign v_3342 = mux_3342(v_3328);
  assign v_3343 = mux_3343(v_3344);
  assign v_3344 = ~v_3328;
  assign v_3345 = v_3346 & 1'h1;
  assign v_3346 = v_3347 & v_3348;
  assign v_3347 = ~act_3327;
  assign v_3348 = v_3349 | v_3353;
  assign v_3349 = v_3350 | v_3351;
  assign v_3350 = mux_3350(v_3284);
  assign v_3351 = mux_3351(v_3352);
  assign v_3352 = ~v_3284;
  assign v_3353 = ~v_3324;
  assign v_3354 = v_3355 | v_3356;
  assign v_3355 = mux_3355(v_3326);
  assign v_3356 = mux_3356(v_3345);
  assign v_3357 = v_3358 & 1'h1;
  assign v_3358 = v_3359 & v_3360;
  assign v_3359 = ~act_3283;
  assign v_3360 = v_3361 | v_3369;
  assign v_3361 = v_3362 | v_3367;
  assign v_3362 = mux_3362(v_3363);
  assign v_3363 = v_3280 & v_3364;
  assign v_3364 = v_3365 & 1'h1;
  assign v_3365 = v_3366 | 1'h0;
  assign v_3366 = ~v_3273;
  assign v_3367 = mux_3367(v_3368);
  assign v_3368 = ~v_3363;
  assign v_3369 = ~v_3280;
  assign v_3370 = v_3371 | v_3372;
  assign v_3371 = mux_3371(v_3282);
  assign v_3372 = mux_3372(v_3357);
  assign v_3374 = v_3375 | v_3450;
  assign v_3375 = act_3376 & 1'h1;
  assign act_3376 = v_3377 | v_3407;
  assign v_3377 = v_3378 & v_3408;
  assign v_3378 = v_3379 & v_3417;
  assign v_3379 = ~v_3380;
  assign v_3381 = v_3382 | v_3401;
  assign v_3382 = act_3383 & 1'h1;
  assign act_3383 = v_3384 | v_3390;
  assign v_3384 = v_3385 & v_3391;
  assign v_3385 = v_3386 & vout_canPeek_3396;
  assign v_3386 = ~vout_canPeek_3387;
  pebbles_core
    pebbles_core_3387
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3388),
       .in0_consume_en(vin0_consume_en_3387),
       .out_canPeek(vout_canPeek_3387),
       .out_peek(vout_peek_3387));
  assign v_3388 = v_3389 | v_3394;
  assign v_3389 = mux_3389(v_3390);
  assign v_3390 = vout_canPeek_3387 & v_3391;
  assign v_3391 = v_3392 & 1'h1;
  assign v_3392 = v_3393 | 1'h0;
  assign v_3393 = ~v_3380;
  assign v_3394 = mux_3394(v_3395);
  assign v_3395 = ~v_3390;
  pebbles_core
    pebbles_core_3396
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3397),
       .in0_consume_en(vin0_consume_en_3396),
       .out_canPeek(vout_canPeek_3396),
       .out_peek(vout_peek_3396));
  assign v_3397 = v_3398 | v_3399;
  assign v_3398 = mux_3398(v_3384);
  assign v_3399 = mux_3399(v_3400);
  assign v_3400 = ~v_3384;
  assign v_3401 = v_3402 & 1'h1;
  assign v_3402 = v_3403 & v_3404;
  assign v_3403 = ~act_3383;
  assign v_3404 = v_3405 | v_3413;
  assign v_3405 = v_3406 | v_3411;
  assign v_3406 = mux_3406(v_3407);
  assign v_3407 = v_3380 & v_3408;
  assign v_3408 = v_3409 & 1'h1;
  assign v_3409 = v_3410 | 1'h0;
  assign v_3410 = ~v_3373;
  assign v_3411 = mux_3411(v_3412);
  assign v_3412 = ~v_3407;
  assign v_3413 = ~v_3380;
  assign v_3414 = v_3415 | v_3416;
  assign v_3415 = mux_3415(v_3382);
  assign v_3416 = mux_3416(v_3401);
  assign v_3418 = v_3419 | v_3438;
  assign v_3419 = act_3420 & 1'h1;
  assign act_3420 = v_3421 | v_3427;
  assign v_3421 = v_3422 & v_3428;
  assign v_3422 = v_3423 & vout_canPeek_3433;
  assign v_3423 = ~vout_canPeek_3424;
  pebbles_core
    pebbles_core_3424
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3425),
       .in0_consume_en(vin0_consume_en_3424),
       .out_canPeek(vout_canPeek_3424),
       .out_peek(vout_peek_3424));
  assign v_3425 = v_3426 | v_3431;
  assign v_3426 = mux_3426(v_3427);
  assign v_3427 = vout_canPeek_3424 & v_3428;
  assign v_3428 = v_3429 & 1'h1;
  assign v_3429 = v_3430 | 1'h0;
  assign v_3430 = ~v_3417;
  assign v_3431 = mux_3431(v_3432);
  assign v_3432 = ~v_3427;
  pebbles_core
    pebbles_core_3433
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3434),
       .in0_consume_en(vin0_consume_en_3433),
       .out_canPeek(vout_canPeek_3433),
       .out_peek(vout_peek_3433));
  assign v_3434 = v_3435 | v_3436;
  assign v_3435 = mux_3435(v_3421);
  assign v_3436 = mux_3436(v_3437);
  assign v_3437 = ~v_3421;
  assign v_3438 = v_3439 & 1'h1;
  assign v_3439 = v_3440 & v_3441;
  assign v_3440 = ~act_3420;
  assign v_3441 = v_3442 | v_3446;
  assign v_3442 = v_3443 | v_3444;
  assign v_3443 = mux_3443(v_3377);
  assign v_3444 = mux_3444(v_3445);
  assign v_3445 = ~v_3377;
  assign v_3446 = ~v_3417;
  assign v_3447 = v_3448 | v_3449;
  assign v_3448 = mux_3448(v_3419);
  assign v_3449 = mux_3449(v_3438);
  assign v_3450 = v_3451 & 1'h1;
  assign v_3451 = v_3452 & v_3453;
  assign v_3452 = ~act_3376;
  assign v_3453 = v_3454 | v_3458;
  assign v_3454 = v_3455 | v_3456;
  assign v_3455 = mux_3455(v_3277);
  assign v_3456 = mux_3456(v_3457);
  assign v_3457 = ~v_3277;
  assign v_3458 = ~v_3373;
  assign v_3459 = v_3460 | v_3461;
  assign v_3460 = mux_3460(v_3375);
  assign v_3461 = mux_3461(v_3450);
  assign v_3462 = v_3463 & 1'h1;
  assign v_3463 = v_3464 & v_3465;
  assign v_3464 = ~act_3276;
  assign v_3465 = v_3466 | v_3470;
  assign v_3466 = v_3467 | v_3468;
  assign v_3467 = mux_3467(v_3065);
  assign v_3468 = mux_3468(v_3469);
  assign v_3469 = ~v_3065;
  assign v_3470 = ~v_3273;
  assign v_3471 = v_3472 | v_3473;
  assign v_3472 = mux_3472(v_3275);
  assign v_3473 = mux_3473(v_3462);
  assign v_3474 = v_3475 & 1'h1;
  assign v_3475 = v_3476 & v_3477;
  assign v_3476 = ~act_3064;
  assign v_3477 = v_3478 | v_3482;
  assign v_3478 = v_3479 | v_3480;
  assign v_3479 = mux_3479(v_2629);
  assign v_3480 = mux_3480(v_3481);
  assign v_3481 = ~v_2629;
  assign v_3482 = ~v_3061;
  assign v_3483 = v_3484 | v_3485;
  assign v_3484 = mux_3484(v_3063);
  assign v_3485 = mux_3485(v_3474);
  assign v_3486 = v_3487 & 1'h1;
  assign v_3487 = v_3488 & v_3489;
  assign v_3488 = ~act_2628;
  assign v_3489 = v_3490 | v_3498;
  assign v_3490 = v_3491 | v_3496;
  assign v_3491 = mux_3491(v_3492);
  assign v_3492 = v_2625 & v_3493;
  assign v_3493 = v_3494 & 1'h1;
  assign v_3494 = v_3495 | 1'h0;
  assign v_3495 = ~v_2618;
  assign v_3496 = mux_3496(v_3497);
  assign v_3497 = ~v_3492;
  assign v_3498 = ~v_2625;
  assign v_3499 = v_3500 | v_3501;
  assign v_3500 = mux_3500(v_2627);
  assign v_3501 = mux_3501(v_3486);
  assign v_3503 = v_3504 | v_4363;
  assign v_3504 = act_3505 & 1'h1;
  assign act_3505 = v_3506 | v_3928;
  assign v_3506 = v_3507 & v_3929;
  assign v_3507 = v_3508 & v_3938;
  assign v_3508 = ~v_3509;
  assign v_3510 = v_3511 | v_3922;
  assign v_3511 = act_3512 & 1'h1;
  assign act_3512 = v_3513 | v_3711;
  assign v_3513 = v_3514 & v_3712;
  assign v_3514 = v_3515 & v_3721;
  assign v_3515 = ~v_3516;
  assign v_3517 = v_3518 | v_3705;
  assign v_3518 = act_3519 & 1'h1;
  assign act_3519 = v_3520 | v_3606;
  assign v_3520 = v_3521 & v_3607;
  assign v_3521 = v_3522 & v_3616;
  assign v_3522 = ~v_3523;
  assign v_3524 = v_3525 | v_3600;
  assign v_3525 = act_3526 & 1'h1;
  assign act_3526 = v_3527 | v_3557;
  assign v_3527 = v_3528 & v_3558;
  assign v_3528 = v_3529 & v_3567;
  assign v_3529 = ~v_3530;
  assign v_3531 = v_3532 | v_3551;
  assign v_3532 = act_3533 & 1'h1;
  assign act_3533 = v_3534 | v_3540;
  assign v_3534 = v_3535 & v_3541;
  assign v_3535 = v_3536 & vout_canPeek_3546;
  assign v_3536 = ~vout_canPeek_3537;
  pebbles_core
    pebbles_core_3537
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3538),
       .in0_consume_en(vin0_consume_en_3537),
       .out_canPeek(vout_canPeek_3537),
       .out_peek(vout_peek_3537));
  assign v_3538 = v_3539 | v_3544;
  assign v_3539 = mux_3539(v_3540);
  assign v_3540 = vout_canPeek_3537 & v_3541;
  assign v_3541 = v_3542 & 1'h1;
  assign v_3542 = v_3543 | 1'h0;
  assign v_3543 = ~v_3530;
  assign v_3544 = mux_3544(v_3545);
  assign v_3545 = ~v_3540;
  pebbles_core
    pebbles_core_3546
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3547),
       .in0_consume_en(vin0_consume_en_3546),
       .out_canPeek(vout_canPeek_3546),
       .out_peek(vout_peek_3546));
  assign v_3547 = v_3548 | v_3549;
  assign v_3548 = mux_3548(v_3534);
  assign v_3549 = mux_3549(v_3550);
  assign v_3550 = ~v_3534;
  assign v_3551 = v_3552 & 1'h1;
  assign v_3552 = v_3553 & v_3554;
  assign v_3553 = ~act_3533;
  assign v_3554 = v_3555 | v_3563;
  assign v_3555 = v_3556 | v_3561;
  assign v_3556 = mux_3556(v_3557);
  assign v_3557 = v_3530 & v_3558;
  assign v_3558 = v_3559 & 1'h1;
  assign v_3559 = v_3560 | 1'h0;
  assign v_3560 = ~v_3523;
  assign v_3561 = mux_3561(v_3562);
  assign v_3562 = ~v_3557;
  assign v_3563 = ~v_3530;
  assign v_3564 = v_3565 | v_3566;
  assign v_3565 = mux_3565(v_3532);
  assign v_3566 = mux_3566(v_3551);
  assign v_3568 = v_3569 | v_3588;
  assign v_3569 = act_3570 & 1'h1;
  assign act_3570 = v_3571 | v_3577;
  assign v_3571 = v_3572 & v_3578;
  assign v_3572 = v_3573 & vout_canPeek_3583;
  assign v_3573 = ~vout_canPeek_3574;
  pebbles_core
    pebbles_core_3574
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3575),
       .in0_consume_en(vin0_consume_en_3574),
       .out_canPeek(vout_canPeek_3574),
       .out_peek(vout_peek_3574));
  assign v_3575 = v_3576 | v_3581;
  assign v_3576 = mux_3576(v_3577);
  assign v_3577 = vout_canPeek_3574 & v_3578;
  assign v_3578 = v_3579 & 1'h1;
  assign v_3579 = v_3580 | 1'h0;
  assign v_3580 = ~v_3567;
  assign v_3581 = mux_3581(v_3582);
  assign v_3582 = ~v_3577;
  pebbles_core
    pebbles_core_3583
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3584),
       .in0_consume_en(vin0_consume_en_3583),
       .out_canPeek(vout_canPeek_3583),
       .out_peek(vout_peek_3583));
  assign v_3584 = v_3585 | v_3586;
  assign v_3585 = mux_3585(v_3571);
  assign v_3586 = mux_3586(v_3587);
  assign v_3587 = ~v_3571;
  assign v_3588 = v_3589 & 1'h1;
  assign v_3589 = v_3590 & v_3591;
  assign v_3590 = ~act_3570;
  assign v_3591 = v_3592 | v_3596;
  assign v_3592 = v_3593 | v_3594;
  assign v_3593 = mux_3593(v_3527);
  assign v_3594 = mux_3594(v_3595);
  assign v_3595 = ~v_3527;
  assign v_3596 = ~v_3567;
  assign v_3597 = v_3598 | v_3599;
  assign v_3598 = mux_3598(v_3569);
  assign v_3599 = mux_3599(v_3588);
  assign v_3600 = v_3601 & 1'h1;
  assign v_3601 = v_3602 & v_3603;
  assign v_3602 = ~act_3526;
  assign v_3603 = v_3604 | v_3612;
  assign v_3604 = v_3605 | v_3610;
  assign v_3605 = mux_3605(v_3606);
  assign v_3606 = v_3523 & v_3607;
  assign v_3607 = v_3608 & 1'h1;
  assign v_3608 = v_3609 | 1'h0;
  assign v_3609 = ~v_3516;
  assign v_3610 = mux_3610(v_3611);
  assign v_3611 = ~v_3606;
  assign v_3612 = ~v_3523;
  assign v_3613 = v_3614 | v_3615;
  assign v_3614 = mux_3614(v_3525);
  assign v_3615 = mux_3615(v_3600);
  assign v_3617 = v_3618 | v_3693;
  assign v_3618 = act_3619 & 1'h1;
  assign act_3619 = v_3620 | v_3650;
  assign v_3620 = v_3621 & v_3651;
  assign v_3621 = v_3622 & v_3660;
  assign v_3622 = ~v_3623;
  assign v_3624 = v_3625 | v_3644;
  assign v_3625 = act_3626 & 1'h1;
  assign act_3626 = v_3627 | v_3633;
  assign v_3627 = v_3628 & v_3634;
  assign v_3628 = v_3629 & vout_canPeek_3639;
  assign v_3629 = ~vout_canPeek_3630;
  pebbles_core
    pebbles_core_3630
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3631),
       .in0_consume_en(vin0_consume_en_3630),
       .out_canPeek(vout_canPeek_3630),
       .out_peek(vout_peek_3630));
  assign v_3631 = v_3632 | v_3637;
  assign v_3632 = mux_3632(v_3633);
  assign v_3633 = vout_canPeek_3630 & v_3634;
  assign v_3634 = v_3635 & 1'h1;
  assign v_3635 = v_3636 | 1'h0;
  assign v_3636 = ~v_3623;
  assign v_3637 = mux_3637(v_3638);
  assign v_3638 = ~v_3633;
  pebbles_core
    pebbles_core_3639
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3640),
       .in0_consume_en(vin0_consume_en_3639),
       .out_canPeek(vout_canPeek_3639),
       .out_peek(vout_peek_3639));
  assign v_3640 = v_3641 | v_3642;
  assign v_3641 = mux_3641(v_3627);
  assign v_3642 = mux_3642(v_3643);
  assign v_3643 = ~v_3627;
  assign v_3644 = v_3645 & 1'h1;
  assign v_3645 = v_3646 & v_3647;
  assign v_3646 = ~act_3626;
  assign v_3647 = v_3648 | v_3656;
  assign v_3648 = v_3649 | v_3654;
  assign v_3649 = mux_3649(v_3650);
  assign v_3650 = v_3623 & v_3651;
  assign v_3651 = v_3652 & 1'h1;
  assign v_3652 = v_3653 | 1'h0;
  assign v_3653 = ~v_3616;
  assign v_3654 = mux_3654(v_3655);
  assign v_3655 = ~v_3650;
  assign v_3656 = ~v_3623;
  assign v_3657 = v_3658 | v_3659;
  assign v_3658 = mux_3658(v_3625);
  assign v_3659 = mux_3659(v_3644);
  assign v_3661 = v_3662 | v_3681;
  assign v_3662 = act_3663 & 1'h1;
  assign act_3663 = v_3664 | v_3670;
  assign v_3664 = v_3665 & v_3671;
  assign v_3665 = v_3666 & vout_canPeek_3676;
  assign v_3666 = ~vout_canPeek_3667;
  pebbles_core
    pebbles_core_3667
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3668),
       .in0_consume_en(vin0_consume_en_3667),
       .out_canPeek(vout_canPeek_3667),
       .out_peek(vout_peek_3667));
  assign v_3668 = v_3669 | v_3674;
  assign v_3669 = mux_3669(v_3670);
  assign v_3670 = vout_canPeek_3667 & v_3671;
  assign v_3671 = v_3672 & 1'h1;
  assign v_3672 = v_3673 | 1'h0;
  assign v_3673 = ~v_3660;
  assign v_3674 = mux_3674(v_3675);
  assign v_3675 = ~v_3670;
  pebbles_core
    pebbles_core_3676
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3677),
       .in0_consume_en(vin0_consume_en_3676),
       .out_canPeek(vout_canPeek_3676),
       .out_peek(vout_peek_3676));
  assign v_3677 = v_3678 | v_3679;
  assign v_3678 = mux_3678(v_3664);
  assign v_3679 = mux_3679(v_3680);
  assign v_3680 = ~v_3664;
  assign v_3681 = v_3682 & 1'h1;
  assign v_3682 = v_3683 & v_3684;
  assign v_3683 = ~act_3663;
  assign v_3684 = v_3685 | v_3689;
  assign v_3685 = v_3686 | v_3687;
  assign v_3686 = mux_3686(v_3620);
  assign v_3687 = mux_3687(v_3688);
  assign v_3688 = ~v_3620;
  assign v_3689 = ~v_3660;
  assign v_3690 = v_3691 | v_3692;
  assign v_3691 = mux_3691(v_3662);
  assign v_3692 = mux_3692(v_3681);
  assign v_3693 = v_3694 & 1'h1;
  assign v_3694 = v_3695 & v_3696;
  assign v_3695 = ~act_3619;
  assign v_3696 = v_3697 | v_3701;
  assign v_3697 = v_3698 | v_3699;
  assign v_3698 = mux_3698(v_3520);
  assign v_3699 = mux_3699(v_3700);
  assign v_3700 = ~v_3520;
  assign v_3701 = ~v_3616;
  assign v_3702 = v_3703 | v_3704;
  assign v_3703 = mux_3703(v_3618);
  assign v_3704 = mux_3704(v_3693);
  assign v_3705 = v_3706 & 1'h1;
  assign v_3706 = v_3707 & v_3708;
  assign v_3707 = ~act_3519;
  assign v_3708 = v_3709 | v_3717;
  assign v_3709 = v_3710 | v_3715;
  assign v_3710 = mux_3710(v_3711);
  assign v_3711 = v_3516 & v_3712;
  assign v_3712 = v_3713 & 1'h1;
  assign v_3713 = v_3714 | 1'h0;
  assign v_3714 = ~v_3509;
  assign v_3715 = mux_3715(v_3716);
  assign v_3716 = ~v_3711;
  assign v_3717 = ~v_3516;
  assign v_3718 = v_3719 | v_3720;
  assign v_3719 = mux_3719(v_3518);
  assign v_3720 = mux_3720(v_3705);
  assign v_3722 = v_3723 | v_3910;
  assign v_3723 = act_3724 & 1'h1;
  assign act_3724 = v_3725 | v_3811;
  assign v_3725 = v_3726 & v_3812;
  assign v_3726 = v_3727 & v_3821;
  assign v_3727 = ~v_3728;
  assign v_3729 = v_3730 | v_3805;
  assign v_3730 = act_3731 & 1'h1;
  assign act_3731 = v_3732 | v_3762;
  assign v_3732 = v_3733 & v_3763;
  assign v_3733 = v_3734 & v_3772;
  assign v_3734 = ~v_3735;
  assign v_3736 = v_3737 | v_3756;
  assign v_3737 = act_3738 & 1'h1;
  assign act_3738 = v_3739 | v_3745;
  assign v_3739 = v_3740 & v_3746;
  assign v_3740 = v_3741 & vout_canPeek_3751;
  assign v_3741 = ~vout_canPeek_3742;
  pebbles_core
    pebbles_core_3742
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3743),
       .in0_consume_en(vin0_consume_en_3742),
       .out_canPeek(vout_canPeek_3742),
       .out_peek(vout_peek_3742));
  assign v_3743 = v_3744 | v_3749;
  assign v_3744 = mux_3744(v_3745);
  assign v_3745 = vout_canPeek_3742 & v_3746;
  assign v_3746 = v_3747 & 1'h1;
  assign v_3747 = v_3748 | 1'h0;
  assign v_3748 = ~v_3735;
  assign v_3749 = mux_3749(v_3750);
  assign v_3750 = ~v_3745;
  pebbles_core
    pebbles_core_3751
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3752),
       .in0_consume_en(vin0_consume_en_3751),
       .out_canPeek(vout_canPeek_3751),
       .out_peek(vout_peek_3751));
  assign v_3752 = v_3753 | v_3754;
  assign v_3753 = mux_3753(v_3739);
  assign v_3754 = mux_3754(v_3755);
  assign v_3755 = ~v_3739;
  assign v_3756 = v_3757 & 1'h1;
  assign v_3757 = v_3758 & v_3759;
  assign v_3758 = ~act_3738;
  assign v_3759 = v_3760 | v_3768;
  assign v_3760 = v_3761 | v_3766;
  assign v_3761 = mux_3761(v_3762);
  assign v_3762 = v_3735 & v_3763;
  assign v_3763 = v_3764 & 1'h1;
  assign v_3764 = v_3765 | 1'h0;
  assign v_3765 = ~v_3728;
  assign v_3766 = mux_3766(v_3767);
  assign v_3767 = ~v_3762;
  assign v_3768 = ~v_3735;
  assign v_3769 = v_3770 | v_3771;
  assign v_3770 = mux_3770(v_3737);
  assign v_3771 = mux_3771(v_3756);
  assign v_3773 = v_3774 | v_3793;
  assign v_3774 = act_3775 & 1'h1;
  assign act_3775 = v_3776 | v_3782;
  assign v_3776 = v_3777 & v_3783;
  assign v_3777 = v_3778 & vout_canPeek_3788;
  assign v_3778 = ~vout_canPeek_3779;
  pebbles_core
    pebbles_core_3779
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3780),
       .in0_consume_en(vin0_consume_en_3779),
       .out_canPeek(vout_canPeek_3779),
       .out_peek(vout_peek_3779));
  assign v_3780 = v_3781 | v_3786;
  assign v_3781 = mux_3781(v_3782);
  assign v_3782 = vout_canPeek_3779 & v_3783;
  assign v_3783 = v_3784 & 1'h1;
  assign v_3784 = v_3785 | 1'h0;
  assign v_3785 = ~v_3772;
  assign v_3786 = mux_3786(v_3787);
  assign v_3787 = ~v_3782;
  pebbles_core
    pebbles_core_3788
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3789),
       .in0_consume_en(vin0_consume_en_3788),
       .out_canPeek(vout_canPeek_3788),
       .out_peek(vout_peek_3788));
  assign v_3789 = v_3790 | v_3791;
  assign v_3790 = mux_3790(v_3776);
  assign v_3791 = mux_3791(v_3792);
  assign v_3792 = ~v_3776;
  assign v_3793 = v_3794 & 1'h1;
  assign v_3794 = v_3795 & v_3796;
  assign v_3795 = ~act_3775;
  assign v_3796 = v_3797 | v_3801;
  assign v_3797 = v_3798 | v_3799;
  assign v_3798 = mux_3798(v_3732);
  assign v_3799 = mux_3799(v_3800);
  assign v_3800 = ~v_3732;
  assign v_3801 = ~v_3772;
  assign v_3802 = v_3803 | v_3804;
  assign v_3803 = mux_3803(v_3774);
  assign v_3804 = mux_3804(v_3793);
  assign v_3805 = v_3806 & 1'h1;
  assign v_3806 = v_3807 & v_3808;
  assign v_3807 = ~act_3731;
  assign v_3808 = v_3809 | v_3817;
  assign v_3809 = v_3810 | v_3815;
  assign v_3810 = mux_3810(v_3811);
  assign v_3811 = v_3728 & v_3812;
  assign v_3812 = v_3813 & 1'h1;
  assign v_3813 = v_3814 | 1'h0;
  assign v_3814 = ~v_3721;
  assign v_3815 = mux_3815(v_3816);
  assign v_3816 = ~v_3811;
  assign v_3817 = ~v_3728;
  assign v_3818 = v_3819 | v_3820;
  assign v_3819 = mux_3819(v_3730);
  assign v_3820 = mux_3820(v_3805);
  assign v_3822 = v_3823 | v_3898;
  assign v_3823 = act_3824 & 1'h1;
  assign act_3824 = v_3825 | v_3855;
  assign v_3825 = v_3826 & v_3856;
  assign v_3826 = v_3827 & v_3865;
  assign v_3827 = ~v_3828;
  assign v_3829 = v_3830 | v_3849;
  assign v_3830 = act_3831 & 1'h1;
  assign act_3831 = v_3832 | v_3838;
  assign v_3832 = v_3833 & v_3839;
  assign v_3833 = v_3834 & vout_canPeek_3844;
  assign v_3834 = ~vout_canPeek_3835;
  pebbles_core
    pebbles_core_3835
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3836),
       .in0_consume_en(vin0_consume_en_3835),
       .out_canPeek(vout_canPeek_3835),
       .out_peek(vout_peek_3835));
  assign v_3836 = v_3837 | v_3842;
  assign v_3837 = mux_3837(v_3838);
  assign v_3838 = vout_canPeek_3835 & v_3839;
  assign v_3839 = v_3840 & 1'h1;
  assign v_3840 = v_3841 | 1'h0;
  assign v_3841 = ~v_3828;
  assign v_3842 = mux_3842(v_3843);
  assign v_3843 = ~v_3838;
  pebbles_core
    pebbles_core_3844
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3845),
       .in0_consume_en(vin0_consume_en_3844),
       .out_canPeek(vout_canPeek_3844),
       .out_peek(vout_peek_3844));
  assign v_3845 = v_3846 | v_3847;
  assign v_3846 = mux_3846(v_3832);
  assign v_3847 = mux_3847(v_3848);
  assign v_3848 = ~v_3832;
  assign v_3849 = v_3850 & 1'h1;
  assign v_3850 = v_3851 & v_3852;
  assign v_3851 = ~act_3831;
  assign v_3852 = v_3853 | v_3861;
  assign v_3853 = v_3854 | v_3859;
  assign v_3854 = mux_3854(v_3855);
  assign v_3855 = v_3828 & v_3856;
  assign v_3856 = v_3857 & 1'h1;
  assign v_3857 = v_3858 | 1'h0;
  assign v_3858 = ~v_3821;
  assign v_3859 = mux_3859(v_3860);
  assign v_3860 = ~v_3855;
  assign v_3861 = ~v_3828;
  assign v_3862 = v_3863 | v_3864;
  assign v_3863 = mux_3863(v_3830);
  assign v_3864 = mux_3864(v_3849);
  assign v_3866 = v_3867 | v_3886;
  assign v_3867 = act_3868 & 1'h1;
  assign act_3868 = v_3869 | v_3875;
  assign v_3869 = v_3870 & v_3876;
  assign v_3870 = v_3871 & vout_canPeek_3881;
  assign v_3871 = ~vout_canPeek_3872;
  pebbles_core
    pebbles_core_3872
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3873),
       .in0_consume_en(vin0_consume_en_3872),
       .out_canPeek(vout_canPeek_3872),
       .out_peek(vout_peek_3872));
  assign v_3873 = v_3874 | v_3879;
  assign v_3874 = mux_3874(v_3875);
  assign v_3875 = vout_canPeek_3872 & v_3876;
  assign v_3876 = v_3877 & 1'h1;
  assign v_3877 = v_3878 | 1'h0;
  assign v_3878 = ~v_3865;
  assign v_3879 = mux_3879(v_3880);
  assign v_3880 = ~v_3875;
  pebbles_core
    pebbles_core_3881
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3882),
       .in0_consume_en(vin0_consume_en_3881),
       .out_canPeek(vout_canPeek_3881),
       .out_peek(vout_peek_3881));
  assign v_3882 = v_3883 | v_3884;
  assign v_3883 = mux_3883(v_3869);
  assign v_3884 = mux_3884(v_3885);
  assign v_3885 = ~v_3869;
  assign v_3886 = v_3887 & 1'h1;
  assign v_3887 = v_3888 & v_3889;
  assign v_3888 = ~act_3868;
  assign v_3889 = v_3890 | v_3894;
  assign v_3890 = v_3891 | v_3892;
  assign v_3891 = mux_3891(v_3825);
  assign v_3892 = mux_3892(v_3893);
  assign v_3893 = ~v_3825;
  assign v_3894 = ~v_3865;
  assign v_3895 = v_3896 | v_3897;
  assign v_3896 = mux_3896(v_3867);
  assign v_3897 = mux_3897(v_3886);
  assign v_3898 = v_3899 & 1'h1;
  assign v_3899 = v_3900 & v_3901;
  assign v_3900 = ~act_3824;
  assign v_3901 = v_3902 | v_3906;
  assign v_3902 = v_3903 | v_3904;
  assign v_3903 = mux_3903(v_3725);
  assign v_3904 = mux_3904(v_3905);
  assign v_3905 = ~v_3725;
  assign v_3906 = ~v_3821;
  assign v_3907 = v_3908 | v_3909;
  assign v_3908 = mux_3908(v_3823);
  assign v_3909 = mux_3909(v_3898);
  assign v_3910 = v_3911 & 1'h1;
  assign v_3911 = v_3912 & v_3913;
  assign v_3912 = ~act_3724;
  assign v_3913 = v_3914 | v_3918;
  assign v_3914 = v_3915 | v_3916;
  assign v_3915 = mux_3915(v_3513);
  assign v_3916 = mux_3916(v_3917);
  assign v_3917 = ~v_3513;
  assign v_3918 = ~v_3721;
  assign v_3919 = v_3920 | v_3921;
  assign v_3920 = mux_3920(v_3723);
  assign v_3921 = mux_3921(v_3910);
  assign v_3922 = v_3923 & 1'h1;
  assign v_3923 = v_3924 & v_3925;
  assign v_3924 = ~act_3512;
  assign v_3925 = v_3926 | v_3934;
  assign v_3926 = v_3927 | v_3932;
  assign v_3927 = mux_3927(v_3928);
  assign v_3928 = v_3509 & v_3929;
  assign v_3929 = v_3930 & 1'h1;
  assign v_3930 = v_3931 | 1'h0;
  assign v_3931 = ~v_3502;
  assign v_3932 = mux_3932(v_3933);
  assign v_3933 = ~v_3928;
  assign v_3934 = ~v_3509;
  assign v_3935 = v_3936 | v_3937;
  assign v_3936 = mux_3936(v_3511);
  assign v_3937 = mux_3937(v_3922);
  assign v_3939 = v_3940 | v_4351;
  assign v_3940 = act_3941 & 1'h1;
  assign act_3941 = v_3942 | v_4140;
  assign v_3942 = v_3943 & v_4141;
  assign v_3943 = v_3944 & v_4150;
  assign v_3944 = ~v_3945;
  assign v_3946 = v_3947 | v_4134;
  assign v_3947 = act_3948 & 1'h1;
  assign act_3948 = v_3949 | v_4035;
  assign v_3949 = v_3950 & v_4036;
  assign v_3950 = v_3951 & v_4045;
  assign v_3951 = ~v_3952;
  assign v_3953 = v_3954 | v_4029;
  assign v_3954 = act_3955 & 1'h1;
  assign act_3955 = v_3956 | v_3986;
  assign v_3956 = v_3957 & v_3987;
  assign v_3957 = v_3958 & v_3996;
  assign v_3958 = ~v_3959;
  assign v_3960 = v_3961 | v_3980;
  assign v_3961 = act_3962 & 1'h1;
  assign act_3962 = v_3963 | v_3969;
  assign v_3963 = v_3964 & v_3970;
  assign v_3964 = v_3965 & vout_canPeek_3975;
  assign v_3965 = ~vout_canPeek_3966;
  pebbles_core
    pebbles_core_3966
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3967),
       .in0_consume_en(vin0_consume_en_3966),
       .out_canPeek(vout_canPeek_3966),
       .out_peek(vout_peek_3966));
  assign v_3967 = v_3968 | v_3973;
  assign v_3968 = mux_3968(v_3969);
  assign v_3969 = vout_canPeek_3966 & v_3970;
  assign v_3970 = v_3971 & 1'h1;
  assign v_3971 = v_3972 | 1'h0;
  assign v_3972 = ~v_3959;
  assign v_3973 = mux_3973(v_3974);
  assign v_3974 = ~v_3969;
  pebbles_core
    pebbles_core_3975
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_3976),
       .in0_consume_en(vin0_consume_en_3975),
       .out_canPeek(vout_canPeek_3975),
       .out_peek(vout_peek_3975));
  assign v_3976 = v_3977 | v_3978;
  assign v_3977 = mux_3977(v_3963);
  assign v_3978 = mux_3978(v_3979);
  assign v_3979 = ~v_3963;
  assign v_3980 = v_3981 & 1'h1;
  assign v_3981 = v_3982 & v_3983;
  assign v_3982 = ~act_3962;
  assign v_3983 = v_3984 | v_3992;
  assign v_3984 = v_3985 | v_3990;
  assign v_3985 = mux_3985(v_3986);
  assign v_3986 = v_3959 & v_3987;
  assign v_3987 = v_3988 & 1'h1;
  assign v_3988 = v_3989 | 1'h0;
  assign v_3989 = ~v_3952;
  assign v_3990 = mux_3990(v_3991);
  assign v_3991 = ~v_3986;
  assign v_3992 = ~v_3959;
  assign v_3993 = v_3994 | v_3995;
  assign v_3994 = mux_3994(v_3961);
  assign v_3995 = mux_3995(v_3980);
  assign v_3997 = v_3998 | v_4017;
  assign v_3998 = act_3999 & 1'h1;
  assign act_3999 = v_4000 | v_4006;
  assign v_4000 = v_4001 & v_4007;
  assign v_4001 = v_4002 & vout_canPeek_4012;
  assign v_4002 = ~vout_canPeek_4003;
  pebbles_core
    pebbles_core_4003
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4004),
       .in0_consume_en(vin0_consume_en_4003),
       .out_canPeek(vout_canPeek_4003),
       .out_peek(vout_peek_4003));
  assign v_4004 = v_4005 | v_4010;
  assign v_4005 = mux_4005(v_4006);
  assign v_4006 = vout_canPeek_4003 & v_4007;
  assign v_4007 = v_4008 & 1'h1;
  assign v_4008 = v_4009 | 1'h0;
  assign v_4009 = ~v_3996;
  assign v_4010 = mux_4010(v_4011);
  assign v_4011 = ~v_4006;
  pebbles_core
    pebbles_core_4012
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4013),
       .in0_consume_en(vin0_consume_en_4012),
       .out_canPeek(vout_canPeek_4012),
       .out_peek(vout_peek_4012));
  assign v_4013 = v_4014 | v_4015;
  assign v_4014 = mux_4014(v_4000);
  assign v_4015 = mux_4015(v_4016);
  assign v_4016 = ~v_4000;
  assign v_4017 = v_4018 & 1'h1;
  assign v_4018 = v_4019 & v_4020;
  assign v_4019 = ~act_3999;
  assign v_4020 = v_4021 | v_4025;
  assign v_4021 = v_4022 | v_4023;
  assign v_4022 = mux_4022(v_3956);
  assign v_4023 = mux_4023(v_4024);
  assign v_4024 = ~v_3956;
  assign v_4025 = ~v_3996;
  assign v_4026 = v_4027 | v_4028;
  assign v_4027 = mux_4027(v_3998);
  assign v_4028 = mux_4028(v_4017);
  assign v_4029 = v_4030 & 1'h1;
  assign v_4030 = v_4031 & v_4032;
  assign v_4031 = ~act_3955;
  assign v_4032 = v_4033 | v_4041;
  assign v_4033 = v_4034 | v_4039;
  assign v_4034 = mux_4034(v_4035);
  assign v_4035 = v_3952 & v_4036;
  assign v_4036 = v_4037 & 1'h1;
  assign v_4037 = v_4038 | 1'h0;
  assign v_4038 = ~v_3945;
  assign v_4039 = mux_4039(v_4040);
  assign v_4040 = ~v_4035;
  assign v_4041 = ~v_3952;
  assign v_4042 = v_4043 | v_4044;
  assign v_4043 = mux_4043(v_3954);
  assign v_4044 = mux_4044(v_4029);
  assign v_4046 = v_4047 | v_4122;
  assign v_4047 = act_4048 & 1'h1;
  assign act_4048 = v_4049 | v_4079;
  assign v_4049 = v_4050 & v_4080;
  assign v_4050 = v_4051 & v_4089;
  assign v_4051 = ~v_4052;
  assign v_4053 = v_4054 | v_4073;
  assign v_4054 = act_4055 & 1'h1;
  assign act_4055 = v_4056 | v_4062;
  assign v_4056 = v_4057 & v_4063;
  assign v_4057 = v_4058 & vout_canPeek_4068;
  assign v_4058 = ~vout_canPeek_4059;
  pebbles_core
    pebbles_core_4059
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4060),
       .in0_consume_en(vin0_consume_en_4059),
       .out_canPeek(vout_canPeek_4059),
       .out_peek(vout_peek_4059));
  assign v_4060 = v_4061 | v_4066;
  assign v_4061 = mux_4061(v_4062);
  assign v_4062 = vout_canPeek_4059 & v_4063;
  assign v_4063 = v_4064 & 1'h1;
  assign v_4064 = v_4065 | 1'h0;
  assign v_4065 = ~v_4052;
  assign v_4066 = mux_4066(v_4067);
  assign v_4067 = ~v_4062;
  pebbles_core
    pebbles_core_4068
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4069),
       .in0_consume_en(vin0_consume_en_4068),
       .out_canPeek(vout_canPeek_4068),
       .out_peek(vout_peek_4068));
  assign v_4069 = v_4070 | v_4071;
  assign v_4070 = mux_4070(v_4056);
  assign v_4071 = mux_4071(v_4072);
  assign v_4072 = ~v_4056;
  assign v_4073 = v_4074 & 1'h1;
  assign v_4074 = v_4075 & v_4076;
  assign v_4075 = ~act_4055;
  assign v_4076 = v_4077 | v_4085;
  assign v_4077 = v_4078 | v_4083;
  assign v_4078 = mux_4078(v_4079);
  assign v_4079 = v_4052 & v_4080;
  assign v_4080 = v_4081 & 1'h1;
  assign v_4081 = v_4082 | 1'h0;
  assign v_4082 = ~v_4045;
  assign v_4083 = mux_4083(v_4084);
  assign v_4084 = ~v_4079;
  assign v_4085 = ~v_4052;
  assign v_4086 = v_4087 | v_4088;
  assign v_4087 = mux_4087(v_4054);
  assign v_4088 = mux_4088(v_4073);
  assign v_4090 = v_4091 | v_4110;
  assign v_4091 = act_4092 & 1'h1;
  assign act_4092 = v_4093 | v_4099;
  assign v_4093 = v_4094 & v_4100;
  assign v_4094 = v_4095 & vout_canPeek_4105;
  assign v_4095 = ~vout_canPeek_4096;
  pebbles_core
    pebbles_core_4096
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4097),
       .in0_consume_en(vin0_consume_en_4096),
       .out_canPeek(vout_canPeek_4096),
       .out_peek(vout_peek_4096));
  assign v_4097 = v_4098 | v_4103;
  assign v_4098 = mux_4098(v_4099);
  assign v_4099 = vout_canPeek_4096 & v_4100;
  assign v_4100 = v_4101 & 1'h1;
  assign v_4101 = v_4102 | 1'h0;
  assign v_4102 = ~v_4089;
  assign v_4103 = mux_4103(v_4104);
  assign v_4104 = ~v_4099;
  pebbles_core
    pebbles_core_4105
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4106),
       .in0_consume_en(vin0_consume_en_4105),
       .out_canPeek(vout_canPeek_4105),
       .out_peek(vout_peek_4105));
  assign v_4106 = v_4107 | v_4108;
  assign v_4107 = mux_4107(v_4093);
  assign v_4108 = mux_4108(v_4109);
  assign v_4109 = ~v_4093;
  assign v_4110 = v_4111 & 1'h1;
  assign v_4111 = v_4112 & v_4113;
  assign v_4112 = ~act_4092;
  assign v_4113 = v_4114 | v_4118;
  assign v_4114 = v_4115 | v_4116;
  assign v_4115 = mux_4115(v_4049);
  assign v_4116 = mux_4116(v_4117);
  assign v_4117 = ~v_4049;
  assign v_4118 = ~v_4089;
  assign v_4119 = v_4120 | v_4121;
  assign v_4120 = mux_4120(v_4091);
  assign v_4121 = mux_4121(v_4110);
  assign v_4122 = v_4123 & 1'h1;
  assign v_4123 = v_4124 & v_4125;
  assign v_4124 = ~act_4048;
  assign v_4125 = v_4126 | v_4130;
  assign v_4126 = v_4127 | v_4128;
  assign v_4127 = mux_4127(v_3949);
  assign v_4128 = mux_4128(v_4129);
  assign v_4129 = ~v_3949;
  assign v_4130 = ~v_4045;
  assign v_4131 = v_4132 | v_4133;
  assign v_4132 = mux_4132(v_4047);
  assign v_4133 = mux_4133(v_4122);
  assign v_4134 = v_4135 & 1'h1;
  assign v_4135 = v_4136 & v_4137;
  assign v_4136 = ~act_3948;
  assign v_4137 = v_4138 | v_4146;
  assign v_4138 = v_4139 | v_4144;
  assign v_4139 = mux_4139(v_4140);
  assign v_4140 = v_3945 & v_4141;
  assign v_4141 = v_4142 & 1'h1;
  assign v_4142 = v_4143 | 1'h0;
  assign v_4143 = ~v_3938;
  assign v_4144 = mux_4144(v_4145);
  assign v_4145 = ~v_4140;
  assign v_4146 = ~v_3945;
  assign v_4147 = v_4148 | v_4149;
  assign v_4148 = mux_4148(v_3947);
  assign v_4149 = mux_4149(v_4134);
  assign v_4151 = v_4152 | v_4339;
  assign v_4152 = act_4153 & 1'h1;
  assign act_4153 = v_4154 | v_4240;
  assign v_4154 = v_4155 & v_4241;
  assign v_4155 = v_4156 & v_4250;
  assign v_4156 = ~v_4157;
  assign v_4158 = v_4159 | v_4234;
  assign v_4159 = act_4160 & 1'h1;
  assign act_4160 = v_4161 | v_4191;
  assign v_4161 = v_4162 & v_4192;
  assign v_4162 = v_4163 & v_4201;
  assign v_4163 = ~v_4164;
  assign v_4165 = v_4166 | v_4185;
  assign v_4166 = act_4167 & 1'h1;
  assign act_4167 = v_4168 | v_4174;
  assign v_4168 = v_4169 & v_4175;
  assign v_4169 = v_4170 & vout_canPeek_4180;
  assign v_4170 = ~vout_canPeek_4171;
  pebbles_core
    pebbles_core_4171
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4172),
       .in0_consume_en(vin0_consume_en_4171),
       .out_canPeek(vout_canPeek_4171),
       .out_peek(vout_peek_4171));
  assign v_4172 = v_4173 | v_4178;
  assign v_4173 = mux_4173(v_4174);
  assign v_4174 = vout_canPeek_4171 & v_4175;
  assign v_4175 = v_4176 & 1'h1;
  assign v_4176 = v_4177 | 1'h0;
  assign v_4177 = ~v_4164;
  assign v_4178 = mux_4178(v_4179);
  assign v_4179 = ~v_4174;
  pebbles_core
    pebbles_core_4180
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4181),
       .in0_consume_en(vin0_consume_en_4180),
       .out_canPeek(vout_canPeek_4180),
       .out_peek(vout_peek_4180));
  assign v_4181 = v_4182 | v_4183;
  assign v_4182 = mux_4182(v_4168);
  assign v_4183 = mux_4183(v_4184);
  assign v_4184 = ~v_4168;
  assign v_4185 = v_4186 & 1'h1;
  assign v_4186 = v_4187 & v_4188;
  assign v_4187 = ~act_4167;
  assign v_4188 = v_4189 | v_4197;
  assign v_4189 = v_4190 | v_4195;
  assign v_4190 = mux_4190(v_4191);
  assign v_4191 = v_4164 & v_4192;
  assign v_4192 = v_4193 & 1'h1;
  assign v_4193 = v_4194 | 1'h0;
  assign v_4194 = ~v_4157;
  assign v_4195 = mux_4195(v_4196);
  assign v_4196 = ~v_4191;
  assign v_4197 = ~v_4164;
  assign v_4198 = v_4199 | v_4200;
  assign v_4199 = mux_4199(v_4166);
  assign v_4200 = mux_4200(v_4185);
  assign v_4202 = v_4203 | v_4222;
  assign v_4203 = act_4204 & 1'h1;
  assign act_4204 = v_4205 | v_4211;
  assign v_4205 = v_4206 & v_4212;
  assign v_4206 = v_4207 & vout_canPeek_4217;
  assign v_4207 = ~vout_canPeek_4208;
  pebbles_core
    pebbles_core_4208
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4209),
       .in0_consume_en(vin0_consume_en_4208),
       .out_canPeek(vout_canPeek_4208),
       .out_peek(vout_peek_4208));
  assign v_4209 = v_4210 | v_4215;
  assign v_4210 = mux_4210(v_4211);
  assign v_4211 = vout_canPeek_4208 & v_4212;
  assign v_4212 = v_4213 & 1'h1;
  assign v_4213 = v_4214 | 1'h0;
  assign v_4214 = ~v_4201;
  assign v_4215 = mux_4215(v_4216);
  assign v_4216 = ~v_4211;
  pebbles_core
    pebbles_core_4217
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4218),
       .in0_consume_en(vin0_consume_en_4217),
       .out_canPeek(vout_canPeek_4217),
       .out_peek(vout_peek_4217));
  assign v_4218 = v_4219 | v_4220;
  assign v_4219 = mux_4219(v_4205);
  assign v_4220 = mux_4220(v_4221);
  assign v_4221 = ~v_4205;
  assign v_4222 = v_4223 & 1'h1;
  assign v_4223 = v_4224 & v_4225;
  assign v_4224 = ~act_4204;
  assign v_4225 = v_4226 | v_4230;
  assign v_4226 = v_4227 | v_4228;
  assign v_4227 = mux_4227(v_4161);
  assign v_4228 = mux_4228(v_4229);
  assign v_4229 = ~v_4161;
  assign v_4230 = ~v_4201;
  assign v_4231 = v_4232 | v_4233;
  assign v_4232 = mux_4232(v_4203);
  assign v_4233 = mux_4233(v_4222);
  assign v_4234 = v_4235 & 1'h1;
  assign v_4235 = v_4236 & v_4237;
  assign v_4236 = ~act_4160;
  assign v_4237 = v_4238 | v_4246;
  assign v_4238 = v_4239 | v_4244;
  assign v_4239 = mux_4239(v_4240);
  assign v_4240 = v_4157 & v_4241;
  assign v_4241 = v_4242 & 1'h1;
  assign v_4242 = v_4243 | 1'h0;
  assign v_4243 = ~v_4150;
  assign v_4244 = mux_4244(v_4245);
  assign v_4245 = ~v_4240;
  assign v_4246 = ~v_4157;
  assign v_4247 = v_4248 | v_4249;
  assign v_4248 = mux_4248(v_4159);
  assign v_4249 = mux_4249(v_4234);
  assign v_4251 = v_4252 | v_4327;
  assign v_4252 = act_4253 & 1'h1;
  assign act_4253 = v_4254 | v_4284;
  assign v_4254 = v_4255 & v_4285;
  assign v_4255 = v_4256 & v_4294;
  assign v_4256 = ~v_4257;
  assign v_4258 = v_4259 | v_4278;
  assign v_4259 = act_4260 & 1'h1;
  assign act_4260 = v_4261 | v_4267;
  assign v_4261 = v_4262 & v_4268;
  assign v_4262 = v_4263 & vout_canPeek_4273;
  assign v_4263 = ~vout_canPeek_4264;
  pebbles_core
    pebbles_core_4264
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4265),
       .in0_consume_en(vin0_consume_en_4264),
       .out_canPeek(vout_canPeek_4264),
       .out_peek(vout_peek_4264));
  assign v_4265 = v_4266 | v_4271;
  assign v_4266 = mux_4266(v_4267);
  assign v_4267 = vout_canPeek_4264 & v_4268;
  assign v_4268 = v_4269 & 1'h1;
  assign v_4269 = v_4270 | 1'h0;
  assign v_4270 = ~v_4257;
  assign v_4271 = mux_4271(v_4272);
  assign v_4272 = ~v_4267;
  pebbles_core
    pebbles_core_4273
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4274),
       .in0_consume_en(vin0_consume_en_4273),
       .out_canPeek(vout_canPeek_4273),
       .out_peek(vout_peek_4273));
  assign v_4274 = v_4275 | v_4276;
  assign v_4275 = mux_4275(v_4261);
  assign v_4276 = mux_4276(v_4277);
  assign v_4277 = ~v_4261;
  assign v_4278 = v_4279 & 1'h1;
  assign v_4279 = v_4280 & v_4281;
  assign v_4280 = ~act_4260;
  assign v_4281 = v_4282 | v_4290;
  assign v_4282 = v_4283 | v_4288;
  assign v_4283 = mux_4283(v_4284);
  assign v_4284 = v_4257 & v_4285;
  assign v_4285 = v_4286 & 1'h1;
  assign v_4286 = v_4287 | 1'h0;
  assign v_4287 = ~v_4250;
  assign v_4288 = mux_4288(v_4289);
  assign v_4289 = ~v_4284;
  assign v_4290 = ~v_4257;
  assign v_4291 = v_4292 | v_4293;
  assign v_4292 = mux_4292(v_4259);
  assign v_4293 = mux_4293(v_4278);
  assign v_4295 = v_4296 | v_4315;
  assign v_4296 = act_4297 & 1'h1;
  assign act_4297 = v_4298 | v_4304;
  assign v_4298 = v_4299 & v_4305;
  assign v_4299 = v_4300 & vout_canPeek_4310;
  assign v_4300 = ~vout_canPeek_4301;
  pebbles_core
    pebbles_core_4301
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4302),
       .in0_consume_en(vin0_consume_en_4301),
       .out_canPeek(vout_canPeek_4301),
       .out_peek(vout_peek_4301));
  assign v_4302 = v_4303 | v_4308;
  assign v_4303 = mux_4303(v_4304);
  assign v_4304 = vout_canPeek_4301 & v_4305;
  assign v_4305 = v_4306 & 1'h1;
  assign v_4306 = v_4307 | 1'h0;
  assign v_4307 = ~v_4294;
  assign v_4308 = mux_4308(v_4309);
  assign v_4309 = ~v_4304;
  pebbles_core
    pebbles_core_4310
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4311),
       .in0_consume_en(vin0_consume_en_4310),
       .out_canPeek(vout_canPeek_4310),
       .out_peek(vout_peek_4310));
  assign v_4311 = v_4312 | v_4313;
  assign v_4312 = mux_4312(v_4298);
  assign v_4313 = mux_4313(v_4314);
  assign v_4314 = ~v_4298;
  assign v_4315 = v_4316 & 1'h1;
  assign v_4316 = v_4317 & v_4318;
  assign v_4317 = ~act_4297;
  assign v_4318 = v_4319 | v_4323;
  assign v_4319 = v_4320 | v_4321;
  assign v_4320 = mux_4320(v_4254);
  assign v_4321 = mux_4321(v_4322);
  assign v_4322 = ~v_4254;
  assign v_4323 = ~v_4294;
  assign v_4324 = v_4325 | v_4326;
  assign v_4325 = mux_4325(v_4296);
  assign v_4326 = mux_4326(v_4315);
  assign v_4327 = v_4328 & 1'h1;
  assign v_4328 = v_4329 & v_4330;
  assign v_4329 = ~act_4253;
  assign v_4330 = v_4331 | v_4335;
  assign v_4331 = v_4332 | v_4333;
  assign v_4332 = mux_4332(v_4154);
  assign v_4333 = mux_4333(v_4334);
  assign v_4334 = ~v_4154;
  assign v_4335 = ~v_4250;
  assign v_4336 = v_4337 | v_4338;
  assign v_4337 = mux_4337(v_4252);
  assign v_4338 = mux_4338(v_4327);
  assign v_4339 = v_4340 & 1'h1;
  assign v_4340 = v_4341 & v_4342;
  assign v_4341 = ~act_4153;
  assign v_4342 = v_4343 | v_4347;
  assign v_4343 = v_4344 | v_4345;
  assign v_4344 = mux_4344(v_3942);
  assign v_4345 = mux_4345(v_4346);
  assign v_4346 = ~v_3942;
  assign v_4347 = ~v_4150;
  assign v_4348 = v_4349 | v_4350;
  assign v_4349 = mux_4349(v_4152);
  assign v_4350 = mux_4350(v_4339);
  assign v_4351 = v_4352 & 1'h1;
  assign v_4352 = v_4353 & v_4354;
  assign v_4353 = ~act_3941;
  assign v_4354 = v_4355 | v_4359;
  assign v_4355 = v_4356 | v_4357;
  assign v_4356 = mux_4356(v_3506);
  assign v_4357 = mux_4357(v_4358);
  assign v_4358 = ~v_3506;
  assign v_4359 = ~v_3938;
  assign v_4360 = v_4361 | v_4362;
  assign v_4361 = mux_4361(v_3940);
  assign v_4362 = mux_4362(v_4351);
  assign v_4363 = v_4364 & 1'h1;
  assign v_4364 = v_4365 & v_4366;
  assign v_4365 = ~act_3505;
  assign v_4366 = v_4367 | v_4371;
  assign v_4367 = v_4368 | v_4369;
  assign v_4368 = mux_4368(v_2622);
  assign v_4369 = mux_4369(v_4370);
  assign v_4370 = ~v_2622;
  assign v_4371 = ~v_3502;
  assign v_4372 = v_4373 | v_4374;
  assign v_4373 = mux_4373(v_3504);
  assign v_4374 = mux_4374(v_4363);
  assign v_4375 = v_4376 & 1'h1;
  assign v_4376 = v_4377 & v_4378;
  assign v_4377 = ~act_2621;
  assign v_4378 = v_4379 | v_22325;
  assign v_4379 = v_4380 | v_22323;
  assign v_4380 = mux_4380(v_4381);
  assign v_4381 = v_2618 & v_4382;
  assign v_4382 = v_4383 & 1'h1;
  assign v_4383 = v_4384 | 1'h0;
  assign v_4384 = ~v_4385;
  assign v_4386 = v_4387 | v_4389;
  assign v_4387 = act_4388 & 1'h1;
  assign act_4388 = v_2615 | v_4381;
  assign v_4389 = v_4390 & 1'h1;
  assign v_4390 = v_4391 & v_4392;
  assign v_4391 = ~act_4388;
  assign v_4392 = v_4393 | v_22319;
  assign v_4393 = v_4394 | v_22317;
  assign v_4394 = mux_4394(v_4395);
  assign v_4395 = v_4396 & v_7954;
  assign v_4396 = v_4397 & v_4385;
  assign v_4397 = ~v_4398;
  assign v_4399 = v_4400 | v_7947;
  assign v_4400 = act_4401 & 1'h1;
  assign act_4401 = v_4402 | v_6168;
  assign v_4402 = v_4403 & v_6169;
  assign v_4403 = v_4404 & v_6178;
  assign v_4404 = ~v_4405;
  assign v_4406 = v_4407 | v_6162;
  assign v_4407 = act_4408 & 1'h1;
  assign act_4408 = v_4409 | v_5279;
  assign v_4409 = v_4410 & v_5280;
  assign v_4410 = v_4411 & v_5289;
  assign v_4411 = ~v_4412;
  assign v_4413 = v_4414 | v_5273;
  assign v_4414 = act_4415 & 1'h1;
  assign act_4415 = v_4416 | v_4838;
  assign v_4416 = v_4417 & v_4839;
  assign v_4417 = v_4418 & v_4848;
  assign v_4418 = ~v_4419;
  assign v_4420 = v_4421 | v_4832;
  assign v_4421 = act_4422 & 1'h1;
  assign act_4422 = v_4423 | v_4621;
  assign v_4423 = v_4424 & v_4622;
  assign v_4424 = v_4425 & v_4631;
  assign v_4425 = ~v_4426;
  assign v_4427 = v_4428 | v_4615;
  assign v_4428 = act_4429 & 1'h1;
  assign act_4429 = v_4430 | v_4516;
  assign v_4430 = v_4431 & v_4517;
  assign v_4431 = v_4432 & v_4526;
  assign v_4432 = ~v_4433;
  assign v_4434 = v_4435 | v_4510;
  assign v_4435 = act_4436 & 1'h1;
  assign act_4436 = v_4437 | v_4467;
  assign v_4437 = v_4438 & v_4468;
  assign v_4438 = v_4439 & v_4477;
  assign v_4439 = ~v_4440;
  assign v_4441 = v_4442 | v_4461;
  assign v_4442 = act_4443 & 1'h1;
  assign act_4443 = v_4444 | v_4450;
  assign v_4444 = v_4445 & v_4451;
  assign v_4445 = v_4446 & vout_canPeek_4456;
  assign v_4446 = ~vout_canPeek_4447;
  pebbles_core
    pebbles_core_4447
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4448),
       .in0_consume_en(vin0_consume_en_4447),
       .out_canPeek(vout_canPeek_4447),
       .out_peek(vout_peek_4447));
  assign v_4448 = v_4449 | v_4454;
  assign v_4449 = mux_4449(v_4450);
  assign v_4450 = vout_canPeek_4447 & v_4451;
  assign v_4451 = v_4452 & 1'h1;
  assign v_4452 = v_4453 | 1'h0;
  assign v_4453 = ~v_4440;
  assign v_4454 = mux_4454(v_4455);
  assign v_4455 = ~v_4450;
  pebbles_core
    pebbles_core_4456
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4457),
       .in0_consume_en(vin0_consume_en_4456),
       .out_canPeek(vout_canPeek_4456),
       .out_peek(vout_peek_4456));
  assign v_4457 = v_4458 | v_4459;
  assign v_4458 = mux_4458(v_4444);
  assign v_4459 = mux_4459(v_4460);
  assign v_4460 = ~v_4444;
  assign v_4461 = v_4462 & 1'h1;
  assign v_4462 = v_4463 & v_4464;
  assign v_4463 = ~act_4443;
  assign v_4464 = v_4465 | v_4473;
  assign v_4465 = v_4466 | v_4471;
  assign v_4466 = mux_4466(v_4467);
  assign v_4467 = v_4440 & v_4468;
  assign v_4468 = v_4469 & 1'h1;
  assign v_4469 = v_4470 | 1'h0;
  assign v_4470 = ~v_4433;
  assign v_4471 = mux_4471(v_4472);
  assign v_4472 = ~v_4467;
  assign v_4473 = ~v_4440;
  assign v_4474 = v_4475 | v_4476;
  assign v_4475 = mux_4475(v_4442);
  assign v_4476 = mux_4476(v_4461);
  assign v_4478 = v_4479 | v_4498;
  assign v_4479 = act_4480 & 1'h1;
  assign act_4480 = v_4481 | v_4487;
  assign v_4481 = v_4482 & v_4488;
  assign v_4482 = v_4483 & vout_canPeek_4493;
  assign v_4483 = ~vout_canPeek_4484;
  pebbles_core
    pebbles_core_4484
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4485),
       .in0_consume_en(vin0_consume_en_4484),
       .out_canPeek(vout_canPeek_4484),
       .out_peek(vout_peek_4484));
  assign v_4485 = v_4486 | v_4491;
  assign v_4486 = mux_4486(v_4487);
  assign v_4487 = vout_canPeek_4484 & v_4488;
  assign v_4488 = v_4489 & 1'h1;
  assign v_4489 = v_4490 | 1'h0;
  assign v_4490 = ~v_4477;
  assign v_4491 = mux_4491(v_4492);
  assign v_4492 = ~v_4487;
  pebbles_core
    pebbles_core_4493
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4494),
       .in0_consume_en(vin0_consume_en_4493),
       .out_canPeek(vout_canPeek_4493),
       .out_peek(vout_peek_4493));
  assign v_4494 = v_4495 | v_4496;
  assign v_4495 = mux_4495(v_4481);
  assign v_4496 = mux_4496(v_4497);
  assign v_4497 = ~v_4481;
  assign v_4498 = v_4499 & 1'h1;
  assign v_4499 = v_4500 & v_4501;
  assign v_4500 = ~act_4480;
  assign v_4501 = v_4502 | v_4506;
  assign v_4502 = v_4503 | v_4504;
  assign v_4503 = mux_4503(v_4437);
  assign v_4504 = mux_4504(v_4505);
  assign v_4505 = ~v_4437;
  assign v_4506 = ~v_4477;
  assign v_4507 = v_4508 | v_4509;
  assign v_4508 = mux_4508(v_4479);
  assign v_4509 = mux_4509(v_4498);
  assign v_4510 = v_4511 & 1'h1;
  assign v_4511 = v_4512 & v_4513;
  assign v_4512 = ~act_4436;
  assign v_4513 = v_4514 | v_4522;
  assign v_4514 = v_4515 | v_4520;
  assign v_4515 = mux_4515(v_4516);
  assign v_4516 = v_4433 & v_4517;
  assign v_4517 = v_4518 & 1'h1;
  assign v_4518 = v_4519 | 1'h0;
  assign v_4519 = ~v_4426;
  assign v_4520 = mux_4520(v_4521);
  assign v_4521 = ~v_4516;
  assign v_4522 = ~v_4433;
  assign v_4523 = v_4524 | v_4525;
  assign v_4524 = mux_4524(v_4435);
  assign v_4525 = mux_4525(v_4510);
  assign v_4527 = v_4528 | v_4603;
  assign v_4528 = act_4529 & 1'h1;
  assign act_4529 = v_4530 | v_4560;
  assign v_4530 = v_4531 & v_4561;
  assign v_4531 = v_4532 & v_4570;
  assign v_4532 = ~v_4533;
  assign v_4534 = v_4535 | v_4554;
  assign v_4535 = act_4536 & 1'h1;
  assign act_4536 = v_4537 | v_4543;
  assign v_4537 = v_4538 & v_4544;
  assign v_4538 = v_4539 & vout_canPeek_4549;
  assign v_4539 = ~vout_canPeek_4540;
  pebbles_core
    pebbles_core_4540
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4541),
       .in0_consume_en(vin0_consume_en_4540),
       .out_canPeek(vout_canPeek_4540),
       .out_peek(vout_peek_4540));
  assign v_4541 = v_4542 | v_4547;
  assign v_4542 = mux_4542(v_4543);
  assign v_4543 = vout_canPeek_4540 & v_4544;
  assign v_4544 = v_4545 & 1'h1;
  assign v_4545 = v_4546 | 1'h0;
  assign v_4546 = ~v_4533;
  assign v_4547 = mux_4547(v_4548);
  assign v_4548 = ~v_4543;
  pebbles_core
    pebbles_core_4549
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4550),
       .in0_consume_en(vin0_consume_en_4549),
       .out_canPeek(vout_canPeek_4549),
       .out_peek(vout_peek_4549));
  assign v_4550 = v_4551 | v_4552;
  assign v_4551 = mux_4551(v_4537);
  assign v_4552 = mux_4552(v_4553);
  assign v_4553 = ~v_4537;
  assign v_4554 = v_4555 & 1'h1;
  assign v_4555 = v_4556 & v_4557;
  assign v_4556 = ~act_4536;
  assign v_4557 = v_4558 | v_4566;
  assign v_4558 = v_4559 | v_4564;
  assign v_4559 = mux_4559(v_4560);
  assign v_4560 = v_4533 & v_4561;
  assign v_4561 = v_4562 & 1'h1;
  assign v_4562 = v_4563 | 1'h0;
  assign v_4563 = ~v_4526;
  assign v_4564 = mux_4564(v_4565);
  assign v_4565 = ~v_4560;
  assign v_4566 = ~v_4533;
  assign v_4567 = v_4568 | v_4569;
  assign v_4568 = mux_4568(v_4535);
  assign v_4569 = mux_4569(v_4554);
  assign v_4571 = v_4572 | v_4591;
  assign v_4572 = act_4573 & 1'h1;
  assign act_4573 = v_4574 | v_4580;
  assign v_4574 = v_4575 & v_4581;
  assign v_4575 = v_4576 & vout_canPeek_4586;
  assign v_4576 = ~vout_canPeek_4577;
  pebbles_core
    pebbles_core_4577
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4578),
       .in0_consume_en(vin0_consume_en_4577),
       .out_canPeek(vout_canPeek_4577),
       .out_peek(vout_peek_4577));
  assign v_4578 = v_4579 | v_4584;
  assign v_4579 = mux_4579(v_4580);
  assign v_4580 = vout_canPeek_4577 & v_4581;
  assign v_4581 = v_4582 & 1'h1;
  assign v_4582 = v_4583 | 1'h0;
  assign v_4583 = ~v_4570;
  assign v_4584 = mux_4584(v_4585);
  assign v_4585 = ~v_4580;
  pebbles_core
    pebbles_core_4586
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4587),
       .in0_consume_en(vin0_consume_en_4586),
       .out_canPeek(vout_canPeek_4586),
       .out_peek(vout_peek_4586));
  assign v_4587 = v_4588 | v_4589;
  assign v_4588 = mux_4588(v_4574);
  assign v_4589 = mux_4589(v_4590);
  assign v_4590 = ~v_4574;
  assign v_4591 = v_4592 & 1'h1;
  assign v_4592 = v_4593 & v_4594;
  assign v_4593 = ~act_4573;
  assign v_4594 = v_4595 | v_4599;
  assign v_4595 = v_4596 | v_4597;
  assign v_4596 = mux_4596(v_4530);
  assign v_4597 = mux_4597(v_4598);
  assign v_4598 = ~v_4530;
  assign v_4599 = ~v_4570;
  assign v_4600 = v_4601 | v_4602;
  assign v_4601 = mux_4601(v_4572);
  assign v_4602 = mux_4602(v_4591);
  assign v_4603 = v_4604 & 1'h1;
  assign v_4604 = v_4605 & v_4606;
  assign v_4605 = ~act_4529;
  assign v_4606 = v_4607 | v_4611;
  assign v_4607 = v_4608 | v_4609;
  assign v_4608 = mux_4608(v_4430);
  assign v_4609 = mux_4609(v_4610);
  assign v_4610 = ~v_4430;
  assign v_4611 = ~v_4526;
  assign v_4612 = v_4613 | v_4614;
  assign v_4613 = mux_4613(v_4528);
  assign v_4614 = mux_4614(v_4603);
  assign v_4615 = v_4616 & 1'h1;
  assign v_4616 = v_4617 & v_4618;
  assign v_4617 = ~act_4429;
  assign v_4618 = v_4619 | v_4627;
  assign v_4619 = v_4620 | v_4625;
  assign v_4620 = mux_4620(v_4621);
  assign v_4621 = v_4426 & v_4622;
  assign v_4622 = v_4623 & 1'h1;
  assign v_4623 = v_4624 | 1'h0;
  assign v_4624 = ~v_4419;
  assign v_4625 = mux_4625(v_4626);
  assign v_4626 = ~v_4621;
  assign v_4627 = ~v_4426;
  assign v_4628 = v_4629 | v_4630;
  assign v_4629 = mux_4629(v_4428);
  assign v_4630 = mux_4630(v_4615);
  assign v_4632 = v_4633 | v_4820;
  assign v_4633 = act_4634 & 1'h1;
  assign act_4634 = v_4635 | v_4721;
  assign v_4635 = v_4636 & v_4722;
  assign v_4636 = v_4637 & v_4731;
  assign v_4637 = ~v_4638;
  assign v_4639 = v_4640 | v_4715;
  assign v_4640 = act_4641 & 1'h1;
  assign act_4641 = v_4642 | v_4672;
  assign v_4642 = v_4643 & v_4673;
  assign v_4643 = v_4644 & v_4682;
  assign v_4644 = ~v_4645;
  assign v_4646 = v_4647 | v_4666;
  assign v_4647 = act_4648 & 1'h1;
  assign act_4648 = v_4649 | v_4655;
  assign v_4649 = v_4650 & v_4656;
  assign v_4650 = v_4651 & vout_canPeek_4661;
  assign v_4651 = ~vout_canPeek_4652;
  pebbles_core
    pebbles_core_4652
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4653),
       .in0_consume_en(vin0_consume_en_4652),
       .out_canPeek(vout_canPeek_4652),
       .out_peek(vout_peek_4652));
  assign v_4653 = v_4654 | v_4659;
  assign v_4654 = mux_4654(v_4655);
  assign v_4655 = vout_canPeek_4652 & v_4656;
  assign v_4656 = v_4657 & 1'h1;
  assign v_4657 = v_4658 | 1'h0;
  assign v_4658 = ~v_4645;
  assign v_4659 = mux_4659(v_4660);
  assign v_4660 = ~v_4655;
  pebbles_core
    pebbles_core_4661
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4662),
       .in0_consume_en(vin0_consume_en_4661),
       .out_canPeek(vout_canPeek_4661),
       .out_peek(vout_peek_4661));
  assign v_4662 = v_4663 | v_4664;
  assign v_4663 = mux_4663(v_4649);
  assign v_4664 = mux_4664(v_4665);
  assign v_4665 = ~v_4649;
  assign v_4666 = v_4667 & 1'h1;
  assign v_4667 = v_4668 & v_4669;
  assign v_4668 = ~act_4648;
  assign v_4669 = v_4670 | v_4678;
  assign v_4670 = v_4671 | v_4676;
  assign v_4671 = mux_4671(v_4672);
  assign v_4672 = v_4645 & v_4673;
  assign v_4673 = v_4674 & 1'h1;
  assign v_4674 = v_4675 | 1'h0;
  assign v_4675 = ~v_4638;
  assign v_4676 = mux_4676(v_4677);
  assign v_4677 = ~v_4672;
  assign v_4678 = ~v_4645;
  assign v_4679 = v_4680 | v_4681;
  assign v_4680 = mux_4680(v_4647);
  assign v_4681 = mux_4681(v_4666);
  assign v_4683 = v_4684 | v_4703;
  assign v_4684 = act_4685 & 1'h1;
  assign act_4685 = v_4686 | v_4692;
  assign v_4686 = v_4687 & v_4693;
  assign v_4687 = v_4688 & vout_canPeek_4698;
  assign v_4688 = ~vout_canPeek_4689;
  pebbles_core
    pebbles_core_4689
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4690),
       .in0_consume_en(vin0_consume_en_4689),
       .out_canPeek(vout_canPeek_4689),
       .out_peek(vout_peek_4689));
  assign v_4690 = v_4691 | v_4696;
  assign v_4691 = mux_4691(v_4692);
  assign v_4692 = vout_canPeek_4689 & v_4693;
  assign v_4693 = v_4694 & 1'h1;
  assign v_4694 = v_4695 | 1'h0;
  assign v_4695 = ~v_4682;
  assign v_4696 = mux_4696(v_4697);
  assign v_4697 = ~v_4692;
  pebbles_core
    pebbles_core_4698
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4699),
       .in0_consume_en(vin0_consume_en_4698),
       .out_canPeek(vout_canPeek_4698),
       .out_peek(vout_peek_4698));
  assign v_4699 = v_4700 | v_4701;
  assign v_4700 = mux_4700(v_4686);
  assign v_4701 = mux_4701(v_4702);
  assign v_4702 = ~v_4686;
  assign v_4703 = v_4704 & 1'h1;
  assign v_4704 = v_4705 & v_4706;
  assign v_4705 = ~act_4685;
  assign v_4706 = v_4707 | v_4711;
  assign v_4707 = v_4708 | v_4709;
  assign v_4708 = mux_4708(v_4642);
  assign v_4709 = mux_4709(v_4710);
  assign v_4710 = ~v_4642;
  assign v_4711 = ~v_4682;
  assign v_4712 = v_4713 | v_4714;
  assign v_4713 = mux_4713(v_4684);
  assign v_4714 = mux_4714(v_4703);
  assign v_4715 = v_4716 & 1'h1;
  assign v_4716 = v_4717 & v_4718;
  assign v_4717 = ~act_4641;
  assign v_4718 = v_4719 | v_4727;
  assign v_4719 = v_4720 | v_4725;
  assign v_4720 = mux_4720(v_4721);
  assign v_4721 = v_4638 & v_4722;
  assign v_4722 = v_4723 & 1'h1;
  assign v_4723 = v_4724 | 1'h0;
  assign v_4724 = ~v_4631;
  assign v_4725 = mux_4725(v_4726);
  assign v_4726 = ~v_4721;
  assign v_4727 = ~v_4638;
  assign v_4728 = v_4729 | v_4730;
  assign v_4729 = mux_4729(v_4640);
  assign v_4730 = mux_4730(v_4715);
  assign v_4732 = v_4733 | v_4808;
  assign v_4733 = act_4734 & 1'h1;
  assign act_4734 = v_4735 | v_4765;
  assign v_4735 = v_4736 & v_4766;
  assign v_4736 = v_4737 & v_4775;
  assign v_4737 = ~v_4738;
  assign v_4739 = v_4740 | v_4759;
  assign v_4740 = act_4741 & 1'h1;
  assign act_4741 = v_4742 | v_4748;
  assign v_4742 = v_4743 & v_4749;
  assign v_4743 = v_4744 & vout_canPeek_4754;
  assign v_4744 = ~vout_canPeek_4745;
  pebbles_core
    pebbles_core_4745
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4746),
       .in0_consume_en(vin0_consume_en_4745),
       .out_canPeek(vout_canPeek_4745),
       .out_peek(vout_peek_4745));
  assign v_4746 = v_4747 | v_4752;
  assign v_4747 = mux_4747(v_4748);
  assign v_4748 = vout_canPeek_4745 & v_4749;
  assign v_4749 = v_4750 & 1'h1;
  assign v_4750 = v_4751 | 1'h0;
  assign v_4751 = ~v_4738;
  assign v_4752 = mux_4752(v_4753);
  assign v_4753 = ~v_4748;
  pebbles_core
    pebbles_core_4754
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4755),
       .in0_consume_en(vin0_consume_en_4754),
       .out_canPeek(vout_canPeek_4754),
       .out_peek(vout_peek_4754));
  assign v_4755 = v_4756 | v_4757;
  assign v_4756 = mux_4756(v_4742);
  assign v_4757 = mux_4757(v_4758);
  assign v_4758 = ~v_4742;
  assign v_4759 = v_4760 & 1'h1;
  assign v_4760 = v_4761 & v_4762;
  assign v_4761 = ~act_4741;
  assign v_4762 = v_4763 | v_4771;
  assign v_4763 = v_4764 | v_4769;
  assign v_4764 = mux_4764(v_4765);
  assign v_4765 = v_4738 & v_4766;
  assign v_4766 = v_4767 & 1'h1;
  assign v_4767 = v_4768 | 1'h0;
  assign v_4768 = ~v_4731;
  assign v_4769 = mux_4769(v_4770);
  assign v_4770 = ~v_4765;
  assign v_4771 = ~v_4738;
  assign v_4772 = v_4773 | v_4774;
  assign v_4773 = mux_4773(v_4740);
  assign v_4774 = mux_4774(v_4759);
  assign v_4776 = v_4777 | v_4796;
  assign v_4777 = act_4778 & 1'h1;
  assign act_4778 = v_4779 | v_4785;
  assign v_4779 = v_4780 & v_4786;
  assign v_4780 = v_4781 & vout_canPeek_4791;
  assign v_4781 = ~vout_canPeek_4782;
  pebbles_core
    pebbles_core_4782
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4783),
       .in0_consume_en(vin0_consume_en_4782),
       .out_canPeek(vout_canPeek_4782),
       .out_peek(vout_peek_4782));
  assign v_4783 = v_4784 | v_4789;
  assign v_4784 = mux_4784(v_4785);
  assign v_4785 = vout_canPeek_4782 & v_4786;
  assign v_4786 = v_4787 & 1'h1;
  assign v_4787 = v_4788 | 1'h0;
  assign v_4788 = ~v_4775;
  assign v_4789 = mux_4789(v_4790);
  assign v_4790 = ~v_4785;
  pebbles_core
    pebbles_core_4791
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4792),
       .in0_consume_en(vin0_consume_en_4791),
       .out_canPeek(vout_canPeek_4791),
       .out_peek(vout_peek_4791));
  assign v_4792 = v_4793 | v_4794;
  assign v_4793 = mux_4793(v_4779);
  assign v_4794 = mux_4794(v_4795);
  assign v_4795 = ~v_4779;
  assign v_4796 = v_4797 & 1'h1;
  assign v_4797 = v_4798 & v_4799;
  assign v_4798 = ~act_4778;
  assign v_4799 = v_4800 | v_4804;
  assign v_4800 = v_4801 | v_4802;
  assign v_4801 = mux_4801(v_4735);
  assign v_4802 = mux_4802(v_4803);
  assign v_4803 = ~v_4735;
  assign v_4804 = ~v_4775;
  assign v_4805 = v_4806 | v_4807;
  assign v_4806 = mux_4806(v_4777);
  assign v_4807 = mux_4807(v_4796);
  assign v_4808 = v_4809 & 1'h1;
  assign v_4809 = v_4810 & v_4811;
  assign v_4810 = ~act_4734;
  assign v_4811 = v_4812 | v_4816;
  assign v_4812 = v_4813 | v_4814;
  assign v_4813 = mux_4813(v_4635);
  assign v_4814 = mux_4814(v_4815);
  assign v_4815 = ~v_4635;
  assign v_4816 = ~v_4731;
  assign v_4817 = v_4818 | v_4819;
  assign v_4818 = mux_4818(v_4733);
  assign v_4819 = mux_4819(v_4808);
  assign v_4820 = v_4821 & 1'h1;
  assign v_4821 = v_4822 & v_4823;
  assign v_4822 = ~act_4634;
  assign v_4823 = v_4824 | v_4828;
  assign v_4824 = v_4825 | v_4826;
  assign v_4825 = mux_4825(v_4423);
  assign v_4826 = mux_4826(v_4827);
  assign v_4827 = ~v_4423;
  assign v_4828 = ~v_4631;
  assign v_4829 = v_4830 | v_4831;
  assign v_4830 = mux_4830(v_4633);
  assign v_4831 = mux_4831(v_4820);
  assign v_4832 = v_4833 & 1'h1;
  assign v_4833 = v_4834 & v_4835;
  assign v_4834 = ~act_4422;
  assign v_4835 = v_4836 | v_4844;
  assign v_4836 = v_4837 | v_4842;
  assign v_4837 = mux_4837(v_4838);
  assign v_4838 = v_4419 & v_4839;
  assign v_4839 = v_4840 & 1'h1;
  assign v_4840 = v_4841 | 1'h0;
  assign v_4841 = ~v_4412;
  assign v_4842 = mux_4842(v_4843);
  assign v_4843 = ~v_4838;
  assign v_4844 = ~v_4419;
  assign v_4845 = v_4846 | v_4847;
  assign v_4846 = mux_4846(v_4421);
  assign v_4847 = mux_4847(v_4832);
  assign v_4849 = v_4850 | v_5261;
  assign v_4850 = act_4851 & 1'h1;
  assign act_4851 = v_4852 | v_5050;
  assign v_4852 = v_4853 & v_5051;
  assign v_4853 = v_4854 & v_5060;
  assign v_4854 = ~v_4855;
  assign v_4856 = v_4857 | v_5044;
  assign v_4857 = act_4858 & 1'h1;
  assign act_4858 = v_4859 | v_4945;
  assign v_4859 = v_4860 & v_4946;
  assign v_4860 = v_4861 & v_4955;
  assign v_4861 = ~v_4862;
  assign v_4863 = v_4864 | v_4939;
  assign v_4864 = act_4865 & 1'h1;
  assign act_4865 = v_4866 | v_4896;
  assign v_4866 = v_4867 & v_4897;
  assign v_4867 = v_4868 & v_4906;
  assign v_4868 = ~v_4869;
  assign v_4870 = v_4871 | v_4890;
  assign v_4871 = act_4872 & 1'h1;
  assign act_4872 = v_4873 | v_4879;
  assign v_4873 = v_4874 & v_4880;
  assign v_4874 = v_4875 & vout_canPeek_4885;
  assign v_4875 = ~vout_canPeek_4876;
  pebbles_core
    pebbles_core_4876
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4877),
       .in0_consume_en(vin0_consume_en_4876),
       .out_canPeek(vout_canPeek_4876),
       .out_peek(vout_peek_4876));
  assign v_4877 = v_4878 | v_4883;
  assign v_4878 = mux_4878(v_4879);
  assign v_4879 = vout_canPeek_4876 & v_4880;
  assign v_4880 = v_4881 & 1'h1;
  assign v_4881 = v_4882 | 1'h0;
  assign v_4882 = ~v_4869;
  assign v_4883 = mux_4883(v_4884);
  assign v_4884 = ~v_4879;
  pebbles_core
    pebbles_core_4885
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4886),
       .in0_consume_en(vin0_consume_en_4885),
       .out_canPeek(vout_canPeek_4885),
       .out_peek(vout_peek_4885));
  assign v_4886 = v_4887 | v_4888;
  assign v_4887 = mux_4887(v_4873);
  assign v_4888 = mux_4888(v_4889);
  assign v_4889 = ~v_4873;
  assign v_4890 = v_4891 & 1'h1;
  assign v_4891 = v_4892 & v_4893;
  assign v_4892 = ~act_4872;
  assign v_4893 = v_4894 | v_4902;
  assign v_4894 = v_4895 | v_4900;
  assign v_4895 = mux_4895(v_4896);
  assign v_4896 = v_4869 & v_4897;
  assign v_4897 = v_4898 & 1'h1;
  assign v_4898 = v_4899 | 1'h0;
  assign v_4899 = ~v_4862;
  assign v_4900 = mux_4900(v_4901);
  assign v_4901 = ~v_4896;
  assign v_4902 = ~v_4869;
  assign v_4903 = v_4904 | v_4905;
  assign v_4904 = mux_4904(v_4871);
  assign v_4905 = mux_4905(v_4890);
  assign v_4907 = v_4908 | v_4927;
  assign v_4908 = act_4909 & 1'h1;
  assign act_4909 = v_4910 | v_4916;
  assign v_4910 = v_4911 & v_4917;
  assign v_4911 = v_4912 & vout_canPeek_4922;
  assign v_4912 = ~vout_canPeek_4913;
  pebbles_core
    pebbles_core_4913
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4914),
       .in0_consume_en(vin0_consume_en_4913),
       .out_canPeek(vout_canPeek_4913),
       .out_peek(vout_peek_4913));
  assign v_4914 = v_4915 | v_4920;
  assign v_4915 = mux_4915(v_4916);
  assign v_4916 = vout_canPeek_4913 & v_4917;
  assign v_4917 = v_4918 & 1'h1;
  assign v_4918 = v_4919 | 1'h0;
  assign v_4919 = ~v_4906;
  assign v_4920 = mux_4920(v_4921);
  assign v_4921 = ~v_4916;
  pebbles_core
    pebbles_core_4922
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4923),
       .in0_consume_en(vin0_consume_en_4922),
       .out_canPeek(vout_canPeek_4922),
       .out_peek(vout_peek_4922));
  assign v_4923 = v_4924 | v_4925;
  assign v_4924 = mux_4924(v_4910);
  assign v_4925 = mux_4925(v_4926);
  assign v_4926 = ~v_4910;
  assign v_4927 = v_4928 & 1'h1;
  assign v_4928 = v_4929 & v_4930;
  assign v_4929 = ~act_4909;
  assign v_4930 = v_4931 | v_4935;
  assign v_4931 = v_4932 | v_4933;
  assign v_4932 = mux_4932(v_4866);
  assign v_4933 = mux_4933(v_4934);
  assign v_4934 = ~v_4866;
  assign v_4935 = ~v_4906;
  assign v_4936 = v_4937 | v_4938;
  assign v_4937 = mux_4937(v_4908);
  assign v_4938 = mux_4938(v_4927);
  assign v_4939 = v_4940 & 1'h1;
  assign v_4940 = v_4941 & v_4942;
  assign v_4941 = ~act_4865;
  assign v_4942 = v_4943 | v_4951;
  assign v_4943 = v_4944 | v_4949;
  assign v_4944 = mux_4944(v_4945);
  assign v_4945 = v_4862 & v_4946;
  assign v_4946 = v_4947 & 1'h1;
  assign v_4947 = v_4948 | 1'h0;
  assign v_4948 = ~v_4855;
  assign v_4949 = mux_4949(v_4950);
  assign v_4950 = ~v_4945;
  assign v_4951 = ~v_4862;
  assign v_4952 = v_4953 | v_4954;
  assign v_4953 = mux_4953(v_4864);
  assign v_4954 = mux_4954(v_4939);
  assign v_4956 = v_4957 | v_5032;
  assign v_4957 = act_4958 & 1'h1;
  assign act_4958 = v_4959 | v_4989;
  assign v_4959 = v_4960 & v_4990;
  assign v_4960 = v_4961 & v_4999;
  assign v_4961 = ~v_4962;
  assign v_4963 = v_4964 | v_4983;
  assign v_4964 = act_4965 & 1'h1;
  assign act_4965 = v_4966 | v_4972;
  assign v_4966 = v_4967 & v_4973;
  assign v_4967 = v_4968 & vout_canPeek_4978;
  assign v_4968 = ~vout_canPeek_4969;
  pebbles_core
    pebbles_core_4969
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4970),
       .in0_consume_en(vin0_consume_en_4969),
       .out_canPeek(vout_canPeek_4969),
       .out_peek(vout_peek_4969));
  assign v_4970 = v_4971 | v_4976;
  assign v_4971 = mux_4971(v_4972);
  assign v_4972 = vout_canPeek_4969 & v_4973;
  assign v_4973 = v_4974 & 1'h1;
  assign v_4974 = v_4975 | 1'h0;
  assign v_4975 = ~v_4962;
  assign v_4976 = mux_4976(v_4977);
  assign v_4977 = ~v_4972;
  pebbles_core
    pebbles_core_4978
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_4979),
       .in0_consume_en(vin0_consume_en_4978),
       .out_canPeek(vout_canPeek_4978),
       .out_peek(vout_peek_4978));
  assign v_4979 = v_4980 | v_4981;
  assign v_4980 = mux_4980(v_4966);
  assign v_4981 = mux_4981(v_4982);
  assign v_4982 = ~v_4966;
  assign v_4983 = v_4984 & 1'h1;
  assign v_4984 = v_4985 & v_4986;
  assign v_4985 = ~act_4965;
  assign v_4986 = v_4987 | v_4995;
  assign v_4987 = v_4988 | v_4993;
  assign v_4988 = mux_4988(v_4989);
  assign v_4989 = v_4962 & v_4990;
  assign v_4990 = v_4991 & 1'h1;
  assign v_4991 = v_4992 | 1'h0;
  assign v_4992 = ~v_4955;
  assign v_4993 = mux_4993(v_4994);
  assign v_4994 = ~v_4989;
  assign v_4995 = ~v_4962;
  assign v_4996 = v_4997 | v_4998;
  assign v_4997 = mux_4997(v_4964);
  assign v_4998 = mux_4998(v_4983);
  assign v_5000 = v_5001 | v_5020;
  assign v_5001 = act_5002 & 1'h1;
  assign act_5002 = v_5003 | v_5009;
  assign v_5003 = v_5004 & v_5010;
  assign v_5004 = v_5005 & vout_canPeek_5015;
  assign v_5005 = ~vout_canPeek_5006;
  pebbles_core
    pebbles_core_5006
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5007),
       .in0_consume_en(vin0_consume_en_5006),
       .out_canPeek(vout_canPeek_5006),
       .out_peek(vout_peek_5006));
  assign v_5007 = v_5008 | v_5013;
  assign v_5008 = mux_5008(v_5009);
  assign v_5009 = vout_canPeek_5006 & v_5010;
  assign v_5010 = v_5011 & 1'h1;
  assign v_5011 = v_5012 | 1'h0;
  assign v_5012 = ~v_4999;
  assign v_5013 = mux_5013(v_5014);
  assign v_5014 = ~v_5009;
  pebbles_core
    pebbles_core_5015
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5016),
       .in0_consume_en(vin0_consume_en_5015),
       .out_canPeek(vout_canPeek_5015),
       .out_peek(vout_peek_5015));
  assign v_5016 = v_5017 | v_5018;
  assign v_5017 = mux_5017(v_5003);
  assign v_5018 = mux_5018(v_5019);
  assign v_5019 = ~v_5003;
  assign v_5020 = v_5021 & 1'h1;
  assign v_5021 = v_5022 & v_5023;
  assign v_5022 = ~act_5002;
  assign v_5023 = v_5024 | v_5028;
  assign v_5024 = v_5025 | v_5026;
  assign v_5025 = mux_5025(v_4959);
  assign v_5026 = mux_5026(v_5027);
  assign v_5027 = ~v_4959;
  assign v_5028 = ~v_4999;
  assign v_5029 = v_5030 | v_5031;
  assign v_5030 = mux_5030(v_5001);
  assign v_5031 = mux_5031(v_5020);
  assign v_5032 = v_5033 & 1'h1;
  assign v_5033 = v_5034 & v_5035;
  assign v_5034 = ~act_4958;
  assign v_5035 = v_5036 | v_5040;
  assign v_5036 = v_5037 | v_5038;
  assign v_5037 = mux_5037(v_4859);
  assign v_5038 = mux_5038(v_5039);
  assign v_5039 = ~v_4859;
  assign v_5040 = ~v_4955;
  assign v_5041 = v_5042 | v_5043;
  assign v_5042 = mux_5042(v_4957);
  assign v_5043 = mux_5043(v_5032);
  assign v_5044 = v_5045 & 1'h1;
  assign v_5045 = v_5046 & v_5047;
  assign v_5046 = ~act_4858;
  assign v_5047 = v_5048 | v_5056;
  assign v_5048 = v_5049 | v_5054;
  assign v_5049 = mux_5049(v_5050);
  assign v_5050 = v_4855 & v_5051;
  assign v_5051 = v_5052 & 1'h1;
  assign v_5052 = v_5053 | 1'h0;
  assign v_5053 = ~v_4848;
  assign v_5054 = mux_5054(v_5055);
  assign v_5055 = ~v_5050;
  assign v_5056 = ~v_4855;
  assign v_5057 = v_5058 | v_5059;
  assign v_5058 = mux_5058(v_4857);
  assign v_5059 = mux_5059(v_5044);
  assign v_5061 = v_5062 | v_5249;
  assign v_5062 = act_5063 & 1'h1;
  assign act_5063 = v_5064 | v_5150;
  assign v_5064 = v_5065 & v_5151;
  assign v_5065 = v_5066 & v_5160;
  assign v_5066 = ~v_5067;
  assign v_5068 = v_5069 | v_5144;
  assign v_5069 = act_5070 & 1'h1;
  assign act_5070 = v_5071 | v_5101;
  assign v_5071 = v_5072 & v_5102;
  assign v_5072 = v_5073 & v_5111;
  assign v_5073 = ~v_5074;
  assign v_5075 = v_5076 | v_5095;
  assign v_5076 = act_5077 & 1'h1;
  assign act_5077 = v_5078 | v_5084;
  assign v_5078 = v_5079 & v_5085;
  assign v_5079 = v_5080 & vout_canPeek_5090;
  assign v_5080 = ~vout_canPeek_5081;
  pebbles_core
    pebbles_core_5081
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5082),
       .in0_consume_en(vin0_consume_en_5081),
       .out_canPeek(vout_canPeek_5081),
       .out_peek(vout_peek_5081));
  assign v_5082 = v_5083 | v_5088;
  assign v_5083 = mux_5083(v_5084);
  assign v_5084 = vout_canPeek_5081 & v_5085;
  assign v_5085 = v_5086 & 1'h1;
  assign v_5086 = v_5087 | 1'h0;
  assign v_5087 = ~v_5074;
  assign v_5088 = mux_5088(v_5089);
  assign v_5089 = ~v_5084;
  pebbles_core
    pebbles_core_5090
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5091),
       .in0_consume_en(vin0_consume_en_5090),
       .out_canPeek(vout_canPeek_5090),
       .out_peek(vout_peek_5090));
  assign v_5091 = v_5092 | v_5093;
  assign v_5092 = mux_5092(v_5078);
  assign v_5093 = mux_5093(v_5094);
  assign v_5094 = ~v_5078;
  assign v_5095 = v_5096 & 1'h1;
  assign v_5096 = v_5097 & v_5098;
  assign v_5097 = ~act_5077;
  assign v_5098 = v_5099 | v_5107;
  assign v_5099 = v_5100 | v_5105;
  assign v_5100 = mux_5100(v_5101);
  assign v_5101 = v_5074 & v_5102;
  assign v_5102 = v_5103 & 1'h1;
  assign v_5103 = v_5104 | 1'h0;
  assign v_5104 = ~v_5067;
  assign v_5105 = mux_5105(v_5106);
  assign v_5106 = ~v_5101;
  assign v_5107 = ~v_5074;
  assign v_5108 = v_5109 | v_5110;
  assign v_5109 = mux_5109(v_5076);
  assign v_5110 = mux_5110(v_5095);
  assign v_5112 = v_5113 | v_5132;
  assign v_5113 = act_5114 & 1'h1;
  assign act_5114 = v_5115 | v_5121;
  assign v_5115 = v_5116 & v_5122;
  assign v_5116 = v_5117 & vout_canPeek_5127;
  assign v_5117 = ~vout_canPeek_5118;
  pebbles_core
    pebbles_core_5118
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5119),
       .in0_consume_en(vin0_consume_en_5118),
       .out_canPeek(vout_canPeek_5118),
       .out_peek(vout_peek_5118));
  assign v_5119 = v_5120 | v_5125;
  assign v_5120 = mux_5120(v_5121);
  assign v_5121 = vout_canPeek_5118 & v_5122;
  assign v_5122 = v_5123 & 1'h1;
  assign v_5123 = v_5124 | 1'h0;
  assign v_5124 = ~v_5111;
  assign v_5125 = mux_5125(v_5126);
  assign v_5126 = ~v_5121;
  pebbles_core
    pebbles_core_5127
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5128),
       .in0_consume_en(vin0_consume_en_5127),
       .out_canPeek(vout_canPeek_5127),
       .out_peek(vout_peek_5127));
  assign v_5128 = v_5129 | v_5130;
  assign v_5129 = mux_5129(v_5115);
  assign v_5130 = mux_5130(v_5131);
  assign v_5131 = ~v_5115;
  assign v_5132 = v_5133 & 1'h1;
  assign v_5133 = v_5134 & v_5135;
  assign v_5134 = ~act_5114;
  assign v_5135 = v_5136 | v_5140;
  assign v_5136 = v_5137 | v_5138;
  assign v_5137 = mux_5137(v_5071);
  assign v_5138 = mux_5138(v_5139);
  assign v_5139 = ~v_5071;
  assign v_5140 = ~v_5111;
  assign v_5141 = v_5142 | v_5143;
  assign v_5142 = mux_5142(v_5113);
  assign v_5143 = mux_5143(v_5132);
  assign v_5144 = v_5145 & 1'h1;
  assign v_5145 = v_5146 & v_5147;
  assign v_5146 = ~act_5070;
  assign v_5147 = v_5148 | v_5156;
  assign v_5148 = v_5149 | v_5154;
  assign v_5149 = mux_5149(v_5150);
  assign v_5150 = v_5067 & v_5151;
  assign v_5151 = v_5152 & 1'h1;
  assign v_5152 = v_5153 | 1'h0;
  assign v_5153 = ~v_5060;
  assign v_5154 = mux_5154(v_5155);
  assign v_5155 = ~v_5150;
  assign v_5156 = ~v_5067;
  assign v_5157 = v_5158 | v_5159;
  assign v_5158 = mux_5158(v_5069);
  assign v_5159 = mux_5159(v_5144);
  assign v_5161 = v_5162 | v_5237;
  assign v_5162 = act_5163 & 1'h1;
  assign act_5163 = v_5164 | v_5194;
  assign v_5164 = v_5165 & v_5195;
  assign v_5165 = v_5166 & v_5204;
  assign v_5166 = ~v_5167;
  assign v_5168 = v_5169 | v_5188;
  assign v_5169 = act_5170 & 1'h1;
  assign act_5170 = v_5171 | v_5177;
  assign v_5171 = v_5172 & v_5178;
  assign v_5172 = v_5173 & vout_canPeek_5183;
  assign v_5173 = ~vout_canPeek_5174;
  pebbles_core
    pebbles_core_5174
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5175),
       .in0_consume_en(vin0_consume_en_5174),
       .out_canPeek(vout_canPeek_5174),
       .out_peek(vout_peek_5174));
  assign v_5175 = v_5176 | v_5181;
  assign v_5176 = mux_5176(v_5177);
  assign v_5177 = vout_canPeek_5174 & v_5178;
  assign v_5178 = v_5179 & 1'h1;
  assign v_5179 = v_5180 | 1'h0;
  assign v_5180 = ~v_5167;
  assign v_5181 = mux_5181(v_5182);
  assign v_5182 = ~v_5177;
  pebbles_core
    pebbles_core_5183
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5184),
       .in0_consume_en(vin0_consume_en_5183),
       .out_canPeek(vout_canPeek_5183),
       .out_peek(vout_peek_5183));
  assign v_5184 = v_5185 | v_5186;
  assign v_5185 = mux_5185(v_5171);
  assign v_5186 = mux_5186(v_5187);
  assign v_5187 = ~v_5171;
  assign v_5188 = v_5189 & 1'h1;
  assign v_5189 = v_5190 & v_5191;
  assign v_5190 = ~act_5170;
  assign v_5191 = v_5192 | v_5200;
  assign v_5192 = v_5193 | v_5198;
  assign v_5193 = mux_5193(v_5194);
  assign v_5194 = v_5167 & v_5195;
  assign v_5195 = v_5196 & 1'h1;
  assign v_5196 = v_5197 | 1'h0;
  assign v_5197 = ~v_5160;
  assign v_5198 = mux_5198(v_5199);
  assign v_5199 = ~v_5194;
  assign v_5200 = ~v_5167;
  assign v_5201 = v_5202 | v_5203;
  assign v_5202 = mux_5202(v_5169);
  assign v_5203 = mux_5203(v_5188);
  assign v_5205 = v_5206 | v_5225;
  assign v_5206 = act_5207 & 1'h1;
  assign act_5207 = v_5208 | v_5214;
  assign v_5208 = v_5209 & v_5215;
  assign v_5209 = v_5210 & vout_canPeek_5220;
  assign v_5210 = ~vout_canPeek_5211;
  pebbles_core
    pebbles_core_5211
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5212),
       .in0_consume_en(vin0_consume_en_5211),
       .out_canPeek(vout_canPeek_5211),
       .out_peek(vout_peek_5211));
  assign v_5212 = v_5213 | v_5218;
  assign v_5213 = mux_5213(v_5214);
  assign v_5214 = vout_canPeek_5211 & v_5215;
  assign v_5215 = v_5216 & 1'h1;
  assign v_5216 = v_5217 | 1'h0;
  assign v_5217 = ~v_5204;
  assign v_5218 = mux_5218(v_5219);
  assign v_5219 = ~v_5214;
  pebbles_core
    pebbles_core_5220
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5221),
       .in0_consume_en(vin0_consume_en_5220),
       .out_canPeek(vout_canPeek_5220),
       .out_peek(vout_peek_5220));
  assign v_5221 = v_5222 | v_5223;
  assign v_5222 = mux_5222(v_5208);
  assign v_5223 = mux_5223(v_5224);
  assign v_5224 = ~v_5208;
  assign v_5225 = v_5226 & 1'h1;
  assign v_5226 = v_5227 & v_5228;
  assign v_5227 = ~act_5207;
  assign v_5228 = v_5229 | v_5233;
  assign v_5229 = v_5230 | v_5231;
  assign v_5230 = mux_5230(v_5164);
  assign v_5231 = mux_5231(v_5232);
  assign v_5232 = ~v_5164;
  assign v_5233 = ~v_5204;
  assign v_5234 = v_5235 | v_5236;
  assign v_5235 = mux_5235(v_5206);
  assign v_5236 = mux_5236(v_5225);
  assign v_5237 = v_5238 & 1'h1;
  assign v_5238 = v_5239 & v_5240;
  assign v_5239 = ~act_5163;
  assign v_5240 = v_5241 | v_5245;
  assign v_5241 = v_5242 | v_5243;
  assign v_5242 = mux_5242(v_5064);
  assign v_5243 = mux_5243(v_5244);
  assign v_5244 = ~v_5064;
  assign v_5245 = ~v_5160;
  assign v_5246 = v_5247 | v_5248;
  assign v_5247 = mux_5247(v_5162);
  assign v_5248 = mux_5248(v_5237);
  assign v_5249 = v_5250 & 1'h1;
  assign v_5250 = v_5251 & v_5252;
  assign v_5251 = ~act_5063;
  assign v_5252 = v_5253 | v_5257;
  assign v_5253 = v_5254 | v_5255;
  assign v_5254 = mux_5254(v_4852);
  assign v_5255 = mux_5255(v_5256);
  assign v_5256 = ~v_4852;
  assign v_5257 = ~v_5060;
  assign v_5258 = v_5259 | v_5260;
  assign v_5259 = mux_5259(v_5062);
  assign v_5260 = mux_5260(v_5249);
  assign v_5261 = v_5262 & 1'h1;
  assign v_5262 = v_5263 & v_5264;
  assign v_5263 = ~act_4851;
  assign v_5264 = v_5265 | v_5269;
  assign v_5265 = v_5266 | v_5267;
  assign v_5266 = mux_5266(v_4416);
  assign v_5267 = mux_5267(v_5268);
  assign v_5268 = ~v_4416;
  assign v_5269 = ~v_4848;
  assign v_5270 = v_5271 | v_5272;
  assign v_5271 = mux_5271(v_4850);
  assign v_5272 = mux_5272(v_5261);
  assign v_5273 = v_5274 & 1'h1;
  assign v_5274 = v_5275 & v_5276;
  assign v_5275 = ~act_4415;
  assign v_5276 = v_5277 | v_5285;
  assign v_5277 = v_5278 | v_5283;
  assign v_5278 = mux_5278(v_5279);
  assign v_5279 = v_4412 & v_5280;
  assign v_5280 = v_5281 & 1'h1;
  assign v_5281 = v_5282 | 1'h0;
  assign v_5282 = ~v_4405;
  assign v_5283 = mux_5283(v_5284);
  assign v_5284 = ~v_5279;
  assign v_5285 = ~v_4412;
  assign v_5286 = v_5287 | v_5288;
  assign v_5287 = mux_5287(v_4414);
  assign v_5288 = mux_5288(v_5273);
  assign v_5290 = v_5291 | v_6150;
  assign v_5291 = act_5292 & 1'h1;
  assign act_5292 = v_5293 | v_5715;
  assign v_5293 = v_5294 & v_5716;
  assign v_5294 = v_5295 & v_5725;
  assign v_5295 = ~v_5296;
  assign v_5297 = v_5298 | v_5709;
  assign v_5298 = act_5299 & 1'h1;
  assign act_5299 = v_5300 | v_5498;
  assign v_5300 = v_5301 & v_5499;
  assign v_5301 = v_5302 & v_5508;
  assign v_5302 = ~v_5303;
  assign v_5304 = v_5305 | v_5492;
  assign v_5305 = act_5306 & 1'h1;
  assign act_5306 = v_5307 | v_5393;
  assign v_5307 = v_5308 & v_5394;
  assign v_5308 = v_5309 & v_5403;
  assign v_5309 = ~v_5310;
  assign v_5311 = v_5312 | v_5387;
  assign v_5312 = act_5313 & 1'h1;
  assign act_5313 = v_5314 | v_5344;
  assign v_5314 = v_5315 & v_5345;
  assign v_5315 = v_5316 & v_5354;
  assign v_5316 = ~v_5317;
  assign v_5318 = v_5319 | v_5338;
  assign v_5319 = act_5320 & 1'h1;
  assign act_5320 = v_5321 | v_5327;
  assign v_5321 = v_5322 & v_5328;
  assign v_5322 = v_5323 & vout_canPeek_5333;
  assign v_5323 = ~vout_canPeek_5324;
  pebbles_core
    pebbles_core_5324
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5325),
       .in0_consume_en(vin0_consume_en_5324),
       .out_canPeek(vout_canPeek_5324),
       .out_peek(vout_peek_5324));
  assign v_5325 = v_5326 | v_5331;
  assign v_5326 = mux_5326(v_5327);
  assign v_5327 = vout_canPeek_5324 & v_5328;
  assign v_5328 = v_5329 & 1'h1;
  assign v_5329 = v_5330 | 1'h0;
  assign v_5330 = ~v_5317;
  assign v_5331 = mux_5331(v_5332);
  assign v_5332 = ~v_5327;
  pebbles_core
    pebbles_core_5333
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5334),
       .in0_consume_en(vin0_consume_en_5333),
       .out_canPeek(vout_canPeek_5333),
       .out_peek(vout_peek_5333));
  assign v_5334 = v_5335 | v_5336;
  assign v_5335 = mux_5335(v_5321);
  assign v_5336 = mux_5336(v_5337);
  assign v_5337 = ~v_5321;
  assign v_5338 = v_5339 & 1'h1;
  assign v_5339 = v_5340 & v_5341;
  assign v_5340 = ~act_5320;
  assign v_5341 = v_5342 | v_5350;
  assign v_5342 = v_5343 | v_5348;
  assign v_5343 = mux_5343(v_5344);
  assign v_5344 = v_5317 & v_5345;
  assign v_5345 = v_5346 & 1'h1;
  assign v_5346 = v_5347 | 1'h0;
  assign v_5347 = ~v_5310;
  assign v_5348 = mux_5348(v_5349);
  assign v_5349 = ~v_5344;
  assign v_5350 = ~v_5317;
  assign v_5351 = v_5352 | v_5353;
  assign v_5352 = mux_5352(v_5319);
  assign v_5353 = mux_5353(v_5338);
  assign v_5355 = v_5356 | v_5375;
  assign v_5356 = act_5357 & 1'h1;
  assign act_5357 = v_5358 | v_5364;
  assign v_5358 = v_5359 & v_5365;
  assign v_5359 = v_5360 & vout_canPeek_5370;
  assign v_5360 = ~vout_canPeek_5361;
  pebbles_core
    pebbles_core_5361
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5362),
       .in0_consume_en(vin0_consume_en_5361),
       .out_canPeek(vout_canPeek_5361),
       .out_peek(vout_peek_5361));
  assign v_5362 = v_5363 | v_5368;
  assign v_5363 = mux_5363(v_5364);
  assign v_5364 = vout_canPeek_5361 & v_5365;
  assign v_5365 = v_5366 & 1'h1;
  assign v_5366 = v_5367 | 1'h0;
  assign v_5367 = ~v_5354;
  assign v_5368 = mux_5368(v_5369);
  assign v_5369 = ~v_5364;
  pebbles_core
    pebbles_core_5370
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5371),
       .in0_consume_en(vin0_consume_en_5370),
       .out_canPeek(vout_canPeek_5370),
       .out_peek(vout_peek_5370));
  assign v_5371 = v_5372 | v_5373;
  assign v_5372 = mux_5372(v_5358);
  assign v_5373 = mux_5373(v_5374);
  assign v_5374 = ~v_5358;
  assign v_5375 = v_5376 & 1'h1;
  assign v_5376 = v_5377 & v_5378;
  assign v_5377 = ~act_5357;
  assign v_5378 = v_5379 | v_5383;
  assign v_5379 = v_5380 | v_5381;
  assign v_5380 = mux_5380(v_5314);
  assign v_5381 = mux_5381(v_5382);
  assign v_5382 = ~v_5314;
  assign v_5383 = ~v_5354;
  assign v_5384 = v_5385 | v_5386;
  assign v_5385 = mux_5385(v_5356);
  assign v_5386 = mux_5386(v_5375);
  assign v_5387 = v_5388 & 1'h1;
  assign v_5388 = v_5389 & v_5390;
  assign v_5389 = ~act_5313;
  assign v_5390 = v_5391 | v_5399;
  assign v_5391 = v_5392 | v_5397;
  assign v_5392 = mux_5392(v_5393);
  assign v_5393 = v_5310 & v_5394;
  assign v_5394 = v_5395 & 1'h1;
  assign v_5395 = v_5396 | 1'h0;
  assign v_5396 = ~v_5303;
  assign v_5397 = mux_5397(v_5398);
  assign v_5398 = ~v_5393;
  assign v_5399 = ~v_5310;
  assign v_5400 = v_5401 | v_5402;
  assign v_5401 = mux_5401(v_5312);
  assign v_5402 = mux_5402(v_5387);
  assign v_5404 = v_5405 | v_5480;
  assign v_5405 = act_5406 & 1'h1;
  assign act_5406 = v_5407 | v_5437;
  assign v_5407 = v_5408 & v_5438;
  assign v_5408 = v_5409 & v_5447;
  assign v_5409 = ~v_5410;
  assign v_5411 = v_5412 | v_5431;
  assign v_5412 = act_5413 & 1'h1;
  assign act_5413 = v_5414 | v_5420;
  assign v_5414 = v_5415 & v_5421;
  assign v_5415 = v_5416 & vout_canPeek_5426;
  assign v_5416 = ~vout_canPeek_5417;
  pebbles_core
    pebbles_core_5417
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5418),
       .in0_consume_en(vin0_consume_en_5417),
       .out_canPeek(vout_canPeek_5417),
       .out_peek(vout_peek_5417));
  assign v_5418 = v_5419 | v_5424;
  assign v_5419 = mux_5419(v_5420);
  assign v_5420 = vout_canPeek_5417 & v_5421;
  assign v_5421 = v_5422 & 1'h1;
  assign v_5422 = v_5423 | 1'h0;
  assign v_5423 = ~v_5410;
  assign v_5424 = mux_5424(v_5425);
  assign v_5425 = ~v_5420;
  pebbles_core
    pebbles_core_5426
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5427),
       .in0_consume_en(vin0_consume_en_5426),
       .out_canPeek(vout_canPeek_5426),
       .out_peek(vout_peek_5426));
  assign v_5427 = v_5428 | v_5429;
  assign v_5428 = mux_5428(v_5414);
  assign v_5429 = mux_5429(v_5430);
  assign v_5430 = ~v_5414;
  assign v_5431 = v_5432 & 1'h1;
  assign v_5432 = v_5433 & v_5434;
  assign v_5433 = ~act_5413;
  assign v_5434 = v_5435 | v_5443;
  assign v_5435 = v_5436 | v_5441;
  assign v_5436 = mux_5436(v_5437);
  assign v_5437 = v_5410 & v_5438;
  assign v_5438 = v_5439 & 1'h1;
  assign v_5439 = v_5440 | 1'h0;
  assign v_5440 = ~v_5403;
  assign v_5441 = mux_5441(v_5442);
  assign v_5442 = ~v_5437;
  assign v_5443 = ~v_5410;
  assign v_5444 = v_5445 | v_5446;
  assign v_5445 = mux_5445(v_5412);
  assign v_5446 = mux_5446(v_5431);
  assign v_5448 = v_5449 | v_5468;
  assign v_5449 = act_5450 & 1'h1;
  assign act_5450 = v_5451 | v_5457;
  assign v_5451 = v_5452 & v_5458;
  assign v_5452 = v_5453 & vout_canPeek_5463;
  assign v_5453 = ~vout_canPeek_5454;
  pebbles_core
    pebbles_core_5454
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5455),
       .in0_consume_en(vin0_consume_en_5454),
       .out_canPeek(vout_canPeek_5454),
       .out_peek(vout_peek_5454));
  assign v_5455 = v_5456 | v_5461;
  assign v_5456 = mux_5456(v_5457);
  assign v_5457 = vout_canPeek_5454 & v_5458;
  assign v_5458 = v_5459 & 1'h1;
  assign v_5459 = v_5460 | 1'h0;
  assign v_5460 = ~v_5447;
  assign v_5461 = mux_5461(v_5462);
  assign v_5462 = ~v_5457;
  pebbles_core
    pebbles_core_5463
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5464),
       .in0_consume_en(vin0_consume_en_5463),
       .out_canPeek(vout_canPeek_5463),
       .out_peek(vout_peek_5463));
  assign v_5464 = v_5465 | v_5466;
  assign v_5465 = mux_5465(v_5451);
  assign v_5466 = mux_5466(v_5467);
  assign v_5467 = ~v_5451;
  assign v_5468 = v_5469 & 1'h1;
  assign v_5469 = v_5470 & v_5471;
  assign v_5470 = ~act_5450;
  assign v_5471 = v_5472 | v_5476;
  assign v_5472 = v_5473 | v_5474;
  assign v_5473 = mux_5473(v_5407);
  assign v_5474 = mux_5474(v_5475);
  assign v_5475 = ~v_5407;
  assign v_5476 = ~v_5447;
  assign v_5477 = v_5478 | v_5479;
  assign v_5478 = mux_5478(v_5449);
  assign v_5479 = mux_5479(v_5468);
  assign v_5480 = v_5481 & 1'h1;
  assign v_5481 = v_5482 & v_5483;
  assign v_5482 = ~act_5406;
  assign v_5483 = v_5484 | v_5488;
  assign v_5484 = v_5485 | v_5486;
  assign v_5485 = mux_5485(v_5307);
  assign v_5486 = mux_5486(v_5487);
  assign v_5487 = ~v_5307;
  assign v_5488 = ~v_5403;
  assign v_5489 = v_5490 | v_5491;
  assign v_5490 = mux_5490(v_5405);
  assign v_5491 = mux_5491(v_5480);
  assign v_5492 = v_5493 & 1'h1;
  assign v_5493 = v_5494 & v_5495;
  assign v_5494 = ~act_5306;
  assign v_5495 = v_5496 | v_5504;
  assign v_5496 = v_5497 | v_5502;
  assign v_5497 = mux_5497(v_5498);
  assign v_5498 = v_5303 & v_5499;
  assign v_5499 = v_5500 & 1'h1;
  assign v_5500 = v_5501 | 1'h0;
  assign v_5501 = ~v_5296;
  assign v_5502 = mux_5502(v_5503);
  assign v_5503 = ~v_5498;
  assign v_5504 = ~v_5303;
  assign v_5505 = v_5506 | v_5507;
  assign v_5506 = mux_5506(v_5305);
  assign v_5507 = mux_5507(v_5492);
  assign v_5509 = v_5510 | v_5697;
  assign v_5510 = act_5511 & 1'h1;
  assign act_5511 = v_5512 | v_5598;
  assign v_5512 = v_5513 & v_5599;
  assign v_5513 = v_5514 & v_5608;
  assign v_5514 = ~v_5515;
  assign v_5516 = v_5517 | v_5592;
  assign v_5517 = act_5518 & 1'h1;
  assign act_5518 = v_5519 | v_5549;
  assign v_5519 = v_5520 & v_5550;
  assign v_5520 = v_5521 & v_5559;
  assign v_5521 = ~v_5522;
  assign v_5523 = v_5524 | v_5543;
  assign v_5524 = act_5525 & 1'h1;
  assign act_5525 = v_5526 | v_5532;
  assign v_5526 = v_5527 & v_5533;
  assign v_5527 = v_5528 & vout_canPeek_5538;
  assign v_5528 = ~vout_canPeek_5529;
  pebbles_core
    pebbles_core_5529
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5530),
       .in0_consume_en(vin0_consume_en_5529),
       .out_canPeek(vout_canPeek_5529),
       .out_peek(vout_peek_5529));
  assign v_5530 = v_5531 | v_5536;
  assign v_5531 = mux_5531(v_5532);
  assign v_5532 = vout_canPeek_5529 & v_5533;
  assign v_5533 = v_5534 & 1'h1;
  assign v_5534 = v_5535 | 1'h0;
  assign v_5535 = ~v_5522;
  assign v_5536 = mux_5536(v_5537);
  assign v_5537 = ~v_5532;
  pebbles_core
    pebbles_core_5538
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5539),
       .in0_consume_en(vin0_consume_en_5538),
       .out_canPeek(vout_canPeek_5538),
       .out_peek(vout_peek_5538));
  assign v_5539 = v_5540 | v_5541;
  assign v_5540 = mux_5540(v_5526);
  assign v_5541 = mux_5541(v_5542);
  assign v_5542 = ~v_5526;
  assign v_5543 = v_5544 & 1'h1;
  assign v_5544 = v_5545 & v_5546;
  assign v_5545 = ~act_5525;
  assign v_5546 = v_5547 | v_5555;
  assign v_5547 = v_5548 | v_5553;
  assign v_5548 = mux_5548(v_5549);
  assign v_5549 = v_5522 & v_5550;
  assign v_5550 = v_5551 & 1'h1;
  assign v_5551 = v_5552 | 1'h0;
  assign v_5552 = ~v_5515;
  assign v_5553 = mux_5553(v_5554);
  assign v_5554 = ~v_5549;
  assign v_5555 = ~v_5522;
  assign v_5556 = v_5557 | v_5558;
  assign v_5557 = mux_5557(v_5524);
  assign v_5558 = mux_5558(v_5543);
  assign v_5560 = v_5561 | v_5580;
  assign v_5561 = act_5562 & 1'h1;
  assign act_5562 = v_5563 | v_5569;
  assign v_5563 = v_5564 & v_5570;
  assign v_5564 = v_5565 & vout_canPeek_5575;
  assign v_5565 = ~vout_canPeek_5566;
  pebbles_core
    pebbles_core_5566
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5567),
       .in0_consume_en(vin0_consume_en_5566),
       .out_canPeek(vout_canPeek_5566),
       .out_peek(vout_peek_5566));
  assign v_5567 = v_5568 | v_5573;
  assign v_5568 = mux_5568(v_5569);
  assign v_5569 = vout_canPeek_5566 & v_5570;
  assign v_5570 = v_5571 & 1'h1;
  assign v_5571 = v_5572 | 1'h0;
  assign v_5572 = ~v_5559;
  assign v_5573 = mux_5573(v_5574);
  assign v_5574 = ~v_5569;
  pebbles_core
    pebbles_core_5575
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5576),
       .in0_consume_en(vin0_consume_en_5575),
       .out_canPeek(vout_canPeek_5575),
       .out_peek(vout_peek_5575));
  assign v_5576 = v_5577 | v_5578;
  assign v_5577 = mux_5577(v_5563);
  assign v_5578 = mux_5578(v_5579);
  assign v_5579 = ~v_5563;
  assign v_5580 = v_5581 & 1'h1;
  assign v_5581 = v_5582 & v_5583;
  assign v_5582 = ~act_5562;
  assign v_5583 = v_5584 | v_5588;
  assign v_5584 = v_5585 | v_5586;
  assign v_5585 = mux_5585(v_5519);
  assign v_5586 = mux_5586(v_5587);
  assign v_5587 = ~v_5519;
  assign v_5588 = ~v_5559;
  assign v_5589 = v_5590 | v_5591;
  assign v_5590 = mux_5590(v_5561);
  assign v_5591 = mux_5591(v_5580);
  assign v_5592 = v_5593 & 1'h1;
  assign v_5593 = v_5594 & v_5595;
  assign v_5594 = ~act_5518;
  assign v_5595 = v_5596 | v_5604;
  assign v_5596 = v_5597 | v_5602;
  assign v_5597 = mux_5597(v_5598);
  assign v_5598 = v_5515 & v_5599;
  assign v_5599 = v_5600 & 1'h1;
  assign v_5600 = v_5601 | 1'h0;
  assign v_5601 = ~v_5508;
  assign v_5602 = mux_5602(v_5603);
  assign v_5603 = ~v_5598;
  assign v_5604 = ~v_5515;
  assign v_5605 = v_5606 | v_5607;
  assign v_5606 = mux_5606(v_5517);
  assign v_5607 = mux_5607(v_5592);
  assign v_5609 = v_5610 | v_5685;
  assign v_5610 = act_5611 & 1'h1;
  assign act_5611 = v_5612 | v_5642;
  assign v_5612 = v_5613 & v_5643;
  assign v_5613 = v_5614 & v_5652;
  assign v_5614 = ~v_5615;
  assign v_5616 = v_5617 | v_5636;
  assign v_5617 = act_5618 & 1'h1;
  assign act_5618 = v_5619 | v_5625;
  assign v_5619 = v_5620 & v_5626;
  assign v_5620 = v_5621 & vout_canPeek_5631;
  assign v_5621 = ~vout_canPeek_5622;
  pebbles_core
    pebbles_core_5622
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5623),
       .in0_consume_en(vin0_consume_en_5622),
       .out_canPeek(vout_canPeek_5622),
       .out_peek(vout_peek_5622));
  assign v_5623 = v_5624 | v_5629;
  assign v_5624 = mux_5624(v_5625);
  assign v_5625 = vout_canPeek_5622 & v_5626;
  assign v_5626 = v_5627 & 1'h1;
  assign v_5627 = v_5628 | 1'h0;
  assign v_5628 = ~v_5615;
  assign v_5629 = mux_5629(v_5630);
  assign v_5630 = ~v_5625;
  pebbles_core
    pebbles_core_5631
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5632),
       .in0_consume_en(vin0_consume_en_5631),
       .out_canPeek(vout_canPeek_5631),
       .out_peek(vout_peek_5631));
  assign v_5632 = v_5633 | v_5634;
  assign v_5633 = mux_5633(v_5619);
  assign v_5634 = mux_5634(v_5635);
  assign v_5635 = ~v_5619;
  assign v_5636 = v_5637 & 1'h1;
  assign v_5637 = v_5638 & v_5639;
  assign v_5638 = ~act_5618;
  assign v_5639 = v_5640 | v_5648;
  assign v_5640 = v_5641 | v_5646;
  assign v_5641 = mux_5641(v_5642);
  assign v_5642 = v_5615 & v_5643;
  assign v_5643 = v_5644 & 1'h1;
  assign v_5644 = v_5645 | 1'h0;
  assign v_5645 = ~v_5608;
  assign v_5646 = mux_5646(v_5647);
  assign v_5647 = ~v_5642;
  assign v_5648 = ~v_5615;
  assign v_5649 = v_5650 | v_5651;
  assign v_5650 = mux_5650(v_5617);
  assign v_5651 = mux_5651(v_5636);
  assign v_5653 = v_5654 | v_5673;
  assign v_5654 = act_5655 & 1'h1;
  assign act_5655 = v_5656 | v_5662;
  assign v_5656 = v_5657 & v_5663;
  assign v_5657 = v_5658 & vout_canPeek_5668;
  assign v_5658 = ~vout_canPeek_5659;
  pebbles_core
    pebbles_core_5659
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5660),
       .in0_consume_en(vin0_consume_en_5659),
       .out_canPeek(vout_canPeek_5659),
       .out_peek(vout_peek_5659));
  assign v_5660 = v_5661 | v_5666;
  assign v_5661 = mux_5661(v_5662);
  assign v_5662 = vout_canPeek_5659 & v_5663;
  assign v_5663 = v_5664 & 1'h1;
  assign v_5664 = v_5665 | 1'h0;
  assign v_5665 = ~v_5652;
  assign v_5666 = mux_5666(v_5667);
  assign v_5667 = ~v_5662;
  pebbles_core
    pebbles_core_5668
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5669),
       .in0_consume_en(vin0_consume_en_5668),
       .out_canPeek(vout_canPeek_5668),
       .out_peek(vout_peek_5668));
  assign v_5669 = v_5670 | v_5671;
  assign v_5670 = mux_5670(v_5656);
  assign v_5671 = mux_5671(v_5672);
  assign v_5672 = ~v_5656;
  assign v_5673 = v_5674 & 1'h1;
  assign v_5674 = v_5675 & v_5676;
  assign v_5675 = ~act_5655;
  assign v_5676 = v_5677 | v_5681;
  assign v_5677 = v_5678 | v_5679;
  assign v_5678 = mux_5678(v_5612);
  assign v_5679 = mux_5679(v_5680);
  assign v_5680 = ~v_5612;
  assign v_5681 = ~v_5652;
  assign v_5682 = v_5683 | v_5684;
  assign v_5683 = mux_5683(v_5654);
  assign v_5684 = mux_5684(v_5673);
  assign v_5685 = v_5686 & 1'h1;
  assign v_5686 = v_5687 & v_5688;
  assign v_5687 = ~act_5611;
  assign v_5688 = v_5689 | v_5693;
  assign v_5689 = v_5690 | v_5691;
  assign v_5690 = mux_5690(v_5512);
  assign v_5691 = mux_5691(v_5692);
  assign v_5692 = ~v_5512;
  assign v_5693 = ~v_5608;
  assign v_5694 = v_5695 | v_5696;
  assign v_5695 = mux_5695(v_5610);
  assign v_5696 = mux_5696(v_5685);
  assign v_5697 = v_5698 & 1'h1;
  assign v_5698 = v_5699 & v_5700;
  assign v_5699 = ~act_5511;
  assign v_5700 = v_5701 | v_5705;
  assign v_5701 = v_5702 | v_5703;
  assign v_5702 = mux_5702(v_5300);
  assign v_5703 = mux_5703(v_5704);
  assign v_5704 = ~v_5300;
  assign v_5705 = ~v_5508;
  assign v_5706 = v_5707 | v_5708;
  assign v_5707 = mux_5707(v_5510);
  assign v_5708 = mux_5708(v_5697);
  assign v_5709 = v_5710 & 1'h1;
  assign v_5710 = v_5711 & v_5712;
  assign v_5711 = ~act_5299;
  assign v_5712 = v_5713 | v_5721;
  assign v_5713 = v_5714 | v_5719;
  assign v_5714 = mux_5714(v_5715);
  assign v_5715 = v_5296 & v_5716;
  assign v_5716 = v_5717 & 1'h1;
  assign v_5717 = v_5718 | 1'h0;
  assign v_5718 = ~v_5289;
  assign v_5719 = mux_5719(v_5720);
  assign v_5720 = ~v_5715;
  assign v_5721 = ~v_5296;
  assign v_5722 = v_5723 | v_5724;
  assign v_5723 = mux_5723(v_5298);
  assign v_5724 = mux_5724(v_5709);
  assign v_5726 = v_5727 | v_6138;
  assign v_5727 = act_5728 & 1'h1;
  assign act_5728 = v_5729 | v_5927;
  assign v_5729 = v_5730 & v_5928;
  assign v_5730 = v_5731 & v_5937;
  assign v_5731 = ~v_5732;
  assign v_5733 = v_5734 | v_5921;
  assign v_5734 = act_5735 & 1'h1;
  assign act_5735 = v_5736 | v_5822;
  assign v_5736 = v_5737 & v_5823;
  assign v_5737 = v_5738 & v_5832;
  assign v_5738 = ~v_5739;
  assign v_5740 = v_5741 | v_5816;
  assign v_5741 = act_5742 & 1'h1;
  assign act_5742 = v_5743 | v_5773;
  assign v_5743 = v_5744 & v_5774;
  assign v_5744 = v_5745 & v_5783;
  assign v_5745 = ~v_5746;
  assign v_5747 = v_5748 | v_5767;
  assign v_5748 = act_5749 & 1'h1;
  assign act_5749 = v_5750 | v_5756;
  assign v_5750 = v_5751 & v_5757;
  assign v_5751 = v_5752 & vout_canPeek_5762;
  assign v_5752 = ~vout_canPeek_5753;
  pebbles_core
    pebbles_core_5753
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5754),
       .in0_consume_en(vin0_consume_en_5753),
       .out_canPeek(vout_canPeek_5753),
       .out_peek(vout_peek_5753));
  assign v_5754 = v_5755 | v_5760;
  assign v_5755 = mux_5755(v_5756);
  assign v_5756 = vout_canPeek_5753 & v_5757;
  assign v_5757 = v_5758 & 1'h1;
  assign v_5758 = v_5759 | 1'h0;
  assign v_5759 = ~v_5746;
  assign v_5760 = mux_5760(v_5761);
  assign v_5761 = ~v_5756;
  pebbles_core
    pebbles_core_5762
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5763),
       .in0_consume_en(vin0_consume_en_5762),
       .out_canPeek(vout_canPeek_5762),
       .out_peek(vout_peek_5762));
  assign v_5763 = v_5764 | v_5765;
  assign v_5764 = mux_5764(v_5750);
  assign v_5765 = mux_5765(v_5766);
  assign v_5766 = ~v_5750;
  assign v_5767 = v_5768 & 1'h1;
  assign v_5768 = v_5769 & v_5770;
  assign v_5769 = ~act_5749;
  assign v_5770 = v_5771 | v_5779;
  assign v_5771 = v_5772 | v_5777;
  assign v_5772 = mux_5772(v_5773);
  assign v_5773 = v_5746 & v_5774;
  assign v_5774 = v_5775 & 1'h1;
  assign v_5775 = v_5776 | 1'h0;
  assign v_5776 = ~v_5739;
  assign v_5777 = mux_5777(v_5778);
  assign v_5778 = ~v_5773;
  assign v_5779 = ~v_5746;
  assign v_5780 = v_5781 | v_5782;
  assign v_5781 = mux_5781(v_5748);
  assign v_5782 = mux_5782(v_5767);
  assign v_5784 = v_5785 | v_5804;
  assign v_5785 = act_5786 & 1'h1;
  assign act_5786 = v_5787 | v_5793;
  assign v_5787 = v_5788 & v_5794;
  assign v_5788 = v_5789 & vout_canPeek_5799;
  assign v_5789 = ~vout_canPeek_5790;
  pebbles_core
    pebbles_core_5790
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5791),
       .in0_consume_en(vin0_consume_en_5790),
       .out_canPeek(vout_canPeek_5790),
       .out_peek(vout_peek_5790));
  assign v_5791 = v_5792 | v_5797;
  assign v_5792 = mux_5792(v_5793);
  assign v_5793 = vout_canPeek_5790 & v_5794;
  assign v_5794 = v_5795 & 1'h1;
  assign v_5795 = v_5796 | 1'h0;
  assign v_5796 = ~v_5783;
  assign v_5797 = mux_5797(v_5798);
  assign v_5798 = ~v_5793;
  pebbles_core
    pebbles_core_5799
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5800),
       .in0_consume_en(vin0_consume_en_5799),
       .out_canPeek(vout_canPeek_5799),
       .out_peek(vout_peek_5799));
  assign v_5800 = v_5801 | v_5802;
  assign v_5801 = mux_5801(v_5787);
  assign v_5802 = mux_5802(v_5803);
  assign v_5803 = ~v_5787;
  assign v_5804 = v_5805 & 1'h1;
  assign v_5805 = v_5806 & v_5807;
  assign v_5806 = ~act_5786;
  assign v_5807 = v_5808 | v_5812;
  assign v_5808 = v_5809 | v_5810;
  assign v_5809 = mux_5809(v_5743);
  assign v_5810 = mux_5810(v_5811);
  assign v_5811 = ~v_5743;
  assign v_5812 = ~v_5783;
  assign v_5813 = v_5814 | v_5815;
  assign v_5814 = mux_5814(v_5785);
  assign v_5815 = mux_5815(v_5804);
  assign v_5816 = v_5817 & 1'h1;
  assign v_5817 = v_5818 & v_5819;
  assign v_5818 = ~act_5742;
  assign v_5819 = v_5820 | v_5828;
  assign v_5820 = v_5821 | v_5826;
  assign v_5821 = mux_5821(v_5822);
  assign v_5822 = v_5739 & v_5823;
  assign v_5823 = v_5824 & 1'h1;
  assign v_5824 = v_5825 | 1'h0;
  assign v_5825 = ~v_5732;
  assign v_5826 = mux_5826(v_5827);
  assign v_5827 = ~v_5822;
  assign v_5828 = ~v_5739;
  assign v_5829 = v_5830 | v_5831;
  assign v_5830 = mux_5830(v_5741);
  assign v_5831 = mux_5831(v_5816);
  assign v_5833 = v_5834 | v_5909;
  assign v_5834 = act_5835 & 1'h1;
  assign act_5835 = v_5836 | v_5866;
  assign v_5836 = v_5837 & v_5867;
  assign v_5837 = v_5838 & v_5876;
  assign v_5838 = ~v_5839;
  assign v_5840 = v_5841 | v_5860;
  assign v_5841 = act_5842 & 1'h1;
  assign act_5842 = v_5843 | v_5849;
  assign v_5843 = v_5844 & v_5850;
  assign v_5844 = v_5845 & vout_canPeek_5855;
  assign v_5845 = ~vout_canPeek_5846;
  pebbles_core
    pebbles_core_5846
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5847),
       .in0_consume_en(vin0_consume_en_5846),
       .out_canPeek(vout_canPeek_5846),
       .out_peek(vout_peek_5846));
  assign v_5847 = v_5848 | v_5853;
  assign v_5848 = mux_5848(v_5849);
  assign v_5849 = vout_canPeek_5846 & v_5850;
  assign v_5850 = v_5851 & 1'h1;
  assign v_5851 = v_5852 | 1'h0;
  assign v_5852 = ~v_5839;
  assign v_5853 = mux_5853(v_5854);
  assign v_5854 = ~v_5849;
  pebbles_core
    pebbles_core_5855
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5856),
       .in0_consume_en(vin0_consume_en_5855),
       .out_canPeek(vout_canPeek_5855),
       .out_peek(vout_peek_5855));
  assign v_5856 = v_5857 | v_5858;
  assign v_5857 = mux_5857(v_5843);
  assign v_5858 = mux_5858(v_5859);
  assign v_5859 = ~v_5843;
  assign v_5860 = v_5861 & 1'h1;
  assign v_5861 = v_5862 & v_5863;
  assign v_5862 = ~act_5842;
  assign v_5863 = v_5864 | v_5872;
  assign v_5864 = v_5865 | v_5870;
  assign v_5865 = mux_5865(v_5866);
  assign v_5866 = v_5839 & v_5867;
  assign v_5867 = v_5868 & 1'h1;
  assign v_5868 = v_5869 | 1'h0;
  assign v_5869 = ~v_5832;
  assign v_5870 = mux_5870(v_5871);
  assign v_5871 = ~v_5866;
  assign v_5872 = ~v_5839;
  assign v_5873 = v_5874 | v_5875;
  assign v_5874 = mux_5874(v_5841);
  assign v_5875 = mux_5875(v_5860);
  assign v_5877 = v_5878 | v_5897;
  assign v_5878 = act_5879 & 1'h1;
  assign act_5879 = v_5880 | v_5886;
  assign v_5880 = v_5881 & v_5887;
  assign v_5881 = v_5882 & vout_canPeek_5892;
  assign v_5882 = ~vout_canPeek_5883;
  pebbles_core
    pebbles_core_5883
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5884),
       .in0_consume_en(vin0_consume_en_5883),
       .out_canPeek(vout_canPeek_5883),
       .out_peek(vout_peek_5883));
  assign v_5884 = v_5885 | v_5890;
  assign v_5885 = mux_5885(v_5886);
  assign v_5886 = vout_canPeek_5883 & v_5887;
  assign v_5887 = v_5888 & 1'h1;
  assign v_5888 = v_5889 | 1'h0;
  assign v_5889 = ~v_5876;
  assign v_5890 = mux_5890(v_5891);
  assign v_5891 = ~v_5886;
  pebbles_core
    pebbles_core_5892
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5893),
       .in0_consume_en(vin0_consume_en_5892),
       .out_canPeek(vout_canPeek_5892),
       .out_peek(vout_peek_5892));
  assign v_5893 = v_5894 | v_5895;
  assign v_5894 = mux_5894(v_5880);
  assign v_5895 = mux_5895(v_5896);
  assign v_5896 = ~v_5880;
  assign v_5897 = v_5898 & 1'h1;
  assign v_5898 = v_5899 & v_5900;
  assign v_5899 = ~act_5879;
  assign v_5900 = v_5901 | v_5905;
  assign v_5901 = v_5902 | v_5903;
  assign v_5902 = mux_5902(v_5836);
  assign v_5903 = mux_5903(v_5904);
  assign v_5904 = ~v_5836;
  assign v_5905 = ~v_5876;
  assign v_5906 = v_5907 | v_5908;
  assign v_5907 = mux_5907(v_5878);
  assign v_5908 = mux_5908(v_5897);
  assign v_5909 = v_5910 & 1'h1;
  assign v_5910 = v_5911 & v_5912;
  assign v_5911 = ~act_5835;
  assign v_5912 = v_5913 | v_5917;
  assign v_5913 = v_5914 | v_5915;
  assign v_5914 = mux_5914(v_5736);
  assign v_5915 = mux_5915(v_5916);
  assign v_5916 = ~v_5736;
  assign v_5917 = ~v_5832;
  assign v_5918 = v_5919 | v_5920;
  assign v_5919 = mux_5919(v_5834);
  assign v_5920 = mux_5920(v_5909);
  assign v_5921 = v_5922 & 1'h1;
  assign v_5922 = v_5923 & v_5924;
  assign v_5923 = ~act_5735;
  assign v_5924 = v_5925 | v_5933;
  assign v_5925 = v_5926 | v_5931;
  assign v_5926 = mux_5926(v_5927);
  assign v_5927 = v_5732 & v_5928;
  assign v_5928 = v_5929 & 1'h1;
  assign v_5929 = v_5930 | 1'h0;
  assign v_5930 = ~v_5725;
  assign v_5931 = mux_5931(v_5932);
  assign v_5932 = ~v_5927;
  assign v_5933 = ~v_5732;
  assign v_5934 = v_5935 | v_5936;
  assign v_5935 = mux_5935(v_5734);
  assign v_5936 = mux_5936(v_5921);
  assign v_5938 = v_5939 | v_6126;
  assign v_5939 = act_5940 & 1'h1;
  assign act_5940 = v_5941 | v_6027;
  assign v_5941 = v_5942 & v_6028;
  assign v_5942 = v_5943 & v_6037;
  assign v_5943 = ~v_5944;
  assign v_5945 = v_5946 | v_6021;
  assign v_5946 = act_5947 & 1'h1;
  assign act_5947 = v_5948 | v_5978;
  assign v_5948 = v_5949 & v_5979;
  assign v_5949 = v_5950 & v_5988;
  assign v_5950 = ~v_5951;
  assign v_5952 = v_5953 | v_5972;
  assign v_5953 = act_5954 & 1'h1;
  assign act_5954 = v_5955 | v_5961;
  assign v_5955 = v_5956 & v_5962;
  assign v_5956 = v_5957 & vout_canPeek_5967;
  assign v_5957 = ~vout_canPeek_5958;
  pebbles_core
    pebbles_core_5958
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5959),
       .in0_consume_en(vin0_consume_en_5958),
       .out_canPeek(vout_canPeek_5958),
       .out_peek(vout_peek_5958));
  assign v_5959 = v_5960 | v_5965;
  assign v_5960 = mux_5960(v_5961);
  assign v_5961 = vout_canPeek_5958 & v_5962;
  assign v_5962 = v_5963 & 1'h1;
  assign v_5963 = v_5964 | 1'h0;
  assign v_5964 = ~v_5951;
  assign v_5965 = mux_5965(v_5966);
  assign v_5966 = ~v_5961;
  pebbles_core
    pebbles_core_5967
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5968),
       .in0_consume_en(vin0_consume_en_5967),
       .out_canPeek(vout_canPeek_5967),
       .out_peek(vout_peek_5967));
  assign v_5968 = v_5969 | v_5970;
  assign v_5969 = mux_5969(v_5955);
  assign v_5970 = mux_5970(v_5971);
  assign v_5971 = ~v_5955;
  assign v_5972 = v_5973 & 1'h1;
  assign v_5973 = v_5974 & v_5975;
  assign v_5974 = ~act_5954;
  assign v_5975 = v_5976 | v_5984;
  assign v_5976 = v_5977 | v_5982;
  assign v_5977 = mux_5977(v_5978);
  assign v_5978 = v_5951 & v_5979;
  assign v_5979 = v_5980 & 1'h1;
  assign v_5980 = v_5981 | 1'h0;
  assign v_5981 = ~v_5944;
  assign v_5982 = mux_5982(v_5983);
  assign v_5983 = ~v_5978;
  assign v_5984 = ~v_5951;
  assign v_5985 = v_5986 | v_5987;
  assign v_5986 = mux_5986(v_5953);
  assign v_5987 = mux_5987(v_5972);
  assign v_5989 = v_5990 | v_6009;
  assign v_5990 = act_5991 & 1'h1;
  assign act_5991 = v_5992 | v_5998;
  assign v_5992 = v_5993 & v_5999;
  assign v_5993 = v_5994 & vout_canPeek_6004;
  assign v_5994 = ~vout_canPeek_5995;
  pebbles_core
    pebbles_core_5995
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_5996),
       .in0_consume_en(vin0_consume_en_5995),
       .out_canPeek(vout_canPeek_5995),
       .out_peek(vout_peek_5995));
  assign v_5996 = v_5997 | v_6002;
  assign v_5997 = mux_5997(v_5998);
  assign v_5998 = vout_canPeek_5995 & v_5999;
  assign v_5999 = v_6000 & 1'h1;
  assign v_6000 = v_6001 | 1'h0;
  assign v_6001 = ~v_5988;
  assign v_6002 = mux_6002(v_6003);
  assign v_6003 = ~v_5998;
  pebbles_core
    pebbles_core_6004
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6005),
       .in0_consume_en(vin0_consume_en_6004),
       .out_canPeek(vout_canPeek_6004),
       .out_peek(vout_peek_6004));
  assign v_6005 = v_6006 | v_6007;
  assign v_6006 = mux_6006(v_5992);
  assign v_6007 = mux_6007(v_6008);
  assign v_6008 = ~v_5992;
  assign v_6009 = v_6010 & 1'h1;
  assign v_6010 = v_6011 & v_6012;
  assign v_6011 = ~act_5991;
  assign v_6012 = v_6013 | v_6017;
  assign v_6013 = v_6014 | v_6015;
  assign v_6014 = mux_6014(v_5948);
  assign v_6015 = mux_6015(v_6016);
  assign v_6016 = ~v_5948;
  assign v_6017 = ~v_5988;
  assign v_6018 = v_6019 | v_6020;
  assign v_6019 = mux_6019(v_5990);
  assign v_6020 = mux_6020(v_6009);
  assign v_6021 = v_6022 & 1'h1;
  assign v_6022 = v_6023 & v_6024;
  assign v_6023 = ~act_5947;
  assign v_6024 = v_6025 | v_6033;
  assign v_6025 = v_6026 | v_6031;
  assign v_6026 = mux_6026(v_6027);
  assign v_6027 = v_5944 & v_6028;
  assign v_6028 = v_6029 & 1'h1;
  assign v_6029 = v_6030 | 1'h0;
  assign v_6030 = ~v_5937;
  assign v_6031 = mux_6031(v_6032);
  assign v_6032 = ~v_6027;
  assign v_6033 = ~v_5944;
  assign v_6034 = v_6035 | v_6036;
  assign v_6035 = mux_6035(v_5946);
  assign v_6036 = mux_6036(v_6021);
  assign v_6038 = v_6039 | v_6114;
  assign v_6039 = act_6040 & 1'h1;
  assign act_6040 = v_6041 | v_6071;
  assign v_6041 = v_6042 & v_6072;
  assign v_6042 = v_6043 & v_6081;
  assign v_6043 = ~v_6044;
  assign v_6045 = v_6046 | v_6065;
  assign v_6046 = act_6047 & 1'h1;
  assign act_6047 = v_6048 | v_6054;
  assign v_6048 = v_6049 & v_6055;
  assign v_6049 = v_6050 & vout_canPeek_6060;
  assign v_6050 = ~vout_canPeek_6051;
  pebbles_core
    pebbles_core_6051
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6052),
       .in0_consume_en(vin0_consume_en_6051),
       .out_canPeek(vout_canPeek_6051),
       .out_peek(vout_peek_6051));
  assign v_6052 = v_6053 | v_6058;
  assign v_6053 = mux_6053(v_6054);
  assign v_6054 = vout_canPeek_6051 & v_6055;
  assign v_6055 = v_6056 & 1'h1;
  assign v_6056 = v_6057 | 1'h0;
  assign v_6057 = ~v_6044;
  assign v_6058 = mux_6058(v_6059);
  assign v_6059 = ~v_6054;
  pebbles_core
    pebbles_core_6060
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6061),
       .in0_consume_en(vin0_consume_en_6060),
       .out_canPeek(vout_canPeek_6060),
       .out_peek(vout_peek_6060));
  assign v_6061 = v_6062 | v_6063;
  assign v_6062 = mux_6062(v_6048);
  assign v_6063 = mux_6063(v_6064);
  assign v_6064 = ~v_6048;
  assign v_6065 = v_6066 & 1'h1;
  assign v_6066 = v_6067 & v_6068;
  assign v_6067 = ~act_6047;
  assign v_6068 = v_6069 | v_6077;
  assign v_6069 = v_6070 | v_6075;
  assign v_6070 = mux_6070(v_6071);
  assign v_6071 = v_6044 & v_6072;
  assign v_6072 = v_6073 & 1'h1;
  assign v_6073 = v_6074 | 1'h0;
  assign v_6074 = ~v_6037;
  assign v_6075 = mux_6075(v_6076);
  assign v_6076 = ~v_6071;
  assign v_6077 = ~v_6044;
  assign v_6078 = v_6079 | v_6080;
  assign v_6079 = mux_6079(v_6046);
  assign v_6080 = mux_6080(v_6065);
  assign v_6082 = v_6083 | v_6102;
  assign v_6083 = act_6084 & 1'h1;
  assign act_6084 = v_6085 | v_6091;
  assign v_6085 = v_6086 & v_6092;
  assign v_6086 = v_6087 & vout_canPeek_6097;
  assign v_6087 = ~vout_canPeek_6088;
  pebbles_core
    pebbles_core_6088
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6089),
       .in0_consume_en(vin0_consume_en_6088),
       .out_canPeek(vout_canPeek_6088),
       .out_peek(vout_peek_6088));
  assign v_6089 = v_6090 | v_6095;
  assign v_6090 = mux_6090(v_6091);
  assign v_6091 = vout_canPeek_6088 & v_6092;
  assign v_6092 = v_6093 & 1'h1;
  assign v_6093 = v_6094 | 1'h0;
  assign v_6094 = ~v_6081;
  assign v_6095 = mux_6095(v_6096);
  assign v_6096 = ~v_6091;
  pebbles_core
    pebbles_core_6097
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6098),
       .in0_consume_en(vin0_consume_en_6097),
       .out_canPeek(vout_canPeek_6097),
       .out_peek(vout_peek_6097));
  assign v_6098 = v_6099 | v_6100;
  assign v_6099 = mux_6099(v_6085);
  assign v_6100 = mux_6100(v_6101);
  assign v_6101 = ~v_6085;
  assign v_6102 = v_6103 & 1'h1;
  assign v_6103 = v_6104 & v_6105;
  assign v_6104 = ~act_6084;
  assign v_6105 = v_6106 | v_6110;
  assign v_6106 = v_6107 | v_6108;
  assign v_6107 = mux_6107(v_6041);
  assign v_6108 = mux_6108(v_6109);
  assign v_6109 = ~v_6041;
  assign v_6110 = ~v_6081;
  assign v_6111 = v_6112 | v_6113;
  assign v_6112 = mux_6112(v_6083);
  assign v_6113 = mux_6113(v_6102);
  assign v_6114 = v_6115 & 1'h1;
  assign v_6115 = v_6116 & v_6117;
  assign v_6116 = ~act_6040;
  assign v_6117 = v_6118 | v_6122;
  assign v_6118 = v_6119 | v_6120;
  assign v_6119 = mux_6119(v_5941);
  assign v_6120 = mux_6120(v_6121);
  assign v_6121 = ~v_5941;
  assign v_6122 = ~v_6037;
  assign v_6123 = v_6124 | v_6125;
  assign v_6124 = mux_6124(v_6039);
  assign v_6125 = mux_6125(v_6114);
  assign v_6126 = v_6127 & 1'h1;
  assign v_6127 = v_6128 & v_6129;
  assign v_6128 = ~act_5940;
  assign v_6129 = v_6130 | v_6134;
  assign v_6130 = v_6131 | v_6132;
  assign v_6131 = mux_6131(v_5729);
  assign v_6132 = mux_6132(v_6133);
  assign v_6133 = ~v_5729;
  assign v_6134 = ~v_5937;
  assign v_6135 = v_6136 | v_6137;
  assign v_6136 = mux_6136(v_5939);
  assign v_6137 = mux_6137(v_6126);
  assign v_6138 = v_6139 & 1'h1;
  assign v_6139 = v_6140 & v_6141;
  assign v_6140 = ~act_5728;
  assign v_6141 = v_6142 | v_6146;
  assign v_6142 = v_6143 | v_6144;
  assign v_6143 = mux_6143(v_5293);
  assign v_6144 = mux_6144(v_6145);
  assign v_6145 = ~v_5293;
  assign v_6146 = ~v_5725;
  assign v_6147 = v_6148 | v_6149;
  assign v_6148 = mux_6148(v_5727);
  assign v_6149 = mux_6149(v_6138);
  assign v_6150 = v_6151 & 1'h1;
  assign v_6151 = v_6152 & v_6153;
  assign v_6152 = ~act_5292;
  assign v_6153 = v_6154 | v_6158;
  assign v_6154 = v_6155 | v_6156;
  assign v_6155 = mux_6155(v_4409);
  assign v_6156 = mux_6156(v_6157);
  assign v_6157 = ~v_4409;
  assign v_6158 = ~v_5289;
  assign v_6159 = v_6160 | v_6161;
  assign v_6160 = mux_6160(v_5291);
  assign v_6161 = mux_6161(v_6150);
  assign v_6162 = v_6163 & 1'h1;
  assign v_6163 = v_6164 & v_6165;
  assign v_6164 = ~act_4408;
  assign v_6165 = v_6166 | v_6174;
  assign v_6166 = v_6167 | v_6172;
  assign v_6167 = mux_6167(v_6168);
  assign v_6168 = v_4405 & v_6169;
  assign v_6169 = v_6170 & 1'h1;
  assign v_6170 = v_6171 | 1'h0;
  assign v_6171 = ~v_4398;
  assign v_6172 = mux_6172(v_6173);
  assign v_6173 = ~v_6168;
  assign v_6174 = ~v_4405;
  assign v_6175 = v_6176 | v_6177;
  assign v_6176 = mux_6176(v_4407);
  assign v_6177 = mux_6177(v_6162);
  assign v_6179 = v_6180 | v_7935;
  assign v_6180 = act_6181 & 1'h1;
  assign act_6181 = v_6182 | v_7052;
  assign v_6182 = v_6183 & v_7053;
  assign v_6183 = v_6184 & v_7062;
  assign v_6184 = ~v_6185;
  assign v_6186 = v_6187 | v_7046;
  assign v_6187 = act_6188 & 1'h1;
  assign act_6188 = v_6189 | v_6611;
  assign v_6189 = v_6190 & v_6612;
  assign v_6190 = v_6191 & v_6621;
  assign v_6191 = ~v_6192;
  assign v_6193 = v_6194 | v_6605;
  assign v_6194 = act_6195 & 1'h1;
  assign act_6195 = v_6196 | v_6394;
  assign v_6196 = v_6197 & v_6395;
  assign v_6197 = v_6198 & v_6404;
  assign v_6198 = ~v_6199;
  assign v_6200 = v_6201 | v_6388;
  assign v_6201 = act_6202 & 1'h1;
  assign act_6202 = v_6203 | v_6289;
  assign v_6203 = v_6204 & v_6290;
  assign v_6204 = v_6205 & v_6299;
  assign v_6205 = ~v_6206;
  assign v_6207 = v_6208 | v_6283;
  assign v_6208 = act_6209 & 1'h1;
  assign act_6209 = v_6210 | v_6240;
  assign v_6210 = v_6211 & v_6241;
  assign v_6211 = v_6212 & v_6250;
  assign v_6212 = ~v_6213;
  assign v_6214 = v_6215 | v_6234;
  assign v_6215 = act_6216 & 1'h1;
  assign act_6216 = v_6217 | v_6223;
  assign v_6217 = v_6218 & v_6224;
  assign v_6218 = v_6219 & vout_canPeek_6229;
  assign v_6219 = ~vout_canPeek_6220;
  pebbles_core
    pebbles_core_6220
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6221),
       .in0_consume_en(vin0_consume_en_6220),
       .out_canPeek(vout_canPeek_6220),
       .out_peek(vout_peek_6220));
  assign v_6221 = v_6222 | v_6227;
  assign v_6222 = mux_6222(v_6223);
  assign v_6223 = vout_canPeek_6220 & v_6224;
  assign v_6224 = v_6225 & 1'h1;
  assign v_6225 = v_6226 | 1'h0;
  assign v_6226 = ~v_6213;
  assign v_6227 = mux_6227(v_6228);
  assign v_6228 = ~v_6223;
  pebbles_core
    pebbles_core_6229
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6230),
       .in0_consume_en(vin0_consume_en_6229),
       .out_canPeek(vout_canPeek_6229),
       .out_peek(vout_peek_6229));
  assign v_6230 = v_6231 | v_6232;
  assign v_6231 = mux_6231(v_6217);
  assign v_6232 = mux_6232(v_6233);
  assign v_6233 = ~v_6217;
  assign v_6234 = v_6235 & 1'h1;
  assign v_6235 = v_6236 & v_6237;
  assign v_6236 = ~act_6216;
  assign v_6237 = v_6238 | v_6246;
  assign v_6238 = v_6239 | v_6244;
  assign v_6239 = mux_6239(v_6240);
  assign v_6240 = v_6213 & v_6241;
  assign v_6241 = v_6242 & 1'h1;
  assign v_6242 = v_6243 | 1'h0;
  assign v_6243 = ~v_6206;
  assign v_6244 = mux_6244(v_6245);
  assign v_6245 = ~v_6240;
  assign v_6246 = ~v_6213;
  assign v_6247 = v_6248 | v_6249;
  assign v_6248 = mux_6248(v_6215);
  assign v_6249 = mux_6249(v_6234);
  assign v_6251 = v_6252 | v_6271;
  assign v_6252 = act_6253 & 1'h1;
  assign act_6253 = v_6254 | v_6260;
  assign v_6254 = v_6255 & v_6261;
  assign v_6255 = v_6256 & vout_canPeek_6266;
  assign v_6256 = ~vout_canPeek_6257;
  pebbles_core
    pebbles_core_6257
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6258),
       .in0_consume_en(vin0_consume_en_6257),
       .out_canPeek(vout_canPeek_6257),
       .out_peek(vout_peek_6257));
  assign v_6258 = v_6259 | v_6264;
  assign v_6259 = mux_6259(v_6260);
  assign v_6260 = vout_canPeek_6257 & v_6261;
  assign v_6261 = v_6262 & 1'h1;
  assign v_6262 = v_6263 | 1'h0;
  assign v_6263 = ~v_6250;
  assign v_6264 = mux_6264(v_6265);
  assign v_6265 = ~v_6260;
  pebbles_core
    pebbles_core_6266
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6267),
       .in0_consume_en(vin0_consume_en_6266),
       .out_canPeek(vout_canPeek_6266),
       .out_peek(vout_peek_6266));
  assign v_6267 = v_6268 | v_6269;
  assign v_6268 = mux_6268(v_6254);
  assign v_6269 = mux_6269(v_6270);
  assign v_6270 = ~v_6254;
  assign v_6271 = v_6272 & 1'h1;
  assign v_6272 = v_6273 & v_6274;
  assign v_6273 = ~act_6253;
  assign v_6274 = v_6275 | v_6279;
  assign v_6275 = v_6276 | v_6277;
  assign v_6276 = mux_6276(v_6210);
  assign v_6277 = mux_6277(v_6278);
  assign v_6278 = ~v_6210;
  assign v_6279 = ~v_6250;
  assign v_6280 = v_6281 | v_6282;
  assign v_6281 = mux_6281(v_6252);
  assign v_6282 = mux_6282(v_6271);
  assign v_6283 = v_6284 & 1'h1;
  assign v_6284 = v_6285 & v_6286;
  assign v_6285 = ~act_6209;
  assign v_6286 = v_6287 | v_6295;
  assign v_6287 = v_6288 | v_6293;
  assign v_6288 = mux_6288(v_6289);
  assign v_6289 = v_6206 & v_6290;
  assign v_6290 = v_6291 & 1'h1;
  assign v_6291 = v_6292 | 1'h0;
  assign v_6292 = ~v_6199;
  assign v_6293 = mux_6293(v_6294);
  assign v_6294 = ~v_6289;
  assign v_6295 = ~v_6206;
  assign v_6296 = v_6297 | v_6298;
  assign v_6297 = mux_6297(v_6208);
  assign v_6298 = mux_6298(v_6283);
  assign v_6300 = v_6301 | v_6376;
  assign v_6301 = act_6302 & 1'h1;
  assign act_6302 = v_6303 | v_6333;
  assign v_6303 = v_6304 & v_6334;
  assign v_6304 = v_6305 & v_6343;
  assign v_6305 = ~v_6306;
  assign v_6307 = v_6308 | v_6327;
  assign v_6308 = act_6309 & 1'h1;
  assign act_6309 = v_6310 | v_6316;
  assign v_6310 = v_6311 & v_6317;
  assign v_6311 = v_6312 & vout_canPeek_6322;
  assign v_6312 = ~vout_canPeek_6313;
  pebbles_core
    pebbles_core_6313
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6314),
       .in0_consume_en(vin0_consume_en_6313),
       .out_canPeek(vout_canPeek_6313),
       .out_peek(vout_peek_6313));
  assign v_6314 = v_6315 | v_6320;
  assign v_6315 = mux_6315(v_6316);
  assign v_6316 = vout_canPeek_6313 & v_6317;
  assign v_6317 = v_6318 & 1'h1;
  assign v_6318 = v_6319 | 1'h0;
  assign v_6319 = ~v_6306;
  assign v_6320 = mux_6320(v_6321);
  assign v_6321 = ~v_6316;
  pebbles_core
    pebbles_core_6322
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6323),
       .in0_consume_en(vin0_consume_en_6322),
       .out_canPeek(vout_canPeek_6322),
       .out_peek(vout_peek_6322));
  assign v_6323 = v_6324 | v_6325;
  assign v_6324 = mux_6324(v_6310);
  assign v_6325 = mux_6325(v_6326);
  assign v_6326 = ~v_6310;
  assign v_6327 = v_6328 & 1'h1;
  assign v_6328 = v_6329 & v_6330;
  assign v_6329 = ~act_6309;
  assign v_6330 = v_6331 | v_6339;
  assign v_6331 = v_6332 | v_6337;
  assign v_6332 = mux_6332(v_6333);
  assign v_6333 = v_6306 & v_6334;
  assign v_6334 = v_6335 & 1'h1;
  assign v_6335 = v_6336 | 1'h0;
  assign v_6336 = ~v_6299;
  assign v_6337 = mux_6337(v_6338);
  assign v_6338 = ~v_6333;
  assign v_6339 = ~v_6306;
  assign v_6340 = v_6341 | v_6342;
  assign v_6341 = mux_6341(v_6308);
  assign v_6342 = mux_6342(v_6327);
  assign v_6344 = v_6345 | v_6364;
  assign v_6345 = act_6346 & 1'h1;
  assign act_6346 = v_6347 | v_6353;
  assign v_6347 = v_6348 & v_6354;
  assign v_6348 = v_6349 & vout_canPeek_6359;
  assign v_6349 = ~vout_canPeek_6350;
  pebbles_core
    pebbles_core_6350
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6351),
       .in0_consume_en(vin0_consume_en_6350),
       .out_canPeek(vout_canPeek_6350),
       .out_peek(vout_peek_6350));
  assign v_6351 = v_6352 | v_6357;
  assign v_6352 = mux_6352(v_6353);
  assign v_6353 = vout_canPeek_6350 & v_6354;
  assign v_6354 = v_6355 & 1'h1;
  assign v_6355 = v_6356 | 1'h0;
  assign v_6356 = ~v_6343;
  assign v_6357 = mux_6357(v_6358);
  assign v_6358 = ~v_6353;
  pebbles_core
    pebbles_core_6359
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6360),
       .in0_consume_en(vin0_consume_en_6359),
       .out_canPeek(vout_canPeek_6359),
       .out_peek(vout_peek_6359));
  assign v_6360 = v_6361 | v_6362;
  assign v_6361 = mux_6361(v_6347);
  assign v_6362 = mux_6362(v_6363);
  assign v_6363 = ~v_6347;
  assign v_6364 = v_6365 & 1'h1;
  assign v_6365 = v_6366 & v_6367;
  assign v_6366 = ~act_6346;
  assign v_6367 = v_6368 | v_6372;
  assign v_6368 = v_6369 | v_6370;
  assign v_6369 = mux_6369(v_6303);
  assign v_6370 = mux_6370(v_6371);
  assign v_6371 = ~v_6303;
  assign v_6372 = ~v_6343;
  assign v_6373 = v_6374 | v_6375;
  assign v_6374 = mux_6374(v_6345);
  assign v_6375 = mux_6375(v_6364);
  assign v_6376 = v_6377 & 1'h1;
  assign v_6377 = v_6378 & v_6379;
  assign v_6378 = ~act_6302;
  assign v_6379 = v_6380 | v_6384;
  assign v_6380 = v_6381 | v_6382;
  assign v_6381 = mux_6381(v_6203);
  assign v_6382 = mux_6382(v_6383);
  assign v_6383 = ~v_6203;
  assign v_6384 = ~v_6299;
  assign v_6385 = v_6386 | v_6387;
  assign v_6386 = mux_6386(v_6301);
  assign v_6387 = mux_6387(v_6376);
  assign v_6388 = v_6389 & 1'h1;
  assign v_6389 = v_6390 & v_6391;
  assign v_6390 = ~act_6202;
  assign v_6391 = v_6392 | v_6400;
  assign v_6392 = v_6393 | v_6398;
  assign v_6393 = mux_6393(v_6394);
  assign v_6394 = v_6199 & v_6395;
  assign v_6395 = v_6396 & 1'h1;
  assign v_6396 = v_6397 | 1'h0;
  assign v_6397 = ~v_6192;
  assign v_6398 = mux_6398(v_6399);
  assign v_6399 = ~v_6394;
  assign v_6400 = ~v_6199;
  assign v_6401 = v_6402 | v_6403;
  assign v_6402 = mux_6402(v_6201);
  assign v_6403 = mux_6403(v_6388);
  assign v_6405 = v_6406 | v_6593;
  assign v_6406 = act_6407 & 1'h1;
  assign act_6407 = v_6408 | v_6494;
  assign v_6408 = v_6409 & v_6495;
  assign v_6409 = v_6410 & v_6504;
  assign v_6410 = ~v_6411;
  assign v_6412 = v_6413 | v_6488;
  assign v_6413 = act_6414 & 1'h1;
  assign act_6414 = v_6415 | v_6445;
  assign v_6415 = v_6416 & v_6446;
  assign v_6416 = v_6417 & v_6455;
  assign v_6417 = ~v_6418;
  assign v_6419 = v_6420 | v_6439;
  assign v_6420 = act_6421 & 1'h1;
  assign act_6421 = v_6422 | v_6428;
  assign v_6422 = v_6423 & v_6429;
  assign v_6423 = v_6424 & vout_canPeek_6434;
  assign v_6424 = ~vout_canPeek_6425;
  pebbles_core
    pebbles_core_6425
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6426),
       .in0_consume_en(vin0_consume_en_6425),
       .out_canPeek(vout_canPeek_6425),
       .out_peek(vout_peek_6425));
  assign v_6426 = v_6427 | v_6432;
  assign v_6427 = mux_6427(v_6428);
  assign v_6428 = vout_canPeek_6425 & v_6429;
  assign v_6429 = v_6430 & 1'h1;
  assign v_6430 = v_6431 | 1'h0;
  assign v_6431 = ~v_6418;
  assign v_6432 = mux_6432(v_6433);
  assign v_6433 = ~v_6428;
  pebbles_core
    pebbles_core_6434
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6435),
       .in0_consume_en(vin0_consume_en_6434),
       .out_canPeek(vout_canPeek_6434),
       .out_peek(vout_peek_6434));
  assign v_6435 = v_6436 | v_6437;
  assign v_6436 = mux_6436(v_6422);
  assign v_6437 = mux_6437(v_6438);
  assign v_6438 = ~v_6422;
  assign v_6439 = v_6440 & 1'h1;
  assign v_6440 = v_6441 & v_6442;
  assign v_6441 = ~act_6421;
  assign v_6442 = v_6443 | v_6451;
  assign v_6443 = v_6444 | v_6449;
  assign v_6444 = mux_6444(v_6445);
  assign v_6445 = v_6418 & v_6446;
  assign v_6446 = v_6447 & 1'h1;
  assign v_6447 = v_6448 | 1'h0;
  assign v_6448 = ~v_6411;
  assign v_6449 = mux_6449(v_6450);
  assign v_6450 = ~v_6445;
  assign v_6451 = ~v_6418;
  assign v_6452 = v_6453 | v_6454;
  assign v_6453 = mux_6453(v_6420);
  assign v_6454 = mux_6454(v_6439);
  assign v_6456 = v_6457 | v_6476;
  assign v_6457 = act_6458 & 1'h1;
  assign act_6458 = v_6459 | v_6465;
  assign v_6459 = v_6460 & v_6466;
  assign v_6460 = v_6461 & vout_canPeek_6471;
  assign v_6461 = ~vout_canPeek_6462;
  pebbles_core
    pebbles_core_6462
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6463),
       .in0_consume_en(vin0_consume_en_6462),
       .out_canPeek(vout_canPeek_6462),
       .out_peek(vout_peek_6462));
  assign v_6463 = v_6464 | v_6469;
  assign v_6464 = mux_6464(v_6465);
  assign v_6465 = vout_canPeek_6462 & v_6466;
  assign v_6466 = v_6467 & 1'h1;
  assign v_6467 = v_6468 | 1'h0;
  assign v_6468 = ~v_6455;
  assign v_6469 = mux_6469(v_6470);
  assign v_6470 = ~v_6465;
  pebbles_core
    pebbles_core_6471
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6472),
       .in0_consume_en(vin0_consume_en_6471),
       .out_canPeek(vout_canPeek_6471),
       .out_peek(vout_peek_6471));
  assign v_6472 = v_6473 | v_6474;
  assign v_6473 = mux_6473(v_6459);
  assign v_6474 = mux_6474(v_6475);
  assign v_6475 = ~v_6459;
  assign v_6476 = v_6477 & 1'h1;
  assign v_6477 = v_6478 & v_6479;
  assign v_6478 = ~act_6458;
  assign v_6479 = v_6480 | v_6484;
  assign v_6480 = v_6481 | v_6482;
  assign v_6481 = mux_6481(v_6415);
  assign v_6482 = mux_6482(v_6483);
  assign v_6483 = ~v_6415;
  assign v_6484 = ~v_6455;
  assign v_6485 = v_6486 | v_6487;
  assign v_6486 = mux_6486(v_6457);
  assign v_6487 = mux_6487(v_6476);
  assign v_6488 = v_6489 & 1'h1;
  assign v_6489 = v_6490 & v_6491;
  assign v_6490 = ~act_6414;
  assign v_6491 = v_6492 | v_6500;
  assign v_6492 = v_6493 | v_6498;
  assign v_6493 = mux_6493(v_6494);
  assign v_6494 = v_6411 & v_6495;
  assign v_6495 = v_6496 & 1'h1;
  assign v_6496 = v_6497 | 1'h0;
  assign v_6497 = ~v_6404;
  assign v_6498 = mux_6498(v_6499);
  assign v_6499 = ~v_6494;
  assign v_6500 = ~v_6411;
  assign v_6501 = v_6502 | v_6503;
  assign v_6502 = mux_6502(v_6413);
  assign v_6503 = mux_6503(v_6488);
  assign v_6505 = v_6506 | v_6581;
  assign v_6506 = act_6507 & 1'h1;
  assign act_6507 = v_6508 | v_6538;
  assign v_6508 = v_6509 & v_6539;
  assign v_6509 = v_6510 & v_6548;
  assign v_6510 = ~v_6511;
  assign v_6512 = v_6513 | v_6532;
  assign v_6513 = act_6514 & 1'h1;
  assign act_6514 = v_6515 | v_6521;
  assign v_6515 = v_6516 & v_6522;
  assign v_6516 = v_6517 & vout_canPeek_6527;
  assign v_6517 = ~vout_canPeek_6518;
  pebbles_core
    pebbles_core_6518
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6519),
       .in0_consume_en(vin0_consume_en_6518),
       .out_canPeek(vout_canPeek_6518),
       .out_peek(vout_peek_6518));
  assign v_6519 = v_6520 | v_6525;
  assign v_6520 = mux_6520(v_6521);
  assign v_6521 = vout_canPeek_6518 & v_6522;
  assign v_6522 = v_6523 & 1'h1;
  assign v_6523 = v_6524 | 1'h0;
  assign v_6524 = ~v_6511;
  assign v_6525 = mux_6525(v_6526);
  assign v_6526 = ~v_6521;
  pebbles_core
    pebbles_core_6527
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6528),
       .in0_consume_en(vin0_consume_en_6527),
       .out_canPeek(vout_canPeek_6527),
       .out_peek(vout_peek_6527));
  assign v_6528 = v_6529 | v_6530;
  assign v_6529 = mux_6529(v_6515);
  assign v_6530 = mux_6530(v_6531);
  assign v_6531 = ~v_6515;
  assign v_6532 = v_6533 & 1'h1;
  assign v_6533 = v_6534 & v_6535;
  assign v_6534 = ~act_6514;
  assign v_6535 = v_6536 | v_6544;
  assign v_6536 = v_6537 | v_6542;
  assign v_6537 = mux_6537(v_6538);
  assign v_6538 = v_6511 & v_6539;
  assign v_6539 = v_6540 & 1'h1;
  assign v_6540 = v_6541 | 1'h0;
  assign v_6541 = ~v_6504;
  assign v_6542 = mux_6542(v_6543);
  assign v_6543 = ~v_6538;
  assign v_6544 = ~v_6511;
  assign v_6545 = v_6546 | v_6547;
  assign v_6546 = mux_6546(v_6513);
  assign v_6547 = mux_6547(v_6532);
  assign v_6549 = v_6550 | v_6569;
  assign v_6550 = act_6551 & 1'h1;
  assign act_6551 = v_6552 | v_6558;
  assign v_6552 = v_6553 & v_6559;
  assign v_6553 = v_6554 & vout_canPeek_6564;
  assign v_6554 = ~vout_canPeek_6555;
  pebbles_core
    pebbles_core_6555
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6556),
       .in0_consume_en(vin0_consume_en_6555),
       .out_canPeek(vout_canPeek_6555),
       .out_peek(vout_peek_6555));
  assign v_6556 = v_6557 | v_6562;
  assign v_6557 = mux_6557(v_6558);
  assign v_6558 = vout_canPeek_6555 & v_6559;
  assign v_6559 = v_6560 & 1'h1;
  assign v_6560 = v_6561 | 1'h0;
  assign v_6561 = ~v_6548;
  assign v_6562 = mux_6562(v_6563);
  assign v_6563 = ~v_6558;
  pebbles_core
    pebbles_core_6564
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6565),
       .in0_consume_en(vin0_consume_en_6564),
       .out_canPeek(vout_canPeek_6564),
       .out_peek(vout_peek_6564));
  assign v_6565 = v_6566 | v_6567;
  assign v_6566 = mux_6566(v_6552);
  assign v_6567 = mux_6567(v_6568);
  assign v_6568 = ~v_6552;
  assign v_6569 = v_6570 & 1'h1;
  assign v_6570 = v_6571 & v_6572;
  assign v_6571 = ~act_6551;
  assign v_6572 = v_6573 | v_6577;
  assign v_6573 = v_6574 | v_6575;
  assign v_6574 = mux_6574(v_6508);
  assign v_6575 = mux_6575(v_6576);
  assign v_6576 = ~v_6508;
  assign v_6577 = ~v_6548;
  assign v_6578 = v_6579 | v_6580;
  assign v_6579 = mux_6579(v_6550);
  assign v_6580 = mux_6580(v_6569);
  assign v_6581 = v_6582 & 1'h1;
  assign v_6582 = v_6583 & v_6584;
  assign v_6583 = ~act_6507;
  assign v_6584 = v_6585 | v_6589;
  assign v_6585 = v_6586 | v_6587;
  assign v_6586 = mux_6586(v_6408);
  assign v_6587 = mux_6587(v_6588);
  assign v_6588 = ~v_6408;
  assign v_6589 = ~v_6504;
  assign v_6590 = v_6591 | v_6592;
  assign v_6591 = mux_6591(v_6506);
  assign v_6592 = mux_6592(v_6581);
  assign v_6593 = v_6594 & 1'h1;
  assign v_6594 = v_6595 & v_6596;
  assign v_6595 = ~act_6407;
  assign v_6596 = v_6597 | v_6601;
  assign v_6597 = v_6598 | v_6599;
  assign v_6598 = mux_6598(v_6196);
  assign v_6599 = mux_6599(v_6600);
  assign v_6600 = ~v_6196;
  assign v_6601 = ~v_6404;
  assign v_6602 = v_6603 | v_6604;
  assign v_6603 = mux_6603(v_6406);
  assign v_6604 = mux_6604(v_6593);
  assign v_6605 = v_6606 & 1'h1;
  assign v_6606 = v_6607 & v_6608;
  assign v_6607 = ~act_6195;
  assign v_6608 = v_6609 | v_6617;
  assign v_6609 = v_6610 | v_6615;
  assign v_6610 = mux_6610(v_6611);
  assign v_6611 = v_6192 & v_6612;
  assign v_6612 = v_6613 & 1'h1;
  assign v_6613 = v_6614 | 1'h0;
  assign v_6614 = ~v_6185;
  assign v_6615 = mux_6615(v_6616);
  assign v_6616 = ~v_6611;
  assign v_6617 = ~v_6192;
  assign v_6618 = v_6619 | v_6620;
  assign v_6619 = mux_6619(v_6194);
  assign v_6620 = mux_6620(v_6605);
  assign v_6622 = v_6623 | v_7034;
  assign v_6623 = act_6624 & 1'h1;
  assign act_6624 = v_6625 | v_6823;
  assign v_6625 = v_6626 & v_6824;
  assign v_6626 = v_6627 & v_6833;
  assign v_6627 = ~v_6628;
  assign v_6629 = v_6630 | v_6817;
  assign v_6630 = act_6631 & 1'h1;
  assign act_6631 = v_6632 | v_6718;
  assign v_6632 = v_6633 & v_6719;
  assign v_6633 = v_6634 & v_6728;
  assign v_6634 = ~v_6635;
  assign v_6636 = v_6637 | v_6712;
  assign v_6637 = act_6638 & 1'h1;
  assign act_6638 = v_6639 | v_6669;
  assign v_6639 = v_6640 & v_6670;
  assign v_6640 = v_6641 & v_6679;
  assign v_6641 = ~v_6642;
  assign v_6643 = v_6644 | v_6663;
  assign v_6644 = act_6645 & 1'h1;
  assign act_6645 = v_6646 | v_6652;
  assign v_6646 = v_6647 & v_6653;
  assign v_6647 = v_6648 & vout_canPeek_6658;
  assign v_6648 = ~vout_canPeek_6649;
  pebbles_core
    pebbles_core_6649
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6650),
       .in0_consume_en(vin0_consume_en_6649),
       .out_canPeek(vout_canPeek_6649),
       .out_peek(vout_peek_6649));
  assign v_6650 = v_6651 | v_6656;
  assign v_6651 = mux_6651(v_6652);
  assign v_6652 = vout_canPeek_6649 & v_6653;
  assign v_6653 = v_6654 & 1'h1;
  assign v_6654 = v_6655 | 1'h0;
  assign v_6655 = ~v_6642;
  assign v_6656 = mux_6656(v_6657);
  assign v_6657 = ~v_6652;
  pebbles_core
    pebbles_core_6658
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6659),
       .in0_consume_en(vin0_consume_en_6658),
       .out_canPeek(vout_canPeek_6658),
       .out_peek(vout_peek_6658));
  assign v_6659 = v_6660 | v_6661;
  assign v_6660 = mux_6660(v_6646);
  assign v_6661 = mux_6661(v_6662);
  assign v_6662 = ~v_6646;
  assign v_6663 = v_6664 & 1'h1;
  assign v_6664 = v_6665 & v_6666;
  assign v_6665 = ~act_6645;
  assign v_6666 = v_6667 | v_6675;
  assign v_6667 = v_6668 | v_6673;
  assign v_6668 = mux_6668(v_6669);
  assign v_6669 = v_6642 & v_6670;
  assign v_6670 = v_6671 & 1'h1;
  assign v_6671 = v_6672 | 1'h0;
  assign v_6672 = ~v_6635;
  assign v_6673 = mux_6673(v_6674);
  assign v_6674 = ~v_6669;
  assign v_6675 = ~v_6642;
  assign v_6676 = v_6677 | v_6678;
  assign v_6677 = mux_6677(v_6644);
  assign v_6678 = mux_6678(v_6663);
  assign v_6680 = v_6681 | v_6700;
  assign v_6681 = act_6682 & 1'h1;
  assign act_6682 = v_6683 | v_6689;
  assign v_6683 = v_6684 & v_6690;
  assign v_6684 = v_6685 & vout_canPeek_6695;
  assign v_6685 = ~vout_canPeek_6686;
  pebbles_core
    pebbles_core_6686
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6687),
       .in0_consume_en(vin0_consume_en_6686),
       .out_canPeek(vout_canPeek_6686),
       .out_peek(vout_peek_6686));
  assign v_6687 = v_6688 | v_6693;
  assign v_6688 = mux_6688(v_6689);
  assign v_6689 = vout_canPeek_6686 & v_6690;
  assign v_6690 = v_6691 & 1'h1;
  assign v_6691 = v_6692 | 1'h0;
  assign v_6692 = ~v_6679;
  assign v_6693 = mux_6693(v_6694);
  assign v_6694 = ~v_6689;
  pebbles_core
    pebbles_core_6695
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6696),
       .in0_consume_en(vin0_consume_en_6695),
       .out_canPeek(vout_canPeek_6695),
       .out_peek(vout_peek_6695));
  assign v_6696 = v_6697 | v_6698;
  assign v_6697 = mux_6697(v_6683);
  assign v_6698 = mux_6698(v_6699);
  assign v_6699 = ~v_6683;
  assign v_6700 = v_6701 & 1'h1;
  assign v_6701 = v_6702 & v_6703;
  assign v_6702 = ~act_6682;
  assign v_6703 = v_6704 | v_6708;
  assign v_6704 = v_6705 | v_6706;
  assign v_6705 = mux_6705(v_6639);
  assign v_6706 = mux_6706(v_6707);
  assign v_6707 = ~v_6639;
  assign v_6708 = ~v_6679;
  assign v_6709 = v_6710 | v_6711;
  assign v_6710 = mux_6710(v_6681);
  assign v_6711 = mux_6711(v_6700);
  assign v_6712 = v_6713 & 1'h1;
  assign v_6713 = v_6714 & v_6715;
  assign v_6714 = ~act_6638;
  assign v_6715 = v_6716 | v_6724;
  assign v_6716 = v_6717 | v_6722;
  assign v_6717 = mux_6717(v_6718);
  assign v_6718 = v_6635 & v_6719;
  assign v_6719 = v_6720 & 1'h1;
  assign v_6720 = v_6721 | 1'h0;
  assign v_6721 = ~v_6628;
  assign v_6722 = mux_6722(v_6723);
  assign v_6723 = ~v_6718;
  assign v_6724 = ~v_6635;
  assign v_6725 = v_6726 | v_6727;
  assign v_6726 = mux_6726(v_6637);
  assign v_6727 = mux_6727(v_6712);
  assign v_6729 = v_6730 | v_6805;
  assign v_6730 = act_6731 & 1'h1;
  assign act_6731 = v_6732 | v_6762;
  assign v_6732 = v_6733 & v_6763;
  assign v_6733 = v_6734 & v_6772;
  assign v_6734 = ~v_6735;
  assign v_6736 = v_6737 | v_6756;
  assign v_6737 = act_6738 & 1'h1;
  assign act_6738 = v_6739 | v_6745;
  assign v_6739 = v_6740 & v_6746;
  assign v_6740 = v_6741 & vout_canPeek_6751;
  assign v_6741 = ~vout_canPeek_6742;
  pebbles_core
    pebbles_core_6742
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6743),
       .in0_consume_en(vin0_consume_en_6742),
       .out_canPeek(vout_canPeek_6742),
       .out_peek(vout_peek_6742));
  assign v_6743 = v_6744 | v_6749;
  assign v_6744 = mux_6744(v_6745);
  assign v_6745 = vout_canPeek_6742 & v_6746;
  assign v_6746 = v_6747 & 1'h1;
  assign v_6747 = v_6748 | 1'h0;
  assign v_6748 = ~v_6735;
  assign v_6749 = mux_6749(v_6750);
  assign v_6750 = ~v_6745;
  pebbles_core
    pebbles_core_6751
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6752),
       .in0_consume_en(vin0_consume_en_6751),
       .out_canPeek(vout_canPeek_6751),
       .out_peek(vout_peek_6751));
  assign v_6752 = v_6753 | v_6754;
  assign v_6753 = mux_6753(v_6739);
  assign v_6754 = mux_6754(v_6755);
  assign v_6755 = ~v_6739;
  assign v_6756 = v_6757 & 1'h1;
  assign v_6757 = v_6758 & v_6759;
  assign v_6758 = ~act_6738;
  assign v_6759 = v_6760 | v_6768;
  assign v_6760 = v_6761 | v_6766;
  assign v_6761 = mux_6761(v_6762);
  assign v_6762 = v_6735 & v_6763;
  assign v_6763 = v_6764 & 1'h1;
  assign v_6764 = v_6765 | 1'h0;
  assign v_6765 = ~v_6728;
  assign v_6766 = mux_6766(v_6767);
  assign v_6767 = ~v_6762;
  assign v_6768 = ~v_6735;
  assign v_6769 = v_6770 | v_6771;
  assign v_6770 = mux_6770(v_6737);
  assign v_6771 = mux_6771(v_6756);
  assign v_6773 = v_6774 | v_6793;
  assign v_6774 = act_6775 & 1'h1;
  assign act_6775 = v_6776 | v_6782;
  assign v_6776 = v_6777 & v_6783;
  assign v_6777 = v_6778 & vout_canPeek_6788;
  assign v_6778 = ~vout_canPeek_6779;
  pebbles_core
    pebbles_core_6779
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6780),
       .in0_consume_en(vin0_consume_en_6779),
       .out_canPeek(vout_canPeek_6779),
       .out_peek(vout_peek_6779));
  assign v_6780 = v_6781 | v_6786;
  assign v_6781 = mux_6781(v_6782);
  assign v_6782 = vout_canPeek_6779 & v_6783;
  assign v_6783 = v_6784 & 1'h1;
  assign v_6784 = v_6785 | 1'h0;
  assign v_6785 = ~v_6772;
  assign v_6786 = mux_6786(v_6787);
  assign v_6787 = ~v_6782;
  pebbles_core
    pebbles_core_6788
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6789),
       .in0_consume_en(vin0_consume_en_6788),
       .out_canPeek(vout_canPeek_6788),
       .out_peek(vout_peek_6788));
  assign v_6789 = v_6790 | v_6791;
  assign v_6790 = mux_6790(v_6776);
  assign v_6791 = mux_6791(v_6792);
  assign v_6792 = ~v_6776;
  assign v_6793 = v_6794 & 1'h1;
  assign v_6794 = v_6795 & v_6796;
  assign v_6795 = ~act_6775;
  assign v_6796 = v_6797 | v_6801;
  assign v_6797 = v_6798 | v_6799;
  assign v_6798 = mux_6798(v_6732);
  assign v_6799 = mux_6799(v_6800);
  assign v_6800 = ~v_6732;
  assign v_6801 = ~v_6772;
  assign v_6802 = v_6803 | v_6804;
  assign v_6803 = mux_6803(v_6774);
  assign v_6804 = mux_6804(v_6793);
  assign v_6805 = v_6806 & 1'h1;
  assign v_6806 = v_6807 & v_6808;
  assign v_6807 = ~act_6731;
  assign v_6808 = v_6809 | v_6813;
  assign v_6809 = v_6810 | v_6811;
  assign v_6810 = mux_6810(v_6632);
  assign v_6811 = mux_6811(v_6812);
  assign v_6812 = ~v_6632;
  assign v_6813 = ~v_6728;
  assign v_6814 = v_6815 | v_6816;
  assign v_6815 = mux_6815(v_6730);
  assign v_6816 = mux_6816(v_6805);
  assign v_6817 = v_6818 & 1'h1;
  assign v_6818 = v_6819 & v_6820;
  assign v_6819 = ~act_6631;
  assign v_6820 = v_6821 | v_6829;
  assign v_6821 = v_6822 | v_6827;
  assign v_6822 = mux_6822(v_6823);
  assign v_6823 = v_6628 & v_6824;
  assign v_6824 = v_6825 & 1'h1;
  assign v_6825 = v_6826 | 1'h0;
  assign v_6826 = ~v_6621;
  assign v_6827 = mux_6827(v_6828);
  assign v_6828 = ~v_6823;
  assign v_6829 = ~v_6628;
  assign v_6830 = v_6831 | v_6832;
  assign v_6831 = mux_6831(v_6630);
  assign v_6832 = mux_6832(v_6817);
  assign v_6834 = v_6835 | v_7022;
  assign v_6835 = act_6836 & 1'h1;
  assign act_6836 = v_6837 | v_6923;
  assign v_6837 = v_6838 & v_6924;
  assign v_6838 = v_6839 & v_6933;
  assign v_6839 = ~v_6840;
  assign v_6841 = v_6842 | v_6917;
  assign v_6842 = act_6843 & 1'h1;
  assign act_6843 = v_6844 | v_6874;
  assign v_6844 = v_6845 & v_6875;
  assign v_6845 = v_6846 & v_6884;
  assign v_6846 = ~v_6847;
  assign v_6848 = v_6849 | v_6868;
  assign v_6849 = act_6850 & 1'h1;
  assign act_6850 = v_6851 | v_6857;
  assign v_6851 = v_6852 & v_6858;
  assign v_6852 = v_6853 & vout_canPeek_6863;
  assign v_6853 = ~vout_canPeek_6854;
  pebbles_core
    pebbles_core_6854
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6855),
       .in0_consume_en(vin0_consume_en_6854),
       .out_canPeek(vout_canPeek_6854),
       .out_peek(vout_peek_6854));
  assign v_6855 = v_6856 | v_6861;
  assign v_6856 = mux_6856(v_6857);
  assign v_6857 = vout_canPeek_6854 & v_6858;
  assign v_6858 = v_6859 & 1'h1;
  assign v_6859 = v_6860 | 1'h0;
  assign v_6860 = ~v_6847;
  assign v_6861 = mux_6861(v_6862);
  assign v_6862 = ~v_6857;
  pebbles_core
    pebbles_core_6863
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6864),
       .in0_consume_en(vin0_consume_en_6863),
       .out_canPeek(vout_canPeek_6863),
       .out_peek(vout_peek_6863));
  assign v_6864 = v_6865 | v_6866;
  assign v_6865 = mux_6865(v_6851);
  assign v_6866 = mux_6866(v_6867);
  assign v_6867 = ~v_6851;
  assign v_6868 = v_6869 & 1'h1;
  assign v_6869 = v_6870 & v_6871;
  assign v_6870 = ~act_6850;
  assign v_6871 = v_6872 | v_6880;
  assign v_6872 = v_6873 | v_6878;
  assign v_6873 = mux_6873(v_6874);
  assign v_6874 = v_6847 & v_6875;
  assign v_6875 = v_6876 & 1'h1;
  assign v_6876 = v_6877 | 1'h0;
  assign v_6877 = ~v_6840;
  assign v_6878 = mux_6878(v_6879);
  assign v_6879 = ~v_6874;
  assign v_6880 = ~v_6847;
  assign v_6881 = v_6882 | v_6883;
  assign v_6882 = mux_6882(v_6849);
  assign v_6883 = mux_6883(v_6868);
  assign v_6885 = v_6886 | v_6905;
  assign v_6886 = act_6887 & 1'h1;
  assign act_6887 = v_6888 | v_6894;
  assign v_6888 = v_6889 & v_6895;
  assign v_6889 = v_6890 & vout_canPeek_6900;
  assign v_6890 = ~vout_canPeek_6891;
  pebbles_core
    pebbles_core_6891
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6892),
       .in0_consume_en(vin0_consume_en_6891),
       .out_canPeek(vout_canPeek_6891),
       .out_peek(vout_peek_6891));
  assign v_6892 = v_6893 | v_6898;
  assign v_6893 = mux_6893(v_6894);
  assign v_6894 = vout_canPeek_6891 & v_6895;
  assign v_6895 = v_6896 & 1'h1;
  assign v_6896 = v_6897 | 1'h0;
  assign v_6897 = ~v_6884;
  assign v_6898 = mux_6898(v_6899);
  assign v_6899 = ~v_6894;
  pebbles_core
    pebbles_core_6900
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6901),
       .in0_consume_en(vin0_consume_en_6900),
       .out_canPeek(vout_canPeek_6900),
       .out_peek(vout_peek_6900));
  assign v_6901 = v_6902 | v_6903;
  assign v_6902 = mux_6902(v_6888);
  assign v_6903 = mux_6903(v_6904);
  assign v_6904 = ~v_6888;
  assign v_6905 = v_6906 & 1'h1;
  assign v_6906 = v_6907 & v_6908;
  assign v_6907 = ~act_6887;
  assign v_6908 = v_6909 | v_6913;
  assign v_6909 = v_6910 | v_6911;
  assign v_6910 = mux_6910(v_6844);
  assign v_6911 = mux_6911(v_6912);
  assign v_6912 = ~v_6844;
  assign v_6913 = ~v_6884;
  assign v_6914 = v_6915 | v_6916;
  assign v_6915 = mux_6915(v_6886);
  assign v_6916 = mux_6916(v_6905);
  assign v_6917 = v_6918 & 1'h1;
  assign v_6918 = v_6919 & v_6920;
  assign v_6919 = ~act_6843;
  assign v_6920 = v_6921 | v_6929;
  assign v_6921 = v_6922 | v_6927;
  assign v_6922 = mux_6922(v_6923);
  assign v_6923 = v_6840 & v_6924;
  assign v_6924 = v_6925 & 1'h1;
  assign v_6925 = v_6926 | 1'h0;
  assign v_6926 = ~v_6833;
  assign v_6927 = mux_6927(v_6928);
  assign v_6928 = ~v_6923;
  assign v_6929 = ~v_6840;
  assign v_6930 = v_6931 | v_6932;
  assign v_6931 = mux_6931(v_6842);
  assign v_6932 = mux_6932(v_6917);
  assign v_6934 = v_6935 | v_7010;
  assign v_6935 = act_6936 & 1'h1;
  assign act_6936 = v_6937 | v_6967;
  assign v_6937 = v_6938 & v_6968;
  assign v_6938 = v_6939 & v_6977;
  assign v_6939 = ~v_6940;
  assign v_6941 = v_6942 | v_6961;
  assign v_6942 = act_6943 & 1'h1;
  assign act_6943 = v_6944 | v_6950;
  assign v_6944 = v_6945 & v_6951;
  assign v_6945 = v_6946 & vout_canPeek_6956;
  assign v_6946 = ~vout_canPeek_6947;
  pebbles_core
    pebbles_core_6947
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6948),
       .in0_consume_en(vin0_consume_en_6947),
       .out_canPeek(vout_canPeek_6947),
       .out_peek(vout_peek_6947));
  assign v_6948 = v_6949 | v_6954;
  assign v_6949 = mux_6949(v_6950);
  assign v_6950 = vout_canPeek_6947 & v_6951;
  assign v_6951 = v_6952 & 1'h1;
  assign v_6952 = v_6953 | 1'h0;
  assign v_6953 = ~v_6940;
  assign v_6954 = mux_6954(v_6955);
  assign v_6955 = ~v_6950;
  pebbles_core
    pebbles_core_6956
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6957),
       .in0_consume_en(vin0_consume_en_6956),
       .out_canPeek(vout_canPeek_6956),
       .out_peek(vout_peek_6956));
  assign v_6957 = v_6958 | v_6959;
  assign v_6958 = mux_6958(v_6944);
  assign v_6959 = mux_6959(v_6960);
  assign v_6960 = ~v_6944;
  assign v_6961 = v_6962 & 1'h1;
  assign v_6962 = v_6963 & v_6964;
  assign v_6963 = ~act_6943;
  assign v_6964 = v_6965 | v_6973;
  assign v_6965 = v_6966 | v_6971;
  assign v_6966 = mux_6966(v_6967);
  assign v_6967 = v_6940 & v_6968;
  assign v_6968 = v_6969 & 1'h1;
  assign v_6969 = v_6970 | 1'h0;
  assign v_6970 = ~v_6933;
  assign v_6971 = mux_6971(v_6972);
  assign v_6972 = ~v_6967;
  assign v_6973 = ~v_6940;
  assign v_6974 = v_6975 | v_6976;
  assign v_6975 = mux_6975(v_6942);
  assign v_6976 = mux_6976(v_6961);
  assign v_6978 = v_6979 | v_6998;
  assign v_6979 = act_6980 & 1'h1;
  assign act_6980 = v_6981 | v_6987;
  assign v_6981 = v_6982 & v_6988;
  assign v_6982 = v_6983 & vout_canPeek_6993;
  assign v_6983 = ~vout_canPeek_6984;
  pebbles_core
    pebbles_core_6984
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6985),
       .in0_consume_en(vin0_consume_en_6984),
       .out_canPeek(vout_canPeek_6984),
       .out_peek(vout_peek_6984));
  assign v_6985 = v_6986 | v_6991;
  assign v_6986 = mux_6986(v_6987);
  assign v_6987 = vout_canPeek_6984 & v_6988;
  assign v_6988 = v_6989 & 1'h1;
  assign v_6989 = v_6990 | 1'h0;
  assign v_6990 = ~v_6977;
  assign v_6991 = mux_6991(v_6992);
  assign v_6992 = ~v_6987;
  pebbles_core
    pebbles_core_6993
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6994),
       .in0_consume_en(vin0_consume_en_6993),
       .out_canPeek(vout_canPeek_6993),
       .out_peek(vout_peek_6993));
  assign v_6994 = v_6995 | v_6996;
  assign v_6995 = mux_6995(v_6981);
  assign v_6996 = mux_6996(v_6997);
  assign v_6997 = ~v_6981;
  assign v_6998 = v_6999 & 1'h1;
  assign v_6999 = v_7000 & v_7001;
  assign v_7000 = ~act_6980;
  assign v_7001 = v_7002 | v_7006;
  assign v_7002 = v_7003 | v_7004;
  assign v_7003 = mux_7003(v_6937);
  assign v_7004 = mux_7004(v_7005);
  assign v_7005 = ~v_6937;
  assign v_7006 = ~v_6977;
  assign v_7007 = v_7008 | v_7009;
  assign v_7008 = mux_7008(v_6979);
  assign v_7009 = mux_7009(v_6998);
  assign v_7010 = v_7011 & 1'h1;
  assign v_7011 = v_7012 & v_7013;
  assign v_7012 = ~act_6936;
  assign v_7013 = v_7014 | v_7018;
  assign v_7014 = v_7015 | v_7016;
  assign v_7015 = mux_7015(v_6837);
  assign v_7016 = mux_7016(v_7017);
  assign v_7017 = ~v_6837;
  assign v_7018 = ~v_6933;
  assign v_7019 = v_7020 | v_7021;
  assign v_7020 = mux_7020(v_6935);
  assign v_7021 = mux_7021(v_7010);
  assign v_7022 = v_7023 & 1'h1;
  assign v_7023 = v_7024 & v_7025;
  assign v_7024 = ~act_6836;
  assign v_7025 = v_7026 | v_7030;
  assign v_7026 = v_7027 | v_7028;
  assign v_7027 = mux_7027(v_6625);
  assign v_7028 = mux_7028(v_7029);
  assign v_7029 = ~v_6625;
  assign v_7030 = ~v_6833;
  assign v_7031 = v_7032 | v_7033;
  assign v_7032 = mux_7032(v_6835);
  assign v_7033 = mux_7033(v_7022);
  assign v_7034 = v_7035 & 1'h1;
  assign v_7035 = v_7036 & v_7037;
  assign v_7036 = ~act_6624;
  assign v_7037 = v_7038 | v_7042;
  assign v_7038 = v_7039 | v_7040;
  assign v_7039 = mux_7039(v_6189);
  assign v_7040 = mux_7040(v_7041);
  assign v_7041 = ~v_6189;
  assign v_7042 = ~v_6621;
  assign v_7043 = v_7044 | v_7045;
  assign v_7044 = mux_7044(v_6623);
  assign v_7045 = mux_7045(v_7034);
  assign v_7046 = v_7047 & 1'h1;
  assign v_7047 = v_7048 & v_7049;
  assign v_7048 = ~act_6188;
  assign v_7049 = v_7050 | v_7058;
  assign v_7050 = v_7051 | v_7056;
  assign v_7051 = mux_7051(v_7052);
  assign v_7052 = v_6185 & v_7053;
  assign v_7053 = v_7054 & 1'h1;
  assign v_7054 = v_7055 | 1'h0;
  assign v_7055 = ~v_6178;
  assign v_7056 = mux_7056(v_7057);
  assign v_7057 = ~v_7052;
  assign v_7058 = ~v_6185;
  assign v_7059 = v_7060 | v_7061;
  assign v_7060 = mux_7060(v_6187);
  assign v_7061 = mux_7061(v_7046);
  assign v_7063 = v_7064 | v_7923;
  assign v_7064 = act_7065 & 1'h1;
  assign act_7065 = v_7066 | v_7488;
  assign v_7066 = v_7067 & v_7489;
  assign v_7067 = v_7068 & v_7498;
  assign v_7068 = ~v_7069;
  assign v_7070 = v_7071 | v_7482;
  assign v_7071 = act_7072 & 1'h1;
  assign act_7072 = v_7073 | v_7271;
  assign v_7073 = v_7074 & v_7272;
  assign v_7074 = v_7075 & v_7281;
  assign v_7075 = ~v_7076;
  assign v_7077 = v_7078 | v_7265;
  assign v_7078 = act_7079 & 1'h1;
  assign act_7079 = v_7080 | v_7166;
  assign v_7080 = v_7081 & v_7167;
  assign v_7081 = v_7082 & v_7176;
  assign v_7082 = ~v_7083;
  assign v_7084 = v_7085 | v_7160;
  assign v_7085 = act_7086 & 1'h1;
  assign act_7086 = v_7087 | v_7117;
  assign v_7087 = v_7088 & v_7118;
  assign v_7088 = v_7089 & v_7127;
  assign v_7089 = ~v_7090;
  assign v_7091 = v_7092 | v_7111;
  assign v_7092 = act_7093 & 1'h1;
  assign act_7093 = v_7094 | v_7100;
  assign v_7094 = v_7095 & v_7101;
  assign v_7095 = v_7096 & vout_canPeek_7106;
  assign v_7096 = ~vout_canPeek_7097;
  pebbles_core
    pebbles_core_7097
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7098),
       .in0_consume_en(vin0_consume_en_7097),
       .out_canPeek(vout_canPeek_7097),
       .out_peek(vout_peek_7097));
  assign v_7098 = v_7099 | v_7104;
  assign v_7099 = mux_7099(v_7100);
  assign v_7100 = vout_canPeek_7097 & v_7101;
  assign v_7101 = v_7102 & 1'h1;
  assign v_7102 = v_7103 | 1'h0;
  assign v_7103 = ~v_7090;
  assign v_7104 = mux_7104(v_7105);
  assign v_7105 = ~v_7100;
  pebbles_core
    pebbles_core_7106
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7107),
       .in0_consume_en(vin0_consume_en_7106),
       .out_canPeek(vout_canPeek_7106),
       .out_peek(vout_peek_7106));
  assign v_7107 = v_7108 | v_7109;
  assign v_7108 = mux_7108(v_7094);
  assign v_7109 = mux_7109(v_7110);
  assign v_7110 = ~v_7094;
  assign v_7111 = v_7112 & 1'h1;
  assign v_7112 = v_7113 & v_7114;
  assign v_7113 = ~act_7093;
  assign v_7114 = v_7115 | v_7123;
  assign v_7115 = v_7116 | v_7121;
  assign v_7116 = mux_7116(v_7117);
  assign v_7117 = v_7090 & v_7118;
  assign v_7118 = v_7119 & 1'h1;
  assign v_7119 = v_7120 | 1'h0;
  assign v_7120 = ~v_7083;
  assign v_7121 = mux_7121(v_7122);
  assign v_7122 = ~v_7117;
  assign v_7123 = ~v_7090;
  assign v_7124 = v_7125 | v_7126;
  assign v_7125 = mux_7125(v_7092);
  assign v_7126 = mux_7126(v_7111);
  assign v_7128 = v_7129 | v_7148;
  assign v_7129 = act_7130 & 1'h1;
  assign act_7130 = v_7131 | v_7137;
  assign v_7131 = v_7132 & v_7138;
  assign v_7132 = v_7133 & vout_canPeek_7143;
  assign v_7133 = ~vout_canPeek_7134;
  pebbles_core
    pebbles_core_7134
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7135),
       .in0_consume_en(vin0_consume_en_7134),
       .out_canPeek(vout_canPeek_7134),
       .out_peek(vout_peek_7134));
  assign v_7135 = v_7136 | v_7141;
  assign v_7136 = mux_7136(v_7137);
  assign v_7137 = vout_canPeek_7134 & v_7138;
  assign v_7138 = v_7139 & 1'h1;
  assign v_7139 = v_7140 | 1'h0;
  assign v_7140 = ~v_7127;
  assign v_7141 = mux_7141(v_7142);
  assign v_7142 = ~v_7137;
  pebbles_core
    pebbles_core_7143
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7144),
       .in0_consume_en(vin0_consume_en_7143),
       .out_canPeek(vout_canPeek_7143),
       .out_peek(vout_peek_7143));
  assign v_7144 = v_7145 | v_7146;
  assign v_7145 = mux_7145(v_7131);
  assign v_7146 = mux_7146(v_7147);
  assign v_7147 = ~v_7131;
  assign v_7148 = v_7149 & 1'h1;
  assign v_7149 = v_7150 & v_7151;
  assign v_7150 = ~act_7130;
  assign v_7151 = v_7152 | v_7156;
  assign v_7152 = v_7153 | v_7154;
  assign v_7153 = mux_7153(v_7087);
  assign v_7154 = mux_7154(v_7155);
  assign v_7155 = ~v_7087;
  assign v_7156 = ~v_7127;
  assign v_7157 = v_7158 | v_7159;
  assign v_7158 = mux_7158(v_7129);
  assign v_7159 = mux_7159(v_7148);
  assign v_7160 = v_7161 & 1'h1;
  assign v_7161 = v_7162 & v_7163;
  assign v_7162 = ~act_7086;
  assign v_7163 = v_7164 | v_7172;
  assign v_7164 = v_7165 | v_7170;
  assign v_7165 = mux_7165(v_7166);
  assign v_7166 = v_7083 & v_7167;
  assign v_7167 = v_7168 & 1'h1;
  assign v_7168 = v_7169 | 1'h0;
  assign v_7169 = ~v_7076;
  assign v_7170 = mux_7170(v_7171);
  assign v_7171 = ~v_7166;
  assign v_7172 = ~v_7083;
  assign v_7173 = v_7174 | v_7175;
  assign v_7174 = mux_7174(v_7085);
  assign v_7175 = mux_7175(v_7160);
  assign v_7177 = v_7178 | v_7253;
  assign v_7178 = act_7179 & 1'h1;
  assign act_7179 = v_7180 | v_7210;
  assign v_7180 = v_7181 & v_7211;
  assign v_7181 = v_7182 & v_7220;
  assign v_7182 = ~v_7183;
  assign v_7184 = v_7185 | v_7204;
  assign v_7185 = act_7186 & 1'h1;
  assign act_7186 = v_7187 | v_7193;
  assign v_7187 = v_7188 & v_7194;
  assign v_7188 = v_7189 & vout_canPeek_7199;
  assign v_7189 = ~vout_canPeek_7190;
  pebbles_core
    pebbles_core_7190
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7191),
       .in0_consume_en(vin0_consume_en_7190),
       .out_canPeek(vout_canPeek_7190),
       .out_peek(vout_peek_7190));
  assign v_7191 = v_7192 | v_7197;
  assign v_7192 = mux_7192(v_7193);
  assign v_7193 = vout_canPeek_7190 & v_7194;
  assign v_7194 = v_7195 & 1'h1;
  assign v_7195 = v_7196 | 1'h0;
  assign v_7196 = ~v_7183;
  assign v_7197 = mux_7197(v_7198);
  assign v_7198 = ~v_7193;
  pebbles_core
    pebbles_core_7199
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7200),
       .in0_consume_en(vin0_consume_en_7199),
       .out_canPeek(vout_canPeek_7199),
       .out_peek(vout_peek_7199));
  assign v_7200 = v_7201 | v_7202;
  assign v_7201 = mux_7201(v_7187);
  assign v_7202 = mux_7202(v_7203);
  assign v_7203 = ~v_7187;
  assign v_7204 = v_7205 & 1'h1;
  assign v_7205 = v_7206 & v_7207;
  assign v_7206 = ~act_7186;
  assign v_7207 = v_7208 | v_7216;
  assign v_7208 = v_7209 | v_7214;
  assign v_7209 = mux_7209(v_7210);
  assign v_7210 = v_7183 & v_7211;
  assign v_7211 = v_7212 & 1'h1;
  assign v_7212 = v_7213 | 1'h0;
  assign v_7213 = ~v_7176;
  assign v_7214 = mux_7214(v_7215);
  assign v_7215 = ~v_7210;
  assign v_7216 = ~v_7183;
  assign v_7217 = v_7218 | v_7219;
  assign v_7218 = mux_7218(v_7185);
  assign v_7219 = mux_7219(v_7204);
  assign v_7221 = v_7222 | v_7241;
  assign v_7222 = act_7223 & 1'h1;
  assign act_7223 = v_7224 | v_7230;
  assign v_7224 = v_7225 & v_7231;
  assign v_7225 = v_7226 & vout_canPeek_7236;
  assign v_7226 = ~vout_canPeek_7227;
  pebbles_core
    pebbles_core_7227
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7228),
       .in0_consume_en(vin0_consume_en_7227),
       .out_canPeek(vout_canPeek_7227),
       .out_peek(vout_peek_7227));
  assign v_7228 = v_7229 | v_7234;
  assign v_7229 = mux_7229(v_7230);
  assign v_7230 = vout_canPeek_7227 & v_7231;
  assign v_7231 = v_7232 & 1'h1;
  assign v_7232 = v_7233 | 1'h0;
  assign v_7233 = ~v_7220;
  assign v_7234 = mux_7234(v_7235);
  assign v_7235 = ~v_7230;
  pebbles_core
    pebbles_core_7236
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7237),
       .in0_consume_en(vin0_consume_en_7236),
       .out_canPeek(vout_canPeek_7236),
       .out_peek(vout_peek_7236));
  assign v_7237 = v_7238 | v_7239;
  assign v_7238 = mux_7238(v_7224);
  assign v_7239 = mux_7239(v_7240);
  assign v_7240 = ~v_7224;
  assign v_7241 = v_7242 & 1'h1;
  assign v_7242 = v_7243 & v_7244;
  assign v_7243 = ~act_7223;
  assign v_7244 = v_7245 | v_7249;
  assign v_7245 = v_7246 | v_7247;
  assign v_7246 = mux_7246(v_7180);
  assign v_7247 = mux_7247(v_7248);
  assign v_7248 = ~v_7180;
  assign v_7249 = ~v_7220;
  assign v_7250 = v_7251 | v_7252;
  assign v_7251 = mux_7251(v_7222);
  assign v_7252 = mux_7252(v_7241);
  assign v_7253 = v_7254 & 1'h1;
  assign v_7254 = v_7255 & v_7256;
  assign v_7255 = ~act_7179;
  assign v_7256 = v_7257 | v_7261;
  assign v_7257 = v_7258 | v_7259;
  assign v_7258 = mux_7258(v_7080);
  assign v_7259 = mux_7259(v_7260);
  assign v_7260 = ~v_7080;
  assign v_7261 = ~v_7176;
  assign v_7262 = v_7263 | v_7264;
  assign v_7263 = mux_7263(v_7178);
  assign v_7264 = mux_7264(v_7253);
  assign v_7265 = v_7266 & 1'h1;
  assign v_7266 = v_7267 & v_7268;
  assign v_7267 = ~act_7079;
  assign v_7268 = v_7269 | v_7277;
  assign v_7269 = v_7270 | v_7275;
  assign v_7270 = mux_7270(v_7271);
  assign v_7271 = v_7076 & v_7272;
  assign v_7272 = v_7273 & 1'h1;
  assign v_7273 = v_7274 | 1'h0;
  assign v_7274 = ~v_7069;
  assign v_7275 = mux_7275(v_7276);
  assign v_7276 = ~v_7271;
  assign v_7277 = ~v_7076;
  assign v_7278 = v_7279 | v_7280;
  assign v_7279 = mux_7279(v_7078);
  assign v_7280 = mux_7280(v_7265);
  assign v_7282 = v_7283 | v_7470;
  assign v_7283 = act_7284 & 1'h1;
  assign act_7284 = v_7285 | v_7371;
  assign v_7285 = v_7286 & v_7372;
  assign v_7286 = v_7287 & v_7381;
  assign v_7287 = ~v_7288;
  assign v_7289 = v_7290 | v_7365;
  assign v_7290 = act_7291 & 1'h1;
  assign act_7291 = v_7292 | v_7322;
  assign v_7292 = v_7293 & v_7323;
  assign v_7293 = v_7294 & v_7332;
  assign v_7294 = ~v_7295;
  assign v_7296 = v_7297 | v_7316;
  assign v_7297 = act_7298 & 1'h1;
  assign act_7298 = v_7299 | v_7305;
  assign v_7299 = v_7300 & v_7306;
  assign v_7300 = v_7301 & vout_canPeek_7311;
  assign v_7301 = ~vout_canPeek_7302;
  pebbles_core
    pebbles_core_7302
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7303),
       .in0_consume_en(vin0_consume_en_7302),
       .out_canPeek(vout_canPeek_7302),
       .out_peek(vout_peek_7302));
  assign v_7303 = v_7304 | v_7309;
  assign v_7304 = mux_7304(v_7305);
  assign v_7305 = vout_canPeek_7302 & v_7306;
  assign v_7306 = v_7307 & 1'h1;
  assign v_7307 = v_7308 | 1'h0;
  assign v_7308 = ~v_7295;
  assign v_7309 = mux_7309(v_7310);
  assign v_7310 = ~v_7305;
  pebbles_core
    pebbles_core_7311
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7312),
       .in0_consume_en(vin0_consume_en_7311),
       .out_canPeek(vout_canPeek_7311),
       .out_peek(vout_peek_7311));
  assign v_7312 = v_7313 | v_7314;
  assign v_7313 = mux_7313(v_7299);
  assign v_7314 = mux_7314(v_7315);
  assign v_7315 = ~v_7299;
  assign v_7316 = v_7317 & 1'h1;
  assign v_7317 = v_7318 & v_7319;
  assign v_7318 = ~act_7298;
  assign v_7319 = v_7320 | v_7328;
  assign v_7320 = v_7321 | v_7326;
  assign v_7321 = mux_7321(v_7322);
  assign v_7322 = v_7295 & v_7323;
  assign v_7323 = v_7324 & 1'h1;
  assign v_7324 = v_7325 | 1'h0;
  assign v_7325 = ~v_7288;
  assign v_7326 = mux_7326(v_7327);
  assign v_7327 = ~v_7322;
  assign v_7328 = ~v_7295;
  assign v_7329 = v_7330 | v_7331;
  assign v_7330 = mux_7330(v_7297);
  assign v_7331 = mux_7331(v_7316);
  assign v_7333 = v_7334 | v_7353;
  assign v_7334 = act_7335 & 1'h1;
  assign act_7335 = v_7336 | v_7342;
  assign v_7336 = v_7337 & v_7343;
  assign v_7337 = v_7338 & vout_canPeek_7348;
  assign v_7338 = ~vout_canPeek_7339;
  pebbles_core
    pebbles_core_7339
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7340),
       .in0_consume_en(vin0_consume_en_7339),
       .out_canPeek(vout_canPeek_7339),
       .out_peek(vout_peek_7339));
  assign v_7340 = v_7341 | v_7346;
  assign v_7341 = mux_7341(v_7342);
  assign v_7342 = vout_canPeek_7339 & v_7343;
  assign v_7343 = v_7344 & 1'h1;
  assign v_7344 = v_7345 | 1'h0;
  assign v_7345 = ~v_7332;
  assign v_7346 = mux_7346(v_7347);
  assign v_7347 = ~v_7342;
  pebbles_core
    pebbles_core_7348
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7349),
       .in0_consume_en(vin0_consume_en_7348),
       .out_canPeek(vout_canPeek_7348),
       .out_peek(vout_peek_7348));
  assign v_7349 = v_7350 | v_7351;
  assign v_7350 = mux_7350(v_7336);
  assign v_7351 = mux_7351(v_7352);
  assign v_7352 = ~v_7336;
  assign v_7353 = v_7354 & 1'h1;
  assign v_7354 = v_7355 & v_7356;
  assign v_7355 = ~act_7335;
  assign v_7356 = v_7357 | v_7361;
  assign v_7357 = v_7358 | v_7359;
  assign v_7358 = mux_7358(v_7292);
  assign v_7359 = mux_7359(v_7360);
  assign v_7360 = ~v_7292;
  assign v_7361 = ~v_7332;
  assign v_7362 = v_7363 | v_7364;
  assign v_7363 = mux_7363(v_7334);
  assign v_7364 = mux_7364(v_7353);
  assign v_7365 = v_7366 & 1'h1;
  assign v_7366 = v_7367 & v_7368;
  assign v_7367 = ~act_7291;
  assign v_7368 = v_7369 | v_7377;
  assign v_7369 = v_7370 | v_7375;
  assign v_7370 = mux_7370(v_7371);
  assign v_7371 = v_7288 & v_7372;
  assign v_7372 = v_7373 & 1'h1;
  assign v_7373 = v_7374 | 1'h0;
  assign v_7374 = ~v_7281;
  assign v_7375 = mux_7375(v_7376);
  assign v_7376 = ~v_7371;
  assign v_7377 = ~v_7288;
  assign v_7378 = v_7379 | v_7380;
  assign v_7379 = mux_7379(v_7290);
  assign v_7380 = mux_7380(v_7365);
  assign v_7382 = v_7383 | v_7458;
  assign v_7383 = act_7384 & 1'h1;
  assign act_7384 = v_7385 | v_7415;
  assign v_7385 = v_7386 & v_7416;
  assign v_7386 = v_7387 & v_7425;
  assign v_7387 = ~v_7388;
  assign v_7389 = v_7390 | v_7409;
  assign v_7390 = act_7391 & 1'h1;
  assign act_7391 = v_7392 | v_7398;
  assign v_7392 = v_7393 & v_7399;
  assign v_7393 = v_7394 & vout_canPeek_7404;
  assign v_7394 = ~vout_canPeek_7395;
  pebbles_core
    pebbles_core_7395
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7396),
       .in0_consume_en(vin0_consume_en_7395),
       .out_canPeek(vout_canPeek_7395),
       .out_peek(vout_peek_7395));
  assign v_7396 = v_7397 | v_7402;
  assign v_7397 = mux_7397(v_7398);
  assign v_7398 = vout_canPeek_7395 & v_7399;
  assign v_7399 = v_7400 & 1'h1;
  assign v_7400 = v_7401 | 1'h0;
  assign v_7401 = ~v_7388;
  assign v_7402 = mux_7402(v_7403);
  assign v_7403 = ~v_7398;
  pebbles_core
    pebbles_core_7404
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7405),
       .in0_consume_en(vin0_consume_en_7404),
       .out_canPeek(vout_canPeek_7404),
       .out_peek(vout_peek_7404));
  assign v_7405 = v_7406 | v_7407;
  assign v_7406 = mux_7406(v_7392);
  assign v_7407 = mux_7407(v_7408);
  assign v_7408 = ~v_7392;
  assign v_7409 = v_7410 & 1'h1;
  assign v_7410 = v_7411 & v_7412;
  assign v_7411 = ~act_7391;
  assign v_7412 = v_7413 | v_7421;
  assign v_7413 = v_7414 | v_7419;
  assign v_7414 = mux_7414(v_7415);
  assign v_7415 = v_7388 & v_7416;
  assign v_7416 = v_7417 & 1'h1;
  assign v_7417 = v_7418 | 1'h0;
  assign v_7418 = ~v_7381;
  assign v_7419 = mux_7419(v_7420);
  assign v_7420 = ~v_7415;
  assign v_7421 = ~v_7388;
  assign v_7422 = v_7423 | v_7424;
  assign v_7423 = mux_7423(v_7390);
  assign v_7424 = mux_7424(v_7409);
  assign v_7426 = v_7427 | v_7446;
  assign v_7427 = act_7428 & 1'h1;
  assign act_7428 = v_7429 | v_7435;
  assign v_7429 = v_7430 & v_7436;
  assign v_7430 = v_7431 & vout_canPeek_7441;
  assign v_7431 = ~vout_canPeek_7432;
  pebbles_core
    pebbles_core_7432
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7433),
       .in0_consume_en(vin0_consume_en_7432),
       .out_canPeek(vout_canPeek_7432),
       .out_peek(vout_peek_7432));
  assign v_7433 = v_7434 | v_7439;
  assign v_7434 = mux_7434(v_7435);
  assign v_7435 = vout_canPeek_7432 & v_7436;
  assign v_7436 = v_7437 & 1'h1;
  assign v_7437 = v_7438 | 1'h0;
  assign v_7438 = ~v_7425;
  assign v_7439 = mux_7439(v_7440);
  assign v_7440 = ~v_7435;
  pebbles_core
    pebbles_core_7441
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7442),
       .in0_consume_en(vin0_consume_en_7441),
       .out_canPeek(vout_canPeek_7441),
       .out_peek(vout_peek_7441));
  assign v_7442 = v_7443 | v_7444;
  assign v_7443 = mux_7443(v_7429);
  assign v_7444 = mux_7444(v_7445);
  assign v_7445 = ~v_7429;
  assign v_7446 = v_7447 & 1'h1;
  assign v_7447 = v_7448 & v_7449;
  assign v_7448 = ~act_7428;
  assign v_7449 = v_7450 | v_7454;
  assign v_7450 = v_7451 | v_7452;
  assign v_7451 = mux_7451(v_7385);
  assign v_7452 = mux_7452(v_7453);
  assign v_7453 = ~v_7385;
  assign v_7454 = ~v_7425;
  assign v_7455 = v_7456 | v_7457;
  assign v_7456 = mux_7456(v_7427);
  assign v_7457 = mux_7457(v_7446);
  assign v_7458 = v_7459 & 1'h1;
  assign v_7459 = v_7460 & v_7461;
  assign v_7460 = ~act_7384;
  assign v_7461 = v_7462 | v_7466;
  assign v_7462 = v_7463 | v_7464;
  assign v_7463 = mux_7463(v_7285);
  assign v_7464 = mux_7464(v_7465);
  assign v_7465 = ~v_7285;
  assign v_7466 = ~v_7381;
  assign v_7467 = v_7468 | v_7469;
  assign v_7468 = mux_7468(v_7383);
  assign v_7469 = mux_7469(v_7458);
  assign v_7470 = v_7471 & 1'h1;
  assign v_7471 = v_7472 & v_7473;
  assign v_7472 = ~act_7284;
  assign v_7473 = v_7474 | v_7478;
  assign v_7474 = v_7475 | v_7476;
  assign v_7475 = mux_7475(v_7073);
  assign v_7476 = mux_7476(v_7477);
  assign v_7477 = ~v_7073;
  assign v_7478 = ~v_7281;
  assign v_7479 = v_7480 | v_7481;
  assign v_7480 = mux_7480(v_7283);
  assign v_7481 = mux_7481(v_7470);
  assign v_7482 = v_7483 & 1'h1;
  assign v_7483 = v_7484 & v_7485;
  assign v_7484 = ~act_7072;
  assign v_7485 = v_7486 | v_7494;
  assign v_7486 = v_7487 | v_7492;
  assign v_7487 = mux_7487(v_7488);
  assign v_7488 = v_7069 & v_7489;
  assign v_7489 = v_7490 & 1'h1;
  assign v_7490 = v_7491 | 1'h0;
  assign v_7491 = ~v_7062;
  assign v_7492 = mux_7492(v_7493);
  assign v_7493 = ~v_7488;
  assign v_7494 = ~v_7069;
  assign v_7495 = v_7496 | v_7497;
  assign v_7496 = mux_7496(v_7071);
  assign v_7497 = mux_7497(v_7482);
  assign v_7499 = v_7500 | v_7911;
  assign v_7500 = act_7501 & 1'h1;
  assign act_7501 = v_7502 | v_7700;
  assign v_7502 = v_7503 & v_7701;
  assign v_7503 = v_7504 & v_7710;
  assign v_7504 = ~v_7505;
  assign v_7506 = v_7507 | v_7694;
  assign v_7507 = act_7508 & 1'h1;
  assign act_7508 = v_7509 | v_7595;
  assign v_7509 = v_7510 & v_7596;
  assign v_7510 = v_7511 & v_7605;
  assign v_7511 = ~v_7512;
  assign v_7513 = v_7514 | v_7589;
  assign v_7514 = act_7515 & 1'h1;
  assign act_7515 = v_7516 | v_7546;
  assign v_7516 = v_7517 & v_7547;
  assign v_7517 = v_7518 & v_7556;
  assign v_7518 = ~v_7519;
  assign v_7520 = v_7521 | v_7540;
  assign v_7521 = act_7522 & 1'h1;
  assign act_7522 = v_7523 | v_7529;
  assign v_7523 = v_7524 & v_7530;
  assign v_7524 = v_7525 & vout_canPeek_7535;
  assign v_7525 = ~vout_canPeek_7526;
  pebbles_core
    pebbles_core_7526
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7527),
       .in0_consume_en(vin0_consume_en_7526),
       .out_canPeek(vout_canPeek_7526),
       .out_peek(vout_peek_7526));
  assign v_7527 = v_7528 | v_7533;
  assign v_7528 = mux_7528(v_7529);
  assign v_7529 = vout_canPeek_7526 & v_7530;
  assign v_7530 = v_7531 & 1'h1;
  assign v_7531 = v_7532 | 1'h0;
  assign v_7532 = ~v_7519;
  assign v_7533 = mux_7533(v_7534);
  assign v_7534 = ~v_7529;
  pebbles_core
    pebbles_core_7535
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7536),
       .in0_consume_en(vin0_consume_en_7535),
       .out_canPeek(vout_canPeek_7535),
       .out_peek(vout_peek_7535));
  assign v_7536 = v_7537 | v_7538;
  assign v_7537 = mux_7537(v_7523);
  assign v_7538 = mux_7538(v_7539);
  assign v_7539 = ~v_7523;
  assign v_7540 = v_7541 & 1'h1;
  assign v_7541 = v_7542 & v_7543;
  assign v_7542 = ~act_7522;
  assign v_7543 = v_7544 | v_7552;
  assign v_7544 = v_7545 | v_7550;
  assign v_7545 = mux_7545(v_7546);
  assign v_7546 = v_7519 & v_7547;
  assign v_7547 = v_7548 & 1'h1;
  assign v_7548 = v_7549 | 1'h0;
  assign v_7549 = ~v_7512;
  assign v_7550 = mux_7550(v_7551);
  assign v_7551 = ~v_7546;
  assign v_7552 = ~v_7519;
  assign v_7553 = v_7554 | v_7555;
  assign v_7554 = mux_7554(v_7521);
  assign v_7555 = mux_7555(v_7540);
  assign v_7557 = v_7558 | v_7577;
  assign v_7558 = act_7559 & 1'h1;
  assign act_7559 = v_7560 | v_7566;
  assign v_7560 = v_7561 & v_7567;
  assign v_7561 = v_7562 & vout_canPeek_7572;
  assign v_7562 = ~vout_canPeek_7563;
  pebbles_core
    pebbles_core_7563
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7564),
       .in0_consume_en(vin0_consume_en_7563),
       .out_canPeek(vout_canPeek_7563),
       .out_peek(vout_peek_7563));
  assign v_7564 = v_7565 | v_7570;
  assign v_7565 = mux_7565(v_7566);
  assign v_7566 = vout_canPeek_7563 & v_7567;
  assign v_7567 = v_7568 & 1'h1;
  assign v_7568 = v_7569 | 1'h0;
  assign v_7569 = ~v_7556;
  assign v_7570 = mux_7570(v_7571);
  assign v_7571 = ~v_7566;
  pebbles_core
    pebbles_core_7572
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7573),
       .in0_consume_en(vin0_consume_en_7572),
       .out_canPeek(vout_canPeek_7572),
       .out_peek(vout_peek_7572));
  assign v_7573 = v_7574 | v_7575;
  assign v_7574 = mux_7574(v_7560);
  assign v_7575 = mux_7575(v_7576);
  assign v_7576 = ~v_7560;
  assign v_7577 = v_7578 & 1'h1;
  assign v_7578 = v_7579 & v_7580;
  assign v_7579 = ~act_7559;
  assign v_7580 = v_7581 | v_7585;
  assign v_7581 = v_7582 | v_7583;
  assign v_7582 = mux_7582(v_7516);
  assign v_7583 = mux_7583(v_7584);
  assign v_7584 = ~v_7516;
  assign v_7585 = ~v_7556;
  assign v_7586 = v_7587 | v_7588;
  assign v_7587 = mux_7587(v_7558);
  assign v_7588 = mux_7588(v_7577);
  assign v_7589 = v_7590 & 1'h1;
  assign v_7590 = v_7591 & v_7592;
  assign v_7591 = ~act_7515;
  assign v_7592 = v_7593 | v_7601;
  assign v_7593 = v_7594 | v_7599;
  assign v_7594 = mux_7594(v_7595);
  assign v_7595 = v_7512 & v_7596;
  assign v_7596 = v_7597 & 1'h1;
  assign v_7597 = v_7598 | 1'h0;
  assign v_7598 = ~v_7505;
  assign v_7599 = mux_7599(v_7600);
  assign v_7600 = ~v_7595;
  assign v_7601 = ~v_7512;
  assign v_7602 = v_7603 | v_7604;
  assign v_7603 = mux_7603(v_7514);
  assign v_7604 = mux_7604(v_7589);
  assign v_7606 = v_7607 | v_7682;
  assign v_7607 = act_7608 & 1'h1;
  assign act_7608 = v_7609 | v_7639;
  assign v_7609 = v_7610 & v_7640;
  assign v_7610 = v_7611 & v_7649;
  assign v_7611 = ~v_7612;
  assign v_7613 = v_7614 | v_7633;
  assign v_7614 = act_7615 & 1'h1;
  assign act_7615 = v_7616 | v_7622;
  assign v_7616 = v_7617 & v_7623;
  assign v_7617 = v_7618 & vout_canPeek_7628;
  assign v_7618 = ~vout_canPeek_7619;
  pebbles_core
    pebbles_core_7619
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7620),
       .in0_consume_en(vin0_consume_en_7619),
       .out_canPeek(vout_canPeek_7619),
       .out_peek(vout_peek_7619));
  assign v_7620 = v_7621 | v_7626;
  assign v_7621 = mux_7621(v_7622);
  assign v_7622 = vout_canPeek_7619 & v_7623;
  assign v_7623 = v_7624 & 1'h1;
  assign v_7624 = v_7625 | 1'h0;
  assign v_7625 = ~v_7612;
  assign v_7626 = mux_7626(v_7627);
  assign v_7627 = ~v_7622;
  pebbles_core
    pebbles_core_7628
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7629),
       .in0_consume_en(vin0_consume_en_7628),
       .out_canPeek(vout_canPeek_7628),
       .out_peek(vout_peek_7628));
  assign v_7629 = v_7630 | v_7631;
  assign v_7630 = mux_7630(v_7616);
  assign v_7631 = mux_7631(v_7632);
  assign v_7632 = ~v_7616;
  assign v_7633 = v_7634 & 1'h1;
  assign v_7634 = v_7635 & v_7636;
  assign v_7635 = ~act_7615;
  assign v_7636 = v_7637 | v_7645;
  assign v_7637 = v_7638 | v_7643;
  assign v_7638 = mux_7638(v_7639);
  assign v_7639 = v_7612 & v_7640;
  assign v_7640 = v_7641 & 1'h1;
  assign v_7641 = v_7642 | 1'h0;
  assign v_7642 = ~v_7605;
  assign v_7643 = mux_7643(v_7644);
  assign v_7644 = ~v_7639;
  assign v_7645 = ~v_7612;
  assign v_7646 = v_7647 | v_7648;
  assign v_7647 = mux_7647(v_7614);
  assign v_7648 = mux_7648(v_7633);
  assign v_7650 = v_7651 | v_7670;
  assign v_7651 = act_7652 & 1'h1;
  assign act_7652 = v_7653 | v_7659;
  assign v_7653 = v_7654 & v_7660;
  assign v_7654 = v_7655 & vout_canPeek_7665;
  assign v_7655 = ~vout_canPeek_7656;
  pebbles_core
    pebbles_core_7656
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7657),
       .in0_consume_en(vin0_consume_en_7656),
       .out_canPeek(vout_canPeek_7656),
       .out_peek(vout_peek_7656));
  assign v_7657 = v_7658 | v_7663;
  assign v_7658 = mux_7658(v_7659);
  assign v_7659 = vout_canPeek_7656 & v_7660;
  assign v_7660 = v_7661 & 1'h1;
  assign v_7661 = v_7662 | 1'h0;
  assign v_7662 = ~v_7649;
  assign v_7663 = mux_7663(v_7664);
  assign v_7664 = ~v_7659;
  pebbles_core
    pebbles_core_7665
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7666),
       .in0_consume_en(vin0_consume_en_7665),
       .out_canPeek(vout_canPeek_7665),
       .out_peek(vout_peek_7665));
  assign v_7666 = v_7667 | v_7668;
  assign v_7667 = mux_7667(v_7653);
  assign v_7668 = mux_7668(v_7669);
  assign v_7669 = ~v_7653;
  assign v_7670 = v_7671 & 1'h1;
  assign v_7671 = v_7672 & v_7673;
  assign v_7672 = ~act_7652;
  assign v_7673 = v_7674 | v_7678;
  assign v_7674 = v_7675 | v_7676;
  assign v_7675 = mux_7675(v_7609);
  assign v_7676 = mux_7676(v_7677);
  assign v_7677 = ~v_7609;
  assign v_7678 = ~v_7649;
  assign v_7679 = v_7680 | v_7681;
  assign v_7680 = mux_7680(v_7651);
  assign v_7681 = mux_7681(v_7670);
  assign v_7682 = v_7683 & 1'h1;
  assign v_7683 = v_7684 & v_7685;
  assign v_7684 = ~act_7608;
  assign v_7685 = v_7686 | v_7690;
  assign v_7686 = v_7687 | v_7688;
  assign v_7687 = mux_7687(v_7509);
  assign v_7688 = mux_7688(v_7689);
  assign v_7689 = ~v_7509;
  assign v_7690 = ~v_7605;
  assign v_7691 = v_7692 | v_7693;
  assign v_7692 = mux_7692(v_7607);
  assign v_7693 = mux_7693(v_7682);
  assign v_7694 = v_7695 & 1'h1;
  assign v_7695 = v_7696 & v_7697;
  assign v_7696 = ~act_7508;
  assign v_7697 = v_7698 | v_7706;
  assign v_7698 = v_7699 | v_7704;
  assign v_7699 = mux_7699(v_7700);
  assign v_7700 = v_7505 & v_7701;
  assign v_7701 = v_7702 & 1'h1;
  assign v_7702 = v_7703 | 1'h0;
  assign v_7703 = ~v_7498;
  assign v_7704 = mux_7704(v_7705);
  assign v_7705 = ~v_7700;
  assign v_7706 = ~v_7505;
  assign v_7707 = v_7708 | v_7709;
  assign v_7708 = mux_7708(v_7507);
  assign v_7709 = mux_7709(v_7694);
  assign v_7711 = v_7712 | v_7899;
  assign v_7712 = act_7713 & 1'h1;
  assign act_7713 = v_7714 | v_7800;
  assign v_7714 = v_7715 & v_7801;
  assign v_7715 = v_7716 & v_7810;
  assign v_7716 = ~v_7717;
  assign v_7718 = v_7719 | v_7794;
  assign v_7719 = act_7720 & 1'h1;
  assign act_7720 = v_7721 | v_7751;
  assign v_7721 = v_7722 & v_7752;
  assign v_7722 = v_7723 & v_7761;
  assign v_7723 = ~v_7724;
  assign v_7725 = v_7726 | v_7745;
  assign v_7726 = act_7727 & 1'h1;
  assign act_7727 = v_7728 | v_7734;
  assign v_7728 = v_7729 & v_7735;
  assign v_7729 = v_7730 & vout_canPeek_7740;
  assign v_7730 = ~vout_canPeek_7731;
  pebbles_core
    pebbles_core_7731
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7732),
       .in0_consume_en(vin0_consume_en_7731),
       .out_canPeek(vout_canPeek_7731),
       .out_peek(vout_peek_7731));
  assign v_7732 = v_7733 | v_7738;
  assign v_7733 = mux_7733(v_7734);
  assign v_7734 = vout_canPeek_7731 & v_7735;
  assign v_7735 = v_7736 & 1'h1;
  assign v_7736 = v_7737 | 1'h0;
  assign v_7737 = ~v_7724;
  assign v_7738 = mux_7738(v_7739);
  assign v_7739 = ~v_7734;
  pebbles_core
    pebbles_core_7740
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7741),
       .in0_consume_en(vin0_consume_en_7740),
       .out_canPeek(vout_canPeek_7740),
       .out_peek(vout_peek_7740));
  assign v_7741 = v_7742 | v_7743;
  assign v_7742 = mux_7742(v_7728);
  assign v_7743 = mux_7743(v_7744);
  assign v_7744 = ~v_7728;
  assign v_7745 = v_7746 & 1'h1;
  assign v_7746 = v_7747 & v_7748;
  assign v_7747 = ~act_7727;
  assign v_7748 = v_7749 | v_7757;
  assign v_7749 = v_7750 | v_7755;
  assign v_7750 = mux_7750(v_7751);
  assign v_7751 = v_7724 & v_7752;
  assign v_7752 = v_7753 & 1'h1;
  assign v_7753 = v_7754 | 1'h0;
  assign v_7754 = ~v_7717;
  assign v_7755 = mux_7755(v_7756);
  assign v_7756 = ~v_7751;
  assign v_7757 = ~v_7724;
  assign v_7758 = v_7759 | v_7760;
  assign v_7759 = mux_7759(v_7726);
  assign v_7760 = mux_7760(v_7745);
  assign v_7762 = v_7763 | v_7782;
  assign v_7763 = act_7764 & 1'h1;
  assign act_7764 = v_7765 | v_7771;
  assign v_7765 = v_7766 & v_7772;
  assign v_7766 = v_7767 & vout_canPeek_7777;
  assign v_7767 = ~vout_canPeek_7768;
  pebbles_core
    pebbles_core_7768
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7769),
       .in0_consume_en(vin0_consume_en_7768),
       .out_canPeek(vout_canPeek_7768),
       .out_peek(vout_peek_7768));
  assign v_7769 = v_7770 | v_7775;
  assign v_7770 = mux_7770(v_7771);
  assign v_7771 = vout_canPeek_7768 & v_7772;
  assign v_7772 = v_7773 & 1'h1;
  assign v_7773 = v_7774 | 1'h0;
  assign v_7774 = ~v_7761;
  assign v_7775 = mux_7775(v_7776);
  assign v_7776 = ~v_7771;
  pebbles_core
    pebbles_core_7777
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7778),
       .in0_consume_en(vin0_consume_en_7777),
       .out_canPeek(vout_canPeek_7777),
       .out_peek(vout_peek_7777));
  assign v_7778 = v_7779 | v_7780;
  assign v_7779 = mux_7779(v_7765);
  assign v_7780 = mux_7780(v_7781);
  assign v_7781 = ~v_7765;
  assign v_7782 = v_7783 & 1'h1;
  assign v_7783 = v_7784 & v_7785;
  assign v_7784 = ~act_7764;
  assign v_7785 = v_7786 | v_7790;
  assign v_7786 = v_7787 | v_7788;
  assign v_7787 = mux_7787(v_7721);
  assign v_7788 = mux_7788(v_7789);
  assign v_7789 = ~v_7721;
  assign v_7790 = ~v_7761;
  assign v_7791 = v_7792 | v_7793;
  assign v_7792 = mux_7792(v_7763);
  assign v_7793 = mux_7793(v_7782);
  assign v_7794 = v_7795 & 1'h1;
  assign v_7795 = v_7796 & v_7797;
  assign v_7796 = ~act_7720;
  assign v_7797 = v_7798 | v_7806;
  assign v_7798 = v_7799 | v_7804;
  assign v_7799 = mux_7799(v_7800);
  assign v_7800 = v_7717 & v_7801;
  assign v_7801 = v_7802 & 1'h1;
  assign v_7802 = v_7803 | 1'h0;
  assign v_7803 = ~v_7710;
  assign v_7804 = mux_7804(v_7805);
  assign v_7805 = ~v_7800;
  assign v_7806 = ~v_7717;
  assign v_7807 = v_7808 | v_7809;
  assign v_7808 = mux_7808(v_7719);
  assign v_7809 = mux_7809(v_7794);
  assign v_7811 = v_7812 | v_7887;
  assign v_7812 = act_7813 & 1'h1;
  assign act_7813 = v_7814 | v_7844;
  assign v_7814 = v_7815 & v_7845;
  assign v_7815 = v_7816 & v_7854;
  assign v_7816 = ~v_7817;
  assign v_7818 = v_7819 | v_7838;
  assign v_7819 = act_7820 & 1'h1;
  assign act_7820 = v_7821 | v_7827;
  assign v_7821 = v_7822 & v_7828;
  assign v_7822 = v_7823 & vout_canPeek_7833;
  assign v_7823 = ~vout_canPeek_7824;
  pebbles_core
    pebbles_core_7824
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7825),
       .in0_consume_en(vin0_consume_en_7824),
       .out_canPeek(vout_canPeek_7824),
       .out_peek(vout_peek_7824));
  assign v_7825 = v_7826 | v_7831;
  assign v_7826 = mux_7826(v_7827);
  assign v_7827 = vout_canPeek_7824 & v_7828;
  assign v_7828 = v_7829 & 1'h1;
  assign v_7829 = v_7830 | 1'h0;
  assign v_7830 = ~v_7817;
  assign v_7831 = mux_7831(v_7832);
  assign v_7832 = ~v_7827;
  pebbles_core
    pebbles_core_7833
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7834),
       .in0_consume_en(vin0_consume_en_7833),
       .out_canPeek(vout_canPeek_7833),
       .out_peek(vout_peek_7833));
  assign v_7834 = v_7835 | v_7836;
  assign v_7835 = mux_7835(v_7821);
  assign v_7836 = mux_7836(v_7837);
  assign v_7837 = ~v_7821;
  assign v_7838 = v_7839 & 1'h1;
  assign v_7839 = v_7840 & v_7841;
  assign v_7840 = ~act_7820;
  assign v_7841 = v_7842 | v_7850;
  assign v_7842 = v_7843 | v_7848;
  assign v_7843 = mux_7843(v_7844);
  assign v_7844 = v_7817 & v_7845;
  assign v_7845 = v_7846 & 1'h1;
  assign v_7846 = v_7847 | 1'h0;
  assign v_7847 = ~v_7810;
  assign v_7848 = mux_7848(v_7849);
  assign v_7849 = ~v_7844;
  assign v_7850 = ~v_7817;
  assign v_7851 = v_7852 | v_7853;
  assign v_7852 = mux_7852(v_7819);
  assign v_7853 = mux_7853(v_7838);
  assign v_7855 = v_7856 | v_7875;
  assign v_7856 = act_7857 & 1'h1;
  assign act_7857 = v_7858 | v_7864;
  assign v_7858 = v_7859 & v_7865;
  assign v_7859 = v_7860 & vout_canPeek_7870;
  assign v_7860 = ~vout_canPeek_7861;
  pebbles_core
    pebbles_core_7861
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7862),
       .in0_consume_en(vin0_consume_en_7861),
       .out_canPeek(vout_canPeek_7861),
       .out_peek(vout_peek_7861));
  assign v_7862 = v_7863 | v_7868;
  assign v_7863 = mux_7863(v_7864);
  assign v_7864 = vout_canPeek_7861 & v_7865;
  assign v_7865 = v_7866 & 1'h1;
  assign v_7866 = v_7867 | 1'h0;
  assign v_7867 = ~v_7854;
  assign v_7868 = mux_7868(v_7869);
  assign v_7869 = ~v_7864;
  pebbles_core
    pebbles_core_7870
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_7871),
       .in0_consume_en(vin0_consume_en_7870),
       .out_canPeek(vout_canPeek_7870),
       .out_peek(vout_peek_7870));
  assign v_7871 = v_7872 | v_7873;
  assign v_7872 = mux_7872(v_7858);
  assign v_7873 = mux_7873(v_7874);
  assign v_7874 = ~v_7858;
  assign v_7875 = v_7876 & 1'h1;
  assign v_7876 = v_7877 & v_7878;
  assign v_7877 = ~act_7857;
  assign v_7878 = v_7879 | v_7883;
  assign v_7879 = v_7880 | v_7881;
  assign v_7880 = mux_7880(v_7814);
  assign v_7881 = mux_7881(v_7882);
  assign v_7882 = ~v_7814;
  assign v_7883 = ~v_7854;
  assign v_7884 = v_7885 | v_7886;
  assign v_7885 = mux_7885(v_7856);
  assign v_7886 = mux_7886(v_7875);
  assign v_7887 = v_7888 & 1'h1;
  assign v_7888 = v_7889 & v_7890;
  assign v_7889 = ~act_7813;
  assign v_7890 = v_7891 | v_7895;
  assign v_7891 = v_7892 | v_7893;
  assign v_7892 = mux_7892(v_7714);
  assign v_7893 = mux_7893(v_7894);
  assign v_7894 = ~v_7714;
  assign v_7895 = ~v_7810;
  assign v_7896 = v_7897 | v_7898;
  assign v_7897 = mux_7897(v_7812);
  assign v_7898 = mux_7898(v_7887);
  assign v_7899 = v_7900 & 1'h1;
  assign v_7900 = v_7901 & v_7902;
  assign v_7901 = ~act_7713;
  assign v_7902 = v_7903 | v_7907;
  assign v_7903 = v_7904 | v_7905;
  assign v_7904 = mux_7904(v_7502);
  assign v_7905 = mux_7905(v_7906);
  assign v_7906 = ~v_7502;
  assign v_7907 = ~v_7710;
  assign v_7908 = v_7909 | v_7910;
  assign v_7909 = mux_7909(v_7712);
  assign v_7910 = mux_7910(v_7899);
  assign v_7911 = v_7912 & 1'h1;
  assign v_7912 = v_7913 & v_7914;
  assign v_7913 = ~act_7501;
  assign v_7914 = v_7915 | v_7919;
  assign v_7915 = v_7916 | v_7917;
  assign v_7916 = mux_7916(v_7066);
  assign v_7917 = mux_7917(v_7918);
  assign v_7918 = ~v_7066;
  assign v_7919 = ~v_7498;
  assign v_7920 = v_7921 | v_7922;
  assign v_7921 = mux_7921(v_7500);
  assign v_7922 = mux_7922(v_7911);
  assign v_7923 = v_7924 & 1'h1;
  assign v_7924 = v_7925 & v_7926;
  assign v_7925 = ~act_7065;
  assign v_7926 = v_7927 | v_7931;
  assign v_7927 = v_7928 | v_7929;
  assign v_7928 = mux_7928(v_6182);
  assign v_7929 = mux_7929(v_7930);
  assign v_7930 = ~v_6182;
  assign v_7931 = ~v_7062;
  assign v_7932 = v_7933 | v_7934;
  assign v_7933 = mux_7933(v_7064);
  assign v_7934 = mux_7934(v_7923);
  assign v_7935 = v_7936 & 1'h1;
  assign v_7936 = v_7937 & v_7938;
  assign v_7937 = ~act_6181;
  assign v_7938 = v_7939 | v_7943;
  assign v_7939 = v_7940 | v_7941;
  assign v_7940 = mux_7940(v_4402);
  assign v_7941 = mux_7941(v_7942);
  assign v_7942 = ~v_4402;
  assign v_7943 = ~v_6178;
  assign v_7944 = v_7945 | v_7946;
  assign v_7945 = mux_7945(v_6180);
  assign v_7946 = mux_7946(v_7935);
  assign v_7947 = v_7948 & 1'h1;
  assign v_7948 = v_7949 & v_7950;
  assign v_7949 = ~act_4401;
  assign v_7950 = v_7951 | v_22313;
  assign v_7951 = v_7952 | v_22311;
  assign v_7952 = mux_7952(v_7953);
  assign v_7953 = v_4398 & v_7954;
  assign v_7954 = v_7955 & 1'h1;
  assign v_7955 = v_7956 | 1'h0;
  assign v_7956 = ~v_7957;
  assign v_7958 = v_7959 | v_7961;
  assign v_7959 = act_7960 & 1'h1;
  assign act_7960 = v_4395 | v_7953;
  assign v_7961 = v_7962 & 1'h1;
  assign v_7962 = v_7963 & v_7964;
  assign v_7963 = ~act_7960;
  assign v_7964 = v_7965 | v_22307;
  assign v_7965 = v_7966 | v_22305;
  assign v_7966 = mux_7966(v_7967);
  assign v_7967 = v_7957 & v_7968;
  assign v_7968 = v_7969 & 1'h1;
  assign v_7969 = v_7970 | 1'h0;
  assign v_7970 = ~v_7971;
  assign v_7972 = v_7973 | v_22291;
  assign v_7973 = act_7974 & 1'h1;
  assign act_7974 = v_7975 | v_7967;
  assign v_7975 = v_7976 & v_7968;
  assign v_7976 = v_7977 & v_7978;
  assign v_7977 = ~v_7957;
  assign v_7979 = v_7980 | v_22279;
  assign v_7980 = act_7981 & 1'h1;
  assign act_7981 = v_7982 | v_15124;
  assign v_7982 = v_7983 & v_15125;
  assign v_7983 = v_7984 & v_15134;
  assign v_7984 = ~v_7985;
  assign v_7986 = v_7987 | v_15118;
  assign v_7987 = act_7988 & 1'h1;
  assign act_7988 = v_7989 | v_11547;
  assign v_7989 = v_7990 & v_11548;
  assign v_7990 = v_7991 & v_11557;
  assign v_7991 = ~v_7992;
  assign v_7993 = v_7994 | v_11541;
  assign v_7994 = act_7995 & 1'h1;
  assign act_7995 = v_7996 | v_9762;
  assign v_7996 = v_7997 & v_9763;
  assign v_7997 = v_7998 & v_9772;
  assign v_7998 = ~v_7999;
  assign v_8000 = v_8001 | v_9756;
  assign v_8001 = act_8002 & 1'h1;
  assign act_8002 = v_8003 | v_8873;
  assign v_8003 = v_8004 & v_8874;
  assign v_8004 = v_8005 & v_8883;
  assign v_8005 = ~v_8006;
  assign v_8007 = v_8008 | v_8867;
  assign v_8008 = act_8009 & 1'h1;
  assign act_8009 = v_8010 | v_8432;
  assign v_8010 = v_8011 & v_8433;
  assign v_8011 = v_8012 & v_8442;
  assign v_8012 = ~v_8013;
  assign v_8014 = v_8015 | v_8426;
  assign v_8015 = act_8016 & 1'h1;
  assign act_8016 = v_8017 | v_8215;
  assign v_8017 = v_8018 & v_8216;
  assign v_8018 = v_8019 & v_8225;
  assign v_8019 = ~v_8020;
  assign v_8021 = v_8022 | v_8209;
  assign v_8022 = act_8023 & 1'h1;
  assign act_8023 = v_8024 | v_8110;
  assign v_8024 = v_8025 & v_8111;
  assign v_8025 = v_8026 & v_8120;
  assign v_8026 = ~v_8027;
  assign v_8028 = v_8029 | v_8104;
  assign v_8029 = act_8030 & 1'h1;
  assign act_8030 = v_8031 | v_8061;
  assign v_8031 = v_8032 & v_8062;
  assign v_8032 = v_8033 & v_8071;
  assign v_8033 = ~v_8034;
  assign v_8035 = v_8036 | v_8055;
  assign v_8036 = act_8037 & 1'h1;
  assign act_8037 = v_8038 | v_8044;
  assign v_8038 = v_8039 & v_8045;
  assign v_8039 = v_8040 & vout_canPeek_8050;
  assign v_8040 = ~vout_canPeek_8041;
  pebbles_core
    pebbles_core_8041
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8042),
       .in0_consume_en(vin0_consume_en_8041),
       .out_canPeek(vout_canPeek_8041),
       .out_peek(vout_peek_8041));
  assign v_8042 = v_8043 | v_8048;
  assign v_8043 = mux_8043(v_8044);
  assign v_8044 = vout_canPeek_8041 & v_8045;
  assign v_8045 = v_8046 & 1'h1;
  assign v_8046 = v_8047 | 1'h0;
  assign v_8047 = ~v_8034;
  assign v_8048 = mux_8048(v_8049);
  assign v_8049 = ~v_8044;
  pebbles_core
    pebbles_core_8050
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8051),
       .in0_consume_en(vin0_consume_en_8050),
       .out_canPeek(vout_canPeek_8050),
       .out_peek(vout_peek_8050));
  assign v_8051 = v_8052 | v_8053;
  assign v_8052 = mux_8052(v_8038);
  assign v_8053 = mux_8053(v_8054);
  assign v_8054 = ~v_8038;
  assign v_8055 = v_8056 & 1'h1;
  assign v_8056 = v_8057 & v_8058;
  assign v_8057 = ~act_8037;
  assign v_8058 = v_8059 | v_8067;
  assign v_8059 = v_8060 | v_8065;
  assign v_8060 = mux_8060(v_8061);
  assign v_8061 = v_8034 & v_8062;
  assign v_8062 = v_8063 & 1'h1;
  assign v_8063 = v_8064 | 1'h0;
  assign v_8064 = ~v_8027;
  assign v_8065 = mux_8065(v_8066);
  assign v_8066 = ~v_8061;
  assign v_8067 = ~v_8034;
  assign v_8068 = v_8069 | v_8070;
  assign v_8069 = mux_8069(v_8036);
  assign v_8070 = mux_8070(v_8055);
  assign v_8072 = v_8073 | v_8092;
  assign v_8073 = act_8074 & 1'h1;
  assign act_8074 = v_8075 | v_8081;
  assign v_8075 = v_8076 & v_8082;
  assign v_8076 = v_8077 & vout_canPeek_8087;
  assign v_8077 = ~vout_canPeek_8078;
  pebbles_core
    pebbles_core_8078
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8079),
       .in0_consume_en(vin0_consume_en_8078),
       .out_canPeek(vout_canPeek_8078),
       .out_peek(vout_peek_8078));
  assign v_8079 = v_8080 | v_8085;
  assign v_8080 = mux_8080(v_8081);
  assign v_8081 = vout_canPeek_8078 & v_8082;
  assign v_8082 = v_8083 & 1'h1;
  assign v_8083 = v_8084 | 1'h0;
  assign v_8084 = ~v_8071;
  assign v_8085 = mux_8085(v_8086);
  assign v_8086 = ~v_8081;
  pebbles_core
    pebbles_core_8087
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8088),
       .in0_consume_en(vin0_consume_en_8087),
       .out_canPeek(vout_canPeek_8087),
       .out_peek(vout_peek_8087));
  assign v_8088 = v_8089 | v_8090;
  assign v_8089 = mux_8089(v_8075);
  assign v_8090 = mux_8090(v_8091);
  assign v_8091 = ~v_8075;
  assign v_8092 = v_8093 & 1'h1;
  assign v_8093 = v_8094 & v_8095;
  assign v_8094 = ~act_8074;
  assign v_8095 = v_8096 | v_8100;
  assign v_8096 = v_8097 | v_8098;
  assign v_8097 = mux_8097(v_8031);
  assign v_8098 = mux_8098(v_8099);
  assign v_8099 = ~v_8031;
  assign v_8100 = ~v_8071;
  assign v_8101 = v_8102 | v_8103;
  assign v_8102 = mux_8102(v_8073);
  assign v_8103 = mux_8103(v_8092);
  assign v_8104 = v_8105 & 1'h1;
  assign v_8105 = v_8106 & v_8107;
  assign v_8106 = ~act_8030;
  assign v_8107 = v_8108 | v_8116;
  assign v_8108 = v_8109 | v_8114;
  assign v_8109 = mux_8109(v_8110);
  assign v_8110 = v_8027 & v_8111;
  assign v_8111 = v_8112 & 1'h1;
  assign v_8112 = v_8113 | 1'h0;
  assign v_8113 = ~v_8020;
  assign v_8114 = mux_8114(v_8115);
  assign v_8115 = ~v_8110;
  assign v_8116 = ~v_8027;
  assign v_8117 = v_8118 | v_8119;
  assign v_8118 = mux_8118(v_8029);
  assign v_8119 = mux_8119(v_8104);
  assign v_8121 = v_8122 | v_8197;
  assign v_8122 = act_8123 & 1'h1;
  assign act_8123 = v_8124 | v_8154;
  assign v_8124 = v_8125 & v_8155;
  assign v_8125 = v_8126 & v_8164;
  assign v_8126 = ~v_8127;
  assign v_8128 = v_8129 | v_8148;
  assign v_8129 = act_8130 & 1'h1;
  assign act_8130 = v_8131 | v_8137;
  assign v_8131 = v_8132 & v_8138;
  assign v_8132 = v_8133 & vout_canPeek_8143;
  assign v_8133 = ~vout_canPeek_8134;
  pebbles_core
    pebbles_core_8134
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8135),
       .in0_consume_en(vin0_consume_en_8134),
       .out_canPeek(vout_canPeek_8134),
       .out_peek(vout_peek_8134));
  assign v_8135 = v_8136 | v_8141;
  assign v_8136 = mux_8136(v_8137);
  assign v_8137 = vout_canPeek_8134 & v_8138;
  assign v_8138 = v_8139 & 1'h1;
  assign v_8139 = v_8140 | 1'h0;
  assign v_8140 = ~v_8127;
  assign v_8141 = mux_8141(v_8142);
  assign v_8142 = ~v_8137;
  pebbles_core
    pebbles_core_8143
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8144),
       .in0_consume_en(vin0_consume_en_8143),
       .out_canPeek(vout_canPeek_8143),
       .out_peek(vout_peek_8143));
  assign v_8144 = v_8145 | v_8146;
  assign v_8145 = mux_8145(v_8131);
  assign v_8146 = mux_8146(v_8147);
  assign v_8147 = ~v_8131;
  assign v_8148 = v_8149 & 1'h1;
  assign v_8149 = v_8150 & v_8151;
  assign v_8150 = ~act_8130;
  assign v_8151 = v_8152 | v_8160;
  assign v_8152 = v_8153 | v_8158;
  assign v_8153 = mux_8153(v_8154);
  assign v_8154 = v_8127 & v_8155;
  assign v_8155 = v_8156 & 1'h1;
  assign v_8156 = v_8157 | 1'h0;
  assign v_8157 = ~v_8120;
  assign v_8158 = mux_8158(v_8159);
  assign v_8159 = ~v_8154;
  assign v_8160 = ~v_8127;
  assign v_8161 = v_8162 | v_8163;
  assign v_8162 = mux_8162(v_8129);
  assign v_8163 = mux_8163(v_8148);
  assign v_8165 = v_8166 | v_8185;
  assign v_8166 = act_8167 & 1'h1;
  assign act_8167 = v_8168 | v_8174;
  assign v_8168 = v_8169 & v_8175;
  assign v_8169 = v_8170 & vout_canPeek_8180;
  assign v_8170 = ~vout_canPeek_8171;
  pebbles_core
    pebbles_core_8171
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8172),
       .in0_consume_en(vin0_consume_en_8171),
       .out_canPeek(vout_canPeek_8171),
       .out_peek(vout_peek_8171));
  assign v_8172 = v_8173 | v_8178;
  assign v_8173 = mux_8173(v_8174);
  assign v_8174 = vout_canPeek_8171 & v_8175;
  assign v_8175 = v_8176 & 1'h1;
  assign v_8176 = v_8177 | 1'h0;
  assign v_8177 = ~v_8164;
  assign v_8178 = mux_8178(v_8179);
  assign v_8179 = ~v_8174;
  pebbles_core
    pebbles_core_8180
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8181),
       .in0_consume_en(vin0_consume_en_8180),
       .out_canPeek(vout_canPeek_8180),
       .out_peek(vout_peek_8180));
  assign v_8181 = v_8182 | v_8183;
  assign v_8182 = mux_8182(v_8168);
  assign v_8183 = mux_8183(v_8184);
  assign v_8184 = ~v_8168;
  assign v_8185 = v_8186 & 1'h1;
  assign v_8186 = v_8187 & v_8188;
  assign v_8187 = ~act_8167;
  assign v_8188 = v_8189 | v_8193;
  assign v_8189 = v_8190 | v_8191;
  assign v_8190 = mux_8190(v_8124);
  assign v_8191 = mux_8191(v_8192);
  assign v_8192 = ~v_8124;
  assign v_8193 = ~v_8164;
  assign v_8194 = v_8195 | v_8196;
  assign v_8195 = mux_8195(v_8166);
  assign v_8196 = mux_8196(v_8185);
  assign v_8197 = v_8198 & 1'h1;
  assign v_8198 = v_8199 & v_8200;
  assign v_8199 = ~act_8123;
  assign v_8200 = v_8201 | v_8205;
  assign v_8201 = v_8202 | v_8203;
  assign v_8202 = mux_8202(v_8024);
  assign v_8203 = mux_8203(v_8204);
  assign v_8204 = ~v_8024;
  assign v_8205 = ~v_8120;
  assign v_8206 = v_8207 | v_8208;
  assign v_8207 = mux_8207(v_8122);
  assign v_8208 = mux_8208(v_8197);
  assign v_8209 = v_8210 & 1'h1;
  assign v_8210 = v_8211 & v_8212;
  assign v_8211 = ~act_8023;
  assign v_8212 = v_8213 | v_8221;
  assign v_8213 = v_8214 | v_8219;
  assign v_8214 = mux_8214(v_8215);
  assign v_8215 = v_8020 & v_8216;
  assign v_8216 = v_8217 & 1'h1;
  assign v_8217 = v_8218 | 1'h0;
  assign v_8218 = ~v_8013;
  assign v_8219 = mux_8219(v_8220);
  assign v_8220 = ~v_8215;
  assign v_8221 = ~v_8020;
  assign v_8222 = v_8223 | v_8224;
  assign v_8223 = mux_8223(v_8022);
  assign v_8224 = mux_8224(v_8209);
  assign v_8226 = v_8227 | v_8414;
  assign v_8227 = act_8228 & 1'h1;
  assign act_8228 = v_8229 | v_8315;
  assign v_8229 = v_8230 & v_8316;
  assign v_8230 = v_8231 & v_8325;
  assign v_8231 = ~v_8232;
  assign v_8233 = v_8234 | v_8309;
  assign v_8234 = act_8235 & 1'h1;
  assign act_8235 = v_8236 | v_8266;
  assign v_8236 = v_8237 & v_8267;
  assign v_8237 = v_8238 & v_8276;
  assign v_8238 = ~v_8239;
  assign v_8240 = v_8241 | v_8260;
  assign v_8241 = act_8242 & 1'h1;
  assign act_8242 = v_8243 | v_8249;
  assign v_8243 = v_8244 & v_8250;
  assign v_8244 = v_8245 & vout_canPeek_8255;
  assign v_8245 = ~vout_canPeek_8246;
  pebbles_core
    pebbles_core_8246
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8247),
       .in0_consume_en(vin0_consume_en_8246),
       .out_canPeek(vout_canPeek_8246),
       .out_peek(vout_peek_8246));
  assign v_8247 = v_8248 | v_8253;
  assign v_8248 = mux_8248(v_8249);
  assign v_8249 = vout_canPeek_8246 & v_8250;
  assign v_8250 = v_8251 & 1'h1;
  assign v_8251 = v_8252 | 1'h0;
  assign v_8252 = ~v_8239;
  assign v_8253 = mux_8253(v_8254);
  assign v_8254 = ~v_8249;
  pebbles_core
    pebbles_core_8255
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8256),
       .in0_consume_en(vin0_consume_en_8255),
       .out_canPeek(vout_canPeek_8255),
       .out_peek(vout_peek_8255));
  assign v_8256 = v_8257 | v_8258;
  assign v_8257 = mux_8257(v_8243);
  assign v_8258 = mux_8258(v_8259);
  assign v_8259 = ~v_8243;
  assign v_8260 = v_8261 & 1'h1;
  assign v_8261 = v_8262 & v_8263;
  assign v_8262 = ~act_8242;
  assign v_8263 = v_8264 | v_8272;
  assign v_8264 = v_8265 | v_8270;
  assign v_8265 = mux_8265(v_8266);
  assign v_8266 = v_8239 & v_8267;
  assign v_8267 = v_8268 & 1'h1;
  assign v_8268 = v_8269 | 1'h0;
  assign v_8269 = ~v_8232;
  assign v_8270 = mux_8270(v_8271);
  assign v_8271 = ~v_8266;
  assign v_8272 = ~v_8239;
  assign v_8273 = v_8274 | v_8275;
  assign v_8274 = mux_8274(v_8241);
  assign v_8275 = mux_8275(v_8260);
  assign v_8277 = v_8278 | v_8297;
  assign v_8278 = act_8279 & 1'h1;
  assign act_8279 = v_8280 | v_8286;
  assign v_8280 = v_8281 & v_8287;
  assign v_8281 = v_8282 & vout_canPeek_8292;
  assign v_8282 = ~vout_canPeek_8283;
  pebbles_core
    pebbles_core_8283
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8284),
       .in0_consume_en(vin0_consume_en_8283),
       .out_canPeek(vout_canPeek_8283),
       .out_peek(vout_peek_8283));
  assign v_8284 = v_8285 | v_8290;
  assign v_8285 = mux_8285(v_8286);
  assign v_8286 = vout_canPeek_8283 & v_8287;
  assign v_8287 = v_8288 & 1'h1;
  assign v_8288 = v_8289 | 1'h0;
  assign v_8289 = ~v_8276;
  assign v_8290 = mux_8290(v_8291);
  assign v_8291 = ~v_8286;
  pebbles_core
    pebbles_core_8292
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8293),
       .in0_consume_en(vin0_consume_en_8292),
       .out_canPeek(vout_canPeek_8292),
       .out_peek(vout_peek_8292));
  assign v_8293 = v_8294 | v_8295;
  assign v_8294 = mux_8294(v_8280);
  assign v_8295 = mux_8295(v_8296);
  assign v_8296 = ~v_8280;
  assign v_8297 = v_8298 & 1'h1;
  assign v_8298 = v_8299 & v_8300;
  assign v_8299 = ~act_8279;
  assign v_8300 = v_8301 | v_8305;
  assign v_8301 = v_8302 | v_8303;
  assign v_8302 = mux_8302(v_8236);
  assign v_8303 = mux_8303(v_8304);
  assign v_8304 = ~v_8236;
  assign v_8305 = ~v_8276;
  assign v_8306 = v_8307 | v_8308;
  assign v_8307 = mux_8307(v_8278);
  assign v_8308 = mux_8308(v_8297);
  assign v_8309 = v_8310 & 1'h1;
  assign v_8310 = v_8311 & v_8312;
  assign v_8311 = ~act_8235;
  assign v_8312 = v_8313 | v_8321;
  assign v_8313 = v_8314 | v_8319;
  assign v_8314 = mux_8314(v_8315);
  assign v_8315 = v_8232 & v_8316;
  assign v_8316 = v_8317 & 1'h1;
  assign v_8317 = v_8318 | 1'h0;
  assign v_8318 = ~v_8225;
  assign v_8319 = mux_8319(v_8320);
  assign v_8320 = ~v_8315;
  assign v_8321 = ~v_8232;
  assign v_8322 = v_8323 | v_8324;
  assign v_8323 = mux_8323(v_8234);
  assign v_8324 = mux_8324(v_8309);
  assign v_8326 = v_8327 | v_8402;
  assign v_8327 = act_8328 & 1'h1;
  assign act_8328 = v_8329 | v_8359;
  assign v_8329 = v_8330 & v_8360;
  assign v_8330 = v_8331 & v_8369;
  assign v_8331 = ~v_8332;
  assign v_8333 = v_8334 | v_8353;
  assign v_8334 = act_8335 & 1'h1;
  assign act_8335 = v_8336 | v_8342;
  assign v_8336 = v_8337 & v_8343;
  assign v_8337 = v_8338 & vout_canPeek_8348;
  assign v_8338 = ~vout_canPeek_8339;
  pebbles_core
    pebbles_core_8339
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8340),
       .in0_consume_en(vin0_consume_en_8339),
       .out_canPeek(vout_canPeek_8339),
       .out_peek(vout_peek_8339));
  assign v_8340 = v_8341 | v_8346;
  assign v_8341 = mux_8341(v_8342);
  assign v_8342 = vout_canPeek_8339 & v_8343;
  assign v_8343 = v_8344 & 1'h1;
  assign v_8344 = v_8345 | 1'h0;
  assign v_8345 = ~v_8332;
  assign v_8346 = mux_8346(v_8347);
  assign v_8347 = ~v_8342;
  pebbles_core
    pebbles_core_8348
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8349),
       .in0_consume_en(vin0_consume_en_8348),
       .out_canPeek(vout_canPeek_8348),
       .out_peek(vout_peek_8348));
  assign v_8349 = v_8350 | v_8351;
  assign v_8350 = mux_8350(v_8336);
  assign v_8351 = mux_8351(v_8352);
  assign v_8352 = ~v_8336;
  assign v_8353 = v_8354 & 1'h1;
  assign v_8354 = v_8355 & v_8356;
  assign v_8355 = ~act_8335;
  assign v_8356 = v_8357 | v_8365;
  assign v_8357 = v_8358 | v_8363;
  assign v_8358 = mux_8358(v_8359);
  assign v_8359 = v_8332 & v_8360;
  assign v_8360 = v_8361 & 1'h1;
  assign v_8361 = v_8362 | 1'h0;
  assign v_8362 = ~v_8325;
  assign v_8363 = mux_8363(v_8364);
  assign v_8364 = ~v_8359;
  assign v_8365 = ~v_8332;
  assign v_8366 = v_8367 | v_8368;
  assign v_8367 = mux_8367(v_8334);
  assign v_8368 = mux_8368(v_8353);
  assign v_8370 = v_8371 | v_8390;
  assign v_8371 = act_8372 & 1'h1;
  assign act_8372 = v_8373 | v_8379;
  assign v_8373 = v_8374 & v_8380;
  assign v_8374 = v_8375 & vout_canPeek_8385;
  assign v_8375 = ~vout_canPeek_8376;
  pebbles_core
    pebbles_core_8376
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8377),
       .in0_consume_en(vin0_consume_en_8376),
       .out_canPeek(vout_canPeek_8376),
       .out_peek(vout_peek_8376));
  assign v_8377 = v_8378 | v_8383;
  assign v_8378 = mux_8378(v_8379);
  assign v_8379 = vout_canPeek_8376 & v_8380;
  assign v_8380 = v_8381 & 1'h1;
  assign v_8381 = v_8382 | 1'h0;
  assign v_8382 = ~v_8369;
  assign v_8383 = mux_8383(v_8384);
  assign v_8384 = ~v_8379;
  pebbles_core
    pebbles_core_8385
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8386),
       .in0_consume_en(vin0_consume_en_8385),
       .out_canPeek(vout_canPeek_8385),
       .out_peek(vout_peek_8385));
  assign v_8386 = v_8387 | v_8388;
  assign v_8387 = mux_8387(v_8373);
  assign v_8388 = mux_8388(v_8389);
  assign v_8389 = ~v_8373;
  assign v_8390 = v_8391 & 1'h1;
  assign v_8391 = v_8392 & v_8393;
  assign v_8392 = ~act_8372;
  assign v_8393 = v_8394 | v_8398;
  assign v_8394 = v_8395 | v_8396;
  assign v_8395 = mux_8395(v_8329);
  assign v_8396 = mux_8396(v_8397);
  assign v_8397 = ~v_8329;
  assign v_8398 = ~v_8369;
  assign v_8399 = v_8400 | v_8401;
  assign v_8400 = mux_8400(v_8371);
  assign v_8401 = mux_8401(v_8390);
  assign v_8402 = v_8403 & 1'h1;
  assign v_8403 = v_8404 & v_8405;
  assign v_8404 = ~act_8328;
  assign v_8405 = v_8406 | v_8410;
  assign v_8406 = v_8407 | v_8408;
  assign v_8407 = mux_8407(v_8229);
  assign v_8408 = mux_8408(v_8409);
  assign v_8409 = ~v_8229;
  assign v_8410 = ~v_8325;
  assign v_8411 = v_8412 | v_8413;
  assign v_8412 = mux_8412(v_8327);
  assign v_8413 = mux_8413(v_8402);
  assign v_8414 = v_8415 & 1'h1;
  assign v_8415 = v_8416 & v_8417;
  assign v_8416 = ~act_8228;
  assign v_8417 = v_8418 | v_8422;
  assign v_8418 = v_8419 | v_8420;
  assign v_8419 = mux_8419(v_8017);
  assign v_8420 = mux_8420(v_8421);
  assign v_8421 = ~v_8017;
  assign v_8422 = ~v_8225;
  assign v_8423 = v_8424 | v_8425;
  assign v_8424 = mux_8424(v_8227);
  assign v_8425 = mux_8425(v_8414);
  assign v_8426 = v_8427 & 1'h1;
  assign v_8427 = v_8428 & v_8429;
  assign v_8428 = ~act_8016;
  assign v_8429 = v_8430 | v_8438;
  assign v_8430 = v_8431 | v_8436;
  assign v_8431 = mux_8431(v_8432);
  assign v_8432 = v_8013 & v_8433;
  assign v_8433 = v_8434 & 1'h1;
  assign v_8434 = v_8435 | 1'h0;
  assign v_8435 = ~v_8006;
  assign v_8436 = mux_8436(v_8437);
  assign v_8437 = ~v_8432;
  assign v_8438 = ~v_8013;
  assign v_8439 = v_8440 | v_8441;
  assign v_8440 = mux_8440(v_8015);
  assign v_8441 = mux_8441(v_8426);
  assign v_8443 = v_8444 | v_8855;
  assign v_8444 = act_8445 & 1'h1;
  assign act_8445 = v_8446 | v_8644;
  assign v_8446 = v_8447 & v_8645;
  assign v_8447 = v_8448 & v_8654;
  assign v_8448 = ~v_8449;
  assign v_8450 = v_8451 | v_8638;
  assign v_8451 = act_8452 & 1'h1;
  assign act_8452 = v_8453 | v_8539;
  assign v_8453 = v_8454 & v_8540;
  assign v_8454 = v_8455 & v_8549;
  assign v_8455 = ~v_8456;
  assign v_8457 = v_8458 | v_8533;
  assign v_8458 = act_8459 & 1'h1;
  assign act_8459 = v_8460 | v_8490;
  assign v_8460 = v_8461 & v_8491;
  assign v_8461 = v_8462 & v_8500;
  assign v_8462 = ~v_8463;
  assign v_8464 = v_8465 | v_8484;
  assign v_8465 = act_8466 & 1'h1;
  assign act_8466 = v_8467 | v_8473;
  assign v_8467 = v_8468 & v_8474;
  assign v_8468 = v_8469 & vout_canPeek_8479;
  assign v_8469 = ~vout_canPeek_8470;
  pebbles_core
    pebbles_core_8470
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8471),
       .in0_consume_en(vin0_consume_en_8470),
       .out_canPeek(vout_canPeek_8470),
       .out_peek(vout_peek_8470));
  assign v_8471 = v_8472 | v_8477;
  assign v_8472 = mux_8472(v_8473);
  assign v_8473 = vout_canPeek_8470 & v_8474;
  assign v_8474 = v_8475 & 1'h1;
  assign v_8475 = v_8476 | 1'h0;
  assign v_8476 = ~v_8463;
  assign v_8477 = mux_8477(v_8478);
  assign v_8478 = ~v_8473;
  pebbles_core
    pebbles_core_8479
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8480),
       .in0_consume_en(vin0_consume_en_8479),
       .out_canPeek(vout_canPeek_8479),
       .out_peek(vout_peek_8479));
  assign v_8480 = v_8481 | v_8482;
  assign v_8481 = mux_8481(v_8467);
  assign v_8482 = mux_8482(v_8483);
  assign v_8483 = ~v_8467;
  assign v_8484 = v_8485 & 1'h1;
  assign v_8485 = v_8486 & v_8487;
  assign v_8486 = ~act_8466;
  assign v_8487 = v_8488 | v_8496;
  assign v_8488 = v_8489 | v_8494;
  assign v_8489 = mux_8489(v_8490);
  assign v_8490 = v_8463 & v_8491;
  assign v_8491 = v_8492 & 1'h1;
  assign v_8492 = v_8493 | 1'h0;
  assign v_8493 = ~v_8456;
  assign v_8494 = mux_8494(v_8495);
  assign v_8495 = ~v_8490;
  assign v_8496 = ~v_8463;
  assign v_8497 = v_8498 | v_8499;
  assign v_8498 = mux_8498(v_8465);
  assign v_8499 = mux_8499(v_8484);
  assign v_8501 = v_8502 | v_8521;
  assign v_8502 = act_8503 & 1'h1;
  assign act_8503 = v_8504 | v_8510;
  assign v_8504 = v_8505 & v_8511;
  assign v_8505 = v_8506 & vout_canPeek_8516;
  assign v_8506 = ~vout_canPeek_8507;
  pebbles_core
    pebbles_core_8507
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8508),
       .in0_consume_en(vin0_consume_en_8507),
       .out_canPeek(vout_canPeek_8507),
       .out_peek(vout_peek_8507));
  assign v_8508 = v_8509 | v_8514;
  assign v_8509 = mux_8509(v_8510);
  assign v_8510 = vout_canPeek_8507 & v_8511;
  assign v_8511 = v_8512 & 1'h1;
  assign v_8512 = v_8513 | 1'h0;
  assign v_8513 = ~v_8500;
  assign v_8514 = mux_8514(v_8515);
  assign v_8515 = ~v_8510;
  pebbles_core
    pebbles_core_8516
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8517),
       .in0_consume_en(vin0_consume_en_8516),
       .out_canPeek(vout_canPeek_8516),
       .out_peek(vout_peek_8516));
  assign v_8517 = v_8518 | v_8519;
  assign v_8518 = mux_8518(v_8504);
  assign v_8519 = mux_8519(v_8520);
  assign v_8520 = ~v_8504;
  assign v_8521 = v_8522 & 1'h1;
  assign v_8522 = v_8523 & v_8524;
  assign v_8523 = ~act_8503;
  assign v_8524 = v_8525 | v_8529;
  assign v_8525 = v_8526 | v_8527;
  assign v_8526 = mux_8526(v_8460);
  assign v_8527 = mux_8527(v_8528);
  assign v_8528 = ~v_8460;
  assign v_8529 = ~v_8500;
  assign v_8530 = v_8531 | v_8532;
  assign v_8531 = mux_8531(v_8502);
  assign v_8532 = mux_8532(v_8521);
  assign v_8533 = v_8534 & 1'h1;
  assign v_8534 = v_8535 & v_8536;
  assign v_8535 = ~act_8459;
  assign v_8536 = v_8537 | v_8545;
  assign v_8537 = v_8538 | v_8543;
  assign v_8538 = mux_8538(v_8539);
  assign v_8539 = v_8456 & v_8540;
  assign v_8540 = v_8541 & 1'h1;
  assign v_8541 = v_8542 | 1'h0;
  assign v_8542 = ~v_8449;
  assign v_8543 = mux_8543(v_8544);
  assign v_8544 = ~v_8539;
  assign v_8545 = ~v_8456;
  assign v_8546 = v_8547 | v_8548;
  assign v_8547 = mux_8547(v_8458);
  assign v_8548 = mux_8548(v_8533);
  assign v_8550 = v_8551 | v_8626;
  assign v_8551 = act_8552 & 1'h1;
  assign act_8552 = v_8553 | v_8583;
  assign v_8553 = v_8554 & v_8584;
  assign v_8554 = v_8555 & v_8593;
  assign v_8555 = ~v_8556;
  assign v_8557 = v_8558 | v_8577;
  assign v_8558 = act_8559 & 1'h1;
  assign act_8559 = v_8560 | v_8566;
  assign v_8560 = v_8561 & v_8567;
  assign v_8561 = v_8562 & vout_canPeek_8572;
  assign v_8562 = ~vout_canPeek_8563;
  pebbles_core
    pebbles_core_8563
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8564),
       .in0_consume_en(vin0_consume_en_8563),
       .out_canPeek(vout_canPeek_8563),
       .out_peek(vout_peek_8563));
  assign v_8564 = v_8565 | v_8570;
  assign v_8565 = mux_8565(v_8566);
  assign v_8566 = vout_canPeek_8563 & v_8567;
  assign v_8567 = v_8568 & 1'h1;
  assign v_8568 = v_8569 | 1'h0;
  assign v_8569 = ~v_8556;
  assign v_8570 = mux_8570(v_8571);
  assign v_8571 = ~v_8566;
  pebbles_core
    pebbles_core_8572
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8573),
       .in0_consume_en(vin0_consume_en_8572),
       .out_canPeek(vout_canPeek_8572),
       .out_peek(vout_peek_8572));
  assign v_8573 = v_8574 | v_8575;
  assign v_8574 = mux_8574(v_8560);
  assign v_8575 = mux_8575(v_8576);
  assign v_8576 = ~v_8560;
  assign v_8577 = v_8578 & 1'h1;
  assign v_8578 = v_8579 & v_8580;
  assign v_8579 = ~act_8559;
  assign v_8580 = v_8581 | v_8589;
  assign v_8581 = v_8582 | v_8587;
  assign v_8582 = mux_8582(v_8583);
  assign v_8583 = v_8556 & v_8584;
  assign v_8584 = v_8585 & 1'h1;
  assign v_8585 = v_8586 | 1'h0;
  assign v_8586 = ~v_8549;
  assign v_8587 = mux_8587(v_8588);
  assign v_8588 = ~v_8583;
  assign v_8589 = ~v_8556;
  assign v_8590 = v_8591 | v_8592;
  assign v_8591 = mux_8591(v_8558);
  assign v_8592 = mux_8592(v_8577);
  assign v_8594 = v_8595 | v_8614;
  assign v_8595 = act_8596 & 1'h1;
  assign act_8596 = v_8597 | v_8603;
  assign v_8597 = v_8598 & v_8604;
  assign v_8598 = v_8599 & vout_canPeek_8609;
  assign v_8599 = ~vout_canPeek_8600;
  pebbles_core
    pebbles_core_8600
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8601),
       .in0_consume_en(vin0_consume_en_8600),
       .out_canPeek(vout_canPeek_8600),
       .out_peek(vout_peek_8600));
  assign v_8601 = v_8602 | v_8607;
  assign v_8602 = mux_8602(v_8603);
  assign v_8603 = vout_canPeek_8600 & v_8604;
  assign v_8604 = v_8605 & 1'h1;
  assign v_8605 = v_8606 | 1'h0;
  assign v_8606 = ~v_8593;
  assign v_8607 = mux_8607(v_8608);
  assign v_8608 = ~v_8603;
  pebbles_core
    pebbles_core_8609
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8610),
       .in0_consume_en(vin0_consume_en_8609),
       .out_canPeek(vout_canPeek_8609),
       .out_peek(vout_peek_8609));
  assign v_8610 = v_8611 | v_8612;
  assign v_8611 = mux_8611(v_8597);
  assign v_8612 = mux_8612(v_8613);
  assign v_8613 = ~v_8597;
  assign v_8614 = v_8615 & 1'h1;
  assign v_8615 = v_8616 & v_8617;
  assign v_8616 = ~act_8596;
  assign v_8617 = v_8618 | v_8622;
  assign v_8618 = v_8619 | v_8620;
  assign v_8619 = mux_8619(v_8553);
  assign v_8620 = mux_8620(v_8621);
  assign v_8621 = ~v_8553;
  assign v_8622 = ~v_8593;
  assign v_8623 = v_8624 | v_8625;
  assign v_8624 = mux_8624(v_8595);
  assign v_8625 = mux_8625(v_8614);
  assign v_8626 = v_8627 & 1'h1;
  assign v_8627 = v_8628 & v_8629;
  assign v_8628 = ~act_8552;
  assign v_8629 = v_8630 | v_8634;
  assign v_8630 = v_8631 | v_8632;
  assign v_8631 = mux_8631(v_8453);
  assign v_8632 = mux_8632(v_8633);
  assign v_8633 = ~v_8453;
  assign v_8634 = ~v_8549;
  assign v_8635 = v_8636 | v_8637;
  assign v_8636 = mux_8636(v_8551);
  assign v_8637 = mux_8637(v_8626);
  assign v_8638 = v_8639 & 1'h1;
  assign v_8639 = v_8640 & v_8641;
  assign v_8640 = ~act_8452;
  assign v_8641 = v_8642 | v_8650;
  assign v_8642 = v_8643 | v_8648;
  assign v_8643 = mux_8643(v_8644);
  assign v_8644 = v_8449 & v_8645;
  assign v_8645 = v_8646 & 1'h1;
  assign v_8646 = v_8647 | 1'h0;
  assign v_8647 = ~v_8442;
  assign v_8648 = mux_8648(v_8649);
  assign v_8649 = ~v_8644;
  assign v_8650 = ~v_8449;
  assign v_8651 = v_8652 | v_8653;
  assign v_8652 = mux_8652(v_8451);
  assign v_8653 = mux_8653(v_8638);
  assign v_8655 = v_8656 | v_8843;
  assign v_8656 = act_8657 & 1'h1;
  assign act_8657 = v_8658 | v_8744;
  assign v_8658 = v_8659 & v_8745;
  assign v_8659 = v_8660 & v_8754;
  assign v_8660 = ~v_8661;
  assign v_8662 = v_8663 | v_8738;
  assign v_8663 = act_8664 & 1'h1;
  assign act_8664 = v_8665 | v_8695;
  assign v_8665 = v_8666 & v_8696;
  assign v_8666 = v_8667 & v_8705;
  assign v_8667 = ~v_8668;
  assign v_8669 = v_8670 | v_8689;
  assign v_8670 = act_8671 & 1'h1;
  assign act_8671 = v_8672 | v_8678;
  assign v_8672 = v_8673 & v_8679;
  assign v_8673 = v_8674 & vout_canPeek_8684;
  assign v_8674 = ~vout_canPeek_8675;
  pebbles_core
    pebbles_core_8675
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8676),
       .in0_consume_en(vin0_consume_en_8675),
       .out_canPeek(vout_canPeek_8675),
       .out_peek(vout_peek_8675));
  assign v_8676 = v_8677 | v_8682;
  assign v_8677 = mux_8677(v_8678);
  assign v_8678 = vout_canPeek_8675 & v_8679;
  assign v_8679 = v_8680 & 1'h1;
  assign v_8680 = v_8681 | 1'h0;
  assign v_8681 = ~v_8668;
  assign v_8682 = mux_8682(v_8683);
  assign v_8683 = ~v_8678;
  pebbles_core
    pebbles_core_8684
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8685),
       .in0_consume_en(vin0_consume_en_8684),
       .out_canPeek(vout_canPeek_8684),
       .out_peek(vout_peek_8684));
  assign v_8685 = v_8686 | v_8687;
  assign v_8686 = mux_8686(v_8672);
  assign v_8687 = mux_8687(v_8688);
  assign v_8688 = ~v_8672;
  assign v_8689 = v_8690 & 1'h1;
  assign v_8690 = v_8691 & v_8692;
  assign v_8691 = ~act_8671;
  assign v_8692 = v_8693 | v_8701;
  assign v_8693 = v_8694 | v_8699;
  assign v_8694 = mux_8694(v_8695);
  assign v_8695 = v_8668 & v_8696;
  assign v_8696 = v_8697 & 1'h1;
  assign v_8697 = v_8698 | 1'h0;
  assign v_8698 = ~v_8661;
  assign v_8699 = mux_8699(v_8700);
  assign v_8700 = ~v_8695;
  assign v_8701 = ~v_8668;
  assign v_8702 = v_8703 | v_8704;
  assign v_8703 = mux_8703(v_8670);
  assign v_8704 = mux_8704(v_8689);
  assign v_8706 = v_8707 | v_8726;
  assign v_8707 = act_8708 & 1'h1;
  assign act_8708 = v_8709 | v_8715;
  assign v_8709 = v_8710 & v_8716;
  assign v_8710 = v_8711 & vout_canPeek_8721;
  assign v_8711 = ~vout_canPeek_8712;
  pebbles_core
    pebbles_core_8712
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8713),
       .in0_consume_en(vin0_consume_en_8712),
       .out_canPeek(vout_canPeek_8712),
       .out_peek(vout_peek_8712));
  assign v_8713 = v_8714 | v_8719;
  assign v_8714 = mux_8714(v_8715);
  assign v_8715 = vout_canPeek_8712 & v_8716;
  assign v_8716 = v_8717 & 1'h1;
  assign v_8717 = v_8718 | 1'h0;
  assign v_8718 = ~v_8705;
  assign v_8719 = mux_8719(v_8720);
  assign v_8720 = ~v_8715;
  pebbles_core
    pebbles_core_8721
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8722),
       .in0_consume_en(vin0_consume_en_8721),
       .out_canPeek(vout_canPeek_8721),
       .out_peek(vout_peek_8721));
  assign v_8722 = v_8723 | v_8724;
  assign v_8723 = mux_8723(v_8709);
  assign v_8724 = mux_8724(v_8725);
  assign v_8725 = ~v_8709;
  assign v_8726 = v_8727 & 1'h1;
  assign v_8727 = v_8728 & v_8729;
  assign v_8728 = ~act_8708;
  assign v_8729 = v_8730 | v_8734;
  assign v_8730 = v_8731 | v_8732;
  assign v_8731 = mux_8731(v_8665);
  assign v_8732 = mux_8732(v_8733);
  assign v_8733 = ~v_8665;
  assign v_8734 = ~v_8705;
  assign v_8735 = v_8736 | v_8737;
  assign v_8736 = mux_8736(v_8707);
  assign v_8737 = mux_8737(v_8726);
  assign v_8738 = v_8739 & 1'h1;
  assign v_8739 = v_8740 & v_8741;
  assign v_8740 = ~act_8664;
  assign v_8741 = v_8742 | v_8750;
  assign v_8742 = v_8743 | v_8748;
  assign v_8743 = mux_8743(v_8744);
  assign v_8744 = v_8661 & v_8745;
  assign v_8745 = v_8746 & 1'h1;
  assign v_8746 = v_8747 | 1'h0;
  assign v_8747 = ~v_8654;
  assign v_8748 = mux_8748(v_8749);
  assign v_8749 = ~v_8744;
  assign v_8750 = ~v_8661;
  assign v_8751 = v_8752 | v_8753;
  assign v_8752 = mux_8752(v_8663);
  assign v_8753 = mux_8753(v_8738);
  assign v_8755 = v_8756 | v_8831;
  assign v_8756 = act_8757 & 1'h1;
  assign act_8757 = v_8758 | v_8788;
  assign v_8758 = v_8759 & v_8789;
  assign v_8759 = v_8760 & v_8798;
  assign v_8760 = ~v_8761;
  assign v_8762 = v_8763 | v_8782;
  assign v_8763 = act_8764 & 1'h1;
  assign act_8764 = v_8765 | v_8771;
  assign v_8765 = v_8766 & v_8772;
  assign v_8766 = v_8767 & vout_canPeek_8777;
  assign v_8767 = ~vout_canPeek_8768;
  pebbles_core
    pebbles_core_8768
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8769),
       .in0_consume_en(vin0_consume_en_8768),
       .out_canPeek(vout_canPeek_8768),
       .out_peek(vout_peek_8768));
  assign v_8769 = v_8770 | v_8775;
  assign v_8770 = mux_8770(v_8771);
  assign v_8771 = vout_canPeek_8768 & v_8772;
  assign v_8772 = v_8773 & 1'h1;
  assign v_8773 = v_8774 | 1'h0;
  assign v_8774 = ~v_8761;
  assign v_8775 = mux_8775(v_8776);
  assign v_8776 = ~v_8771;
  pebbles_core
    pebbles_core_8777
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8778),
       .in0_consume_en(vin0_consume_en_8777),
       .out_canPeek(vout_canPeek_8777),
       .out_peek(vout_peek_8777));
  assign v_8778 = v_8779 | v_8780;
  assign v_8779 = mux_8779(v_8765);
  assign v_8780 = mux_8780(v_8781);
  assign v_8781 = ~v_8765;
  assign v_8782 = v_8783 & 1'h1;
  assign v_8783 = v_8784 & v_8785;
  assign v_8784 = ~act_8764;
  assign v_8785 = v_8786 | v_8794;
  assign v_8786 = v_8787 | v_8792;
  assign v_8787 = mux_8787(v_8788);
  assign v_8788 = v_8761 & v_8789;
  assign v_8789 = v_8790 & 1'h1;
  assign v_8790 = v_8791 | 1'h0;
  assign v_8791 = ~v_8754;
  assign v_8792 = mux_8792(v_8793);
  assign v_8793 = ~v_8788;
  assign v_8794 = ~v_8761;
  assign v_8795 = v_8796 | v_8797;
  assign v_8796 = mux_8796(v_8763);
  assign v_8797 = mux_8797(v_8782);
  assign v_8799 = v_8800 | v_8819;
  assign v_8800 = act_8801 & 1'h1;
  assign act_8801 = v_8802 | v_8808;
  assign v_8802 = v_8803 & v_8809;
  assign v_8803 = v_8804 & vout_canPeek_8814;
  assign v_8804 = ~vout_canPeek_8805;
  pebbles_core
    pebbles_core_8805
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8806),
       .in0_consume_en(vin0_consume_en_8805),
       .out_canPeek(vout_canPeek_8805),
       .out_peek(vout_peek_8805));
  assign v_8806 = v_8807 | v_8812;
  assign v_8807 = mux_8807(v_8808);
  assign v_8808 = vout_canPeek_8805 & v_8809;
  assign v_8809 = v_8810 & 1'h1;
  assign v_8810 = v_8811 | 1'h0;
  assign v_8811 = ~v_8798;
  assign v_8812 = mux_8812(v_8813);
  assign v_8813 = ~v_8808;
  pebbles_core
    pebbles_core_8814
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8815),
       .in0_consume_en(vin0_consume_en_8814),
       .out_canPeek(vout_canPeek_8814),
       .out_peek(vout_peek_8814));
  assign v_8815 = v_8816 | v_8817;
  assign v_8816 = mux_8816(v_8802);
  assign v_8817 = mux_8817(v_8818);
  assign v_8818 = ~v_8802;
  assign v_8819 = v_8820 & 1'h1;
  assign v_8820 = v_8821 & v_8822;
  assign v_8821 = ~act_8801;
  assign v_8822 = v_8823 | v_8827;
  assign v_8823 = v_8824 | v_8825;
  assign v_8824 = mux_8824(v_8758);
  assign v_8825 = mux_8825(v_8826);
  assign v_8826 = ~v_8758;
  assign v_8827 = ~v_8798;
  assign v_8828 = v_8829 | v_8830;
  assign v_8829 = mux_8829(v_8800);
  assign v_8830 = mux_8830(v_8819);
  assign v_8831 = v_8832 & 1'h1;
  assign v_8832 = v_8833 & v_8834;
  assign v_8833 = ~act_8757;
  assign v_8834 = v_8835 | v_8839;
  assign v_8835 = v_8836 | v_8837;
  assign v_8836 = mux_8836(v_8658);
  assign v_8837 = mux_8837(v_8838);
  assign v_8838 = ~v_8658;
  assign v_8839 = ~v_8754;
  assign v_8840 = v_8841 | v_8842;
  assign v_8841 = mux_8841(v_8756);
  assign v_8842 = mux_8842(v_8831);
  assign v_8843 = v_8844 & 1'h1;
  assign v_8844 = v_8845 & v_8846;
  assign v_8845 = ~act_8657;
  assign v_8846 = v_8847 | v_8851;
  assign v_8847 = v_8848 | v_8849;
  assign v_8848 = mux_8848(v_8446);
  assign v_8849 = mux_8849(v_8850);
  assign v_8850 = ~v_8446;
  assign v_8851 = ~v_8654;
  assign v_8852 = v_8853 | v_8854;
  assign v_8853 = mux_8853(v_8656);
  assign v_8854 = mux_8854(v_8843);
  assign v_8855 = v_8856 & 1'h1;
  assign v_8856 = v_8857 & v_8858;
  assign v_8857 = ~act_8445;
  assign v_8858 = v_8859 | v_8863;
  assign v_8859 = v_8860 | v_8861;
  assign v_8860 = mux_8860(v_8010);
  assign v_8861 = mux_8861(v_8862);
  assign v_8862 = ~v_8010;
  assign v_8863 = ~v_8442;
  assign v_8864 = v_8865 | v_8866;
  assign v_8865 = mux_8865(v_8444);
  assign v_8866 = mux_8866(v_8855);
  assign v_8867 = v_8868 & 1'h1;
  assign v_8868 = v_8869 & v_8870;
  assign v_8869 = ~act_8009;
  assign v_8870 = v_8871 | v_8879;
  assign v_8871 = v_8872 | v_8877;
  assign v_8872 = mux_8872(v_8873);
  assign v_8873 = v_8006 & v_8874;
  assign v_8874 = v_8875 & 1'h1;
  assign v_8875 = v_8876 | 1'h0;
  assign v_8876 = ~v_7999;
  assign v_8877 = mux_8877(v_8878);
  assign v_8878 = ~v_8873;
  assign v_8879 = ~v_8006;
  assign v_8880 = v_8881 | v_8882;
  assign v_8881 = mux_8881(v_8008);
  assign v_8882 = mux_8882(v_8867);
  assign v_8884 = v_8885 | v_9744;
  assign v_8885 = act_8886 & 1'h1;
  assign act_8886 = v_8887 | v_9309;
  assign v_8887 = v_8888 & v_9310;
  assign v_8888 = v_8889 & v_9319;
  assign v_8889 = ~v_8890;
  assign v_8891 = v_8892 | v_9303;
  assign v_8892 = act_8893 & 1'h1;
  assign act_8893 = v_8894 | v_9092;
  assign v_8894 = v_8895 & v_9093;
  assign v_8895 = v_8896 & v_9102;
  assign v_8896 = ~v_8897;
  assign v_8898 = v_8899 | v_9086;
  assign v_8899 = act_8900 & 1'h1;
  assign act_8900 = v_8901 | v_8987;
  assign v_8901 = v_8902 & v_8988;
  assign v_8902 = v_8903 & v_8997;
  assign v_8903 = ~v_8904;
  assign v_8905 = v_8906 | v_8981;
  assign v_8906 = act_8907 & 1'h1;
  assign act_8907 = v_8908 | v_8938;
  assign v_8908 = v_8909 & v_8939;
  assign v_8909 = v_8910 & v_8948;
  assign v_8910 = ~v_8911;
  assign v_8912 = v_8913 | v_8932;
  assign v_8913 = act_8914 & 1'h1;
  assign act_8914 = v_8915 | v_8921;
  assign v_8915 = v_8916 & v_8922;
  assign v_8916 = v_8917 & vout_canPeek_8927;
  assign v_8917 = ~vout_canPeek_8918;
  pebbles_core
    pebbles_core_8918
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8919),
       .in0_consume_en(vin0_consume_en_8918),
       .out_canPeek(vout_canPeek_8918),
       .out_peek(vout_peek_8918));
  assign v_8919 = v_8920 | v_8925;
  assign v_8920 = mux_8920(v_8921);
  assign v_8921 = vout_canPeek_8918 & v_8922;
  assign v_8922 = v_8923 & 1'h1;
  assign v_8923 = v_8924 | 1'h0;
  assign v_8924 = ~v_8911;
  assign v_8925 = mux_8925(v_8926);
  assign v_8926 = ~v_8921;
  pebbles_core
    pebbles_core_8927
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8928),
       .in0_consume_en(vin0_consume_en_8927),
       .out_canPeek(vout_canPeek_8927),
       .out_peek(vout_peek_8927));
  assign v_8928 = v_8929 | v_8930;
  assign v_8929 = mux_8929(v_8915);
  assign v_8930 = mux_8930(v_8931);
  assign v_8931 = ~v_8915;
  assign v_8932 = v_8933 & 1'h1;
  assign v_8933 = v_8934 & v_8935;
  assign v_8934 = ~act_8914;
  assign v_8935 = v_8936 | v_8944;
  assign v_8936 = v_8937 | v_8942;
  assign v_8937 = mux_8937(v_8938);
  assign v_8938 = v_8911 & v_8939;
  assign v_8939 = v_8940 & 1'h1;
  assign v_8940 = v_8941 | 1'h0;
  assign v_8941 = ~v_8904;
  assign v_8942 = mux_8942(v_8943);
  assign v_8943 = ~v_8938;
  assign v_8944 = ~v_8911;
  assign v_8945 = v_8946 | v_8947;
  assign v_8946 = mux_8946(v_8913);
  assign v_8947 = mux_8947(v_8932);
  assign v_8949 = v_8950 | v_8969;
  assign v_8950 = act_8951 & 1'h1;
  assign act_8951 = v_8952 | v_8958;
  assign v_8952 = v_8953 & v_8959;
  assign v_8953 = v_8954 & vout_canPeek_8964;
  assign v_8954 = ~vout_canPeek_8955;
  pebbles_core
    pebbles_core_8955
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8956),
       .in0_consume_en(vin0_consume_en_8955),
       .out_canPeek(vout_canPeek_8955),
       .out_peek(vout_peek_8955));
  assign v_8956 = v_8957 | v_8962;
  assign v_8957 = mux_8957(v_8958);
  assign v_8958 = vout_canPeek_8955 & v_8959;
  assign v_8959 = v_8960 & 1'h1;
  assign v_8960 = v_8961 | 1'h0;
  assign v_8961 = ~v_8948;
  assign v_8962 = mux_8962(v_8963);
  assign v_8963 = ~v_8958;
  pebbles_core
    pebbles_core_8964
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_8965),
       .in0_consume_en(vin0_consume_en_8964),
       .out_canPeek(vout_canPeek_8964),
       .out_peek(vout_peek_8964));
  assign v_8965 = v_8966 | v_8967;
  assign v_8966 = mux_8966(v_8952);
  assign v_8967 = mux_8967(v_8968);
  assign v_8968 = ~v_8952;
  assign v_8969 = v_8970 & 1'h1;
  assign v_8970 = v_8971 & v_8972;
  assign v_8971 = ~act_8951;
  assign v_8972 = v_8973 | v_8977;
  assign v_8973 = v_8974 | v_8975;
  assign v_8974 = mux_8974(v_8908);
  assign v_8975 = mux_8975(v_8976);
  assign v_8976 = ~v_8908;
  assign v_8977 = ~v_8948;
  assign v_8978 = v_8979 | v_8980;
  assign v_8979 = mux_8979(v_8950);
  assign v_8980 = mux_8980(v_8969);
  assign v_8981 = v_8982 & 1'h1;
  assign v_8982 = v_8983 & v_8984;
  assign v_8983 = ~act_8907;
  assign v_8984 = v_8985 | v_8993;
  assign v_8985 = v_8986 | v_8991;
  assign v_8986 = mux_8986(v_8987);
  assign v_8987 = v_8904 & v_8988;
  assign v_8988 = v_8989 & 1'h1;
  assign v_8989 = v_8990 | 1'h0;
  assign v_8990 = ~v_8897;
  assign v_8991 = mux_8991(v_8992);
  assign v_8992 = ~v_8987;
  assign v_8993 = ~v_8904;
  assign v_8994 = v_8995 | v_8996;
  assign v_8995 = mux_8995(v_8906);
  assign v_8996 = mux_8996(v_8981);
  assign v_8998 = v_8999 | v_9074;
  assign v_8999 = act_9000 & 1'h1;
  assign act_9000 = v_9001 | v_9031;
  assign v_9001 = v_9002 & v_9032;
  assign v_9002 = v_9003 & v_9041;
  assign v_9003 = ~v_9004;
  assign v_9005 = v_9006 | v_9025;
  assign v_9006 = act_9007 & 1'h1;
  assign act_9007 = v_9008 | v_9014;
  assign v_9008 = v_9009 & v_9015;
  assign v_9009 = v_9010 & vout_canPeek_9020;
  assign v_9010 = ~vout_canPeek_9011;
  pebbles_core
    pebbles_core_9011
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9012),
       .in0_consume_en(vin0_consume_en_9011),
       .out_canPeek(vout_canPeek_9011),
       .out_peek(vout_peek_9011));
  assign v_9012 = v_9013 | v_9018;
  assign v_9013 = mux_9013(v_9014);
  assign v_9014 = vout_canPeek_9011 & v_9015;
  assign v_9015 = v_9016 & 1'h1;
  assign v_9016 = v_9017 | 1'h0;
  assign v_9017 = ~v_9004;
  assign v_9018 = mux_9018(v_9019);
  assign v_9019 = ~v_9014;
  pebbles_core
    pebbles_core_9020
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9021),
       .in0_consume_en(vin0_consume_en_9020),
       .out_canPeek(vout_canPeek_9020),
       .out_peek(vout_peek_9020));
  assign v_9021 = v_9022 | v_9023;
  assign v_9022 = mux_9022(v_9008);
  assign v_9023 = mux_9023(v_9024);
  assign v_9024 = ~v_9008;
  assign v_9025 = v_9026 & 1'h1;
  assign v_9026 = v_9027 & v_9028;
  assign v_9027 = ~act_9007;
  assign v_9028 = v_9029 | v_9037;
  assign v_9029 = v_9030 | v_9035;
  assign v_9030 = mux_9030(v_9031);
  assign v_9031 = v_9004 & v_9032;
  assign v_9032 = v_9033 & 1'h1;
  assign v_9033 = v_9034 | 1'h0;
  assign v_9034 = ~v_8997;
  assign v_9035 = mux_9035(v_9036);
  assign v_9036 = ~v_9031;
  assign v_9037 = ~v_9004;
  assign v_9038 = v_9039 | v_9040;
  assign v_9039 = mux_9039(v_9006);
  assign v_9040 = mux_9040(v_9025);
  assign v_9042 = v_9043 | v_9062;
  assign v_9043 = act_9044 & 1'h1;
  assign act_9044 = v_9045 | v_9051;
  assign v_9045 = v_9046 & v_9052;
  assign v_9046 = v_9047 & vout_canPeek_9057;
  assign v_9047 = ~vout_canPeek_9048;
  pebbles_core
    pebbles_core_9048
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9049),
       .in0_consume_en(vin0_consume_en_9048),
       .out_canPeek(vout_canPeek_9048),
       .out_peek(vout_peek_9048));
  assign v_9049 = v_9050 | v_9055;
  assign v_9050 = mux_9050(v_9051);
  assign v_9051 = vout_canPeek_9048 & v_9052;
  assign v_9052 = v_9053 & 1'h1;
  assign v_9053 = v_9054 | 1'h0;
  assign v_9054 = ~v_9041;
  assign v_9055 = mux_9055(v_9056);
  assign v_9056 = ~v_9051;
  pebbles_core
    pebbles_core_9057
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9058),
       .in0_consume_en(vin0_consume_en_9057),
       .out_canPeek(vout_canPeek_9057),
       .out_peek(vout_peek_9057));
  assign v_9058 = v_9059 | v_9060;
  assign v_9059 = mux_9059(v_9045);
  assign v_9060 = mux_9060(v_9061);
  assign v_9061 = ~v_9045;
  assign v_9062 = v_9063 & 1'h1;
  assign v_9063 = v_9064 & v_9065;
  assign v_9064 = ~act_9044;
  assign v_9065 = v_9066 | v_9070;
  assign v_9066 = v_9067 | v_9068;
  assign v_9067 = mux_9067(v_9001);
  assign v_9068 = mux_9068(v_9069);
  assign v_9069 = ~v_9001;
  assign v_9070 = ~v_9041;
  assign v_9071 = v_9072 | v_9073;
  assign v_9072 = mux_9072(v_9043);
  assign v_9073 = mux_9073(v_9062);
  assign v_9074 = v_9075 & 1'h1;
  assign v_9075 = v_9076 & v_9077;
  assign v_9076 = ~act_9000;
  assign v_9077 = v_9078 | v_9082;
  assign v_9078 = v_9079 | v_9080;
  assign v_9079 = mux_9079(v_8901);
  assign v_9080 = mux_9080(v_9081);
  assign v_9081 = ~v_8901;
  assign v_9082 = ~v_8997;
  assign v_9083 = v_9084 | v_9085;
  assign v_9084 = mux_9084(v_8999);
  assign v_9085 = mux_9085(v_9074);
  assign v_9086 = v_9087 & 1'h1;
  assign v_9087 = v_9088 & v_9089;
  assign v_9088 = ~act_8900;
  assign v_9089 = v_9090 | v_9098;
  assign v_9090 = v_9091 | v_9096;
  assign v_9091 = mux_9091(v_9092);
  assign v_9092 = v_8897 & v_9093;
  assign v_9093 = v_9094 & 1'h1;
  assign v_9094 = v_9095 | 1'h0;
  assign v_9095 = ~v_8890;
  assign v_9096 = mux_9096(v_9097);
  assign v_9097 = ~v_9092;
  assign v_9098 = ~v_8897;
  assign v_9099 = v_9100 | v_9101;
  assign v_9100 = mux_9100(v_8899);
  assign v_9101 = mux_9101(v_9086);
  assign v_9103 = v_9104 | v_9291;
  assign v_9104 = act_9105 & 1'h1;
  assign act_9105 = v_9106 | v_9192;
  assign v_9106 = v_9107 & v_9193;
  assign v_9107 = v_9108 & v_9202;
  assign v_9108 = ~v_9109;
  assign v_9110 = v_9111 | v_9186;
  assign v_9111 = act_9112 & 1'h1;
  assign act_9112 = v_9113 | v_9143;
  assign v_9113 = v_9114 & v_9144;
  assign v_9114 = v_9115 & v_9153;
  assign v_9115 = ~v_9116;
  assign v_9117 = v_9118 | v_9137;
  assign v_9118 = act_9119 & 1'h1;
  assign act_9119 = v_9120 | v_9126;
  assign v_9120 = v_9121 & v_9127;
  assign v_9121 = v_9122 & vout_canPeek_9132;
  assign v_9122 = ~vout_canPeek_9123;
  pebbles_core
    pebbles_core_9123
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9124),
       .in0_consume_en(vin0_consume_en_9123),
       .out_canPeek(vout_canPeek_9123),
       .out_peek(vout_peek_9123));
  assign v_9124 = v_9125 | v_9130;
  assign v_9125 = mux_9125(v_9126);
  assign v_9126 = vout_canPeek_9123 & v_9127;
  assign v_9127 = v_9128 & 1'h1;
  assign v_9128 = v_9129 | 1'h0;
  assign v_9129 = ~v_9116;
  assign v_9130 = mux_9130(v_9131);
  assign v_9131 = ~v_9126;
  pebbles_core
    pebbles_core_9132
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9133),
       .in0_consume_en(vin0_consume_en_9132),
       .out_canPeek(vout_canPeek_9132),
       .out_peek(vout_peek_9132));
  assign v_9133 = v_9134 | v_9135;
  assign v_9134 = mux_9134(v_9120);
  assign v_9135 = mux_9135(v_9136);
  assign v_9136 = ~v_9120;
  assign v_9137 = v_9138 & 1'h1;
  assign v_9138 = v_9139 & v_9140;
  assign v_9139 = ~act_9119;
  assign v_9140 = v_9141 | v_9149;
  assign v_9141 = v_9142 | v_9147;
  assign v_9142 = mux_9142(v_9143);
  assign v_9143 = v_9116 & v_9144;
  assign v_9144 = v_9145 & 1'h1;
  assign v_9145 = v_9146 | 1'h0;
  assign v_9146 = ~v_9109;
  assign v_9147 = mux_9147(v_9148);
  assign v_9148 = ~v_9143;
  assign v_9149 = ~v_9116;
  assign v_9150 = v_9151 | v_9152;
  assign v_9151 = mux_9151(v_9118);
  assign v_9152 = mux_9152(v_9137);
  assign v_9154 = v_9155 | v_9174;
  assign v_9155 = act_9156 & 1'h1;
  assign act_9156 = v_9157 | v_9163;
  assign v_9157 = v_9158 & v_9164;
  assign v_9158 = v_9159 & vout_canPeek_9169;
  assign v_9159 = ~vout_canPeek_9160;
  pebbles_core
    pebbles_core_9160
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9161),
       .in0_consume_en(vin0_consume_en_9160),
       .out_canPeek(vout_canPeek_9160),
       .out_peek(vout_peek_9160));
  assign v_9161 = v_9162 | v_9167;
  assign v_9162 = mux_9162(v_9163);
  assign v_9163 = vout_canPeek_9160 & v_9164;
  assign v_9164 = v_9165 & 1'h1;
  assign v_9165 = v_9166 | 1'h0;
  assign v_9166 = ~v_9153;
  assign v_9167 = mux_9167(v_9168);
  assign v_9168 = ~v_9163;
  pebbles_core
    pebbles_core_9169
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9170),
       .in0_consume_en(vin0_consume_en_9169),
       .out_canPeek(vout_canPeek_9169),
       .out_peek(vout_peek_9169));
  assign v_9170 = v_9171 | v_9172;
  assign v_9171 = mux_9171(v_9157);
  assign v_9172 = mux_9172(v_9173);
  assign v_9173 = ~v_9157;
  assign v_9174 = v_9175 & 1'h1;
  assign v_9175 = v_9176 & v_9177;
  assign v_9176 = ~act_9156;
  assign v_9177 = v_9178 | v_9182;
  assign v_9178 = v_9179 | v_9180;
  assign v_9179 = mux_9179(v_9113);
  assign v_9180 = mux_9180(v_9181);
  assign v_9181 = ~v_9113;
  assign v_9182 = ~v_9153;
  assign v_9183 = v_9184 | v_9185;
  assign v_9184 = mux_9184(v_9155);
  assign v_9185 = mux_9185(v_9174);
  assign v_9186 = v_9187 & 1'h1;
  assign v_9187 = v_9188 & v_9189;
  assign v_9188 = ~act_9112;
  assign v_9189 = v_9190 | v_9198;
  assign v_9190 = v_9191 | v_9196;
  assign v_9191 = mux_9191(v_9192);
  assign v_9192 = v_9109 & v_9193;
  assign v_9193 = v_9194 & 1'h1;
  assign v_9194 = v_9195 | 1'h0;
  assign v_9195 = ~v_9102;
  assign v_9196 = mux_9196(v_9197);
  assign v_9197 = ~v_9192;
  assign v_9198 = ~v_9109;
  assign v_9199 = v_9200 | v_9201;
  assign v_9200 = mux_9200(v_9111);
  assign v_9201 = mux_9201(v_9186);
  assign v_9203 = v_9204 | v_9279;
  assign v_9204 = act_9205 & 1'h1;
  assign act_9205 = v_9206 | v_9236;
  assign v_9206 = v_9207 & v_9237;
  assign v_9207 = v_9208 & v_9246;
  assign v_9208 = ~v_9209;
  assign v_9210 = v_9211 | v_9230;
  assign v_9211 = act_9212 & 1'h1;
  assign act_9212 = v_9213 | v_9219;
  assign v_9213 = v_9214 & v_9220;
  assign v_9214 = v_9215 & vout_canPeek_9225;
  assign v_9215 = ~vout_canPeek_9216;
  pebbles_core
    pebbles_core_9216
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9217),
       .in0_consume_en(vin0_consume_en_9216),
       .out_canPeek(vout_canPeek_9216),
       .out_peek(vout_peek_9216));
  assign v_9217 = v_9218 | v_9223;
  assign v_9218 = mux_9218(v_9219);
  assign v_9219 = vout_canPeek_9216 & v_9220;
  assign v_9220 = v_9221 & 1'h1;
  assign v_9221 = v_9222 | 1'h0;
  assign v_9222 = ~v_9209;
  assign v_9223 = mux_9223(v_9224);
  assign v_9224 = ~v_9219;
  pebbles_core
    pebbles_core_9225
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9226),
       .in0_consume_en(vin0_consume_en_9225),
       .out_canPeek(vout_canPeek_9225),
       .out_peek(vout_peek_9225));
  assign v_9226 = v_9227 | v_9228;
  assign v_9227 = mux_9227(v_9213);
  assign v_9228 = mux_9228(v_9229);
  assign v_9229 = ~v_9213;
  assign v_9230 = v_9231 & 1'h1;
  assign v_9231 = v_9232 & v_9233;
  assign v_9232 = ~act_9212;
  assign v_9233 = v_9234 | v_9242;
  assign v_9234 = v_9235 | v_9240;
  assign v_9235 = mux_9235(v_9236);
  assign v_9236 = v_9209 & v_9237;
  assign v_9237 = v_9238 & 1'h1;
  assign v_9238 = v_9239 | 1'h0;
  assign v_9239 = ~v_9202;
  assign v_9240 = mux_9240(v_9241);
  assign v_9241 = ~v_9236;
  assign v_9242 = ~v_9209;
  assign v_9243 = v_9244 | v_9245;
  assign v_9244 = mux_9244(v_9211);
  assign v_9245 = mux_9245(v_9230);
  assign v_9247 = v_9248 | v_9267;
  assign v_9248 = act_9249 & 1'h1;
  assign act_9249 = v_9250 | v_9256;
  assign v_9250 = v_9251 & v_9257;
  assign v_9251 = v_9252 & vout_canPeek_9262;
  assign v_9252 = ~vout_canPeek_9253;
  pebbles_core
    pebbles_core_9253
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9254),
       .in0_consume_en(vin0_consume_en_9253),
       .out_canPeek(vout_canPeek_9253),
       .out_peek(vout_peek_9253));
  assign v_9254 = v_9255 | v_9260;
  assign v_9255 = mux_9255(v_9256);
  assign v_9256 = vout_canPeek_9253 & v_9257;
  assign v_9257 = v_9258 & 1'h1;
  assign v_9258 = v_9259 | 1'h0;
  assign v_9259 = ~v_9246;
  assign v_9260 = mux_9260(v_9261);
  assign v_9261 = ~v_9256;
  pebbles_core
    pebbles_core_9262
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9263),
       .in0_consume_en(vin0_consume_en_9262),
       .out_canPeek(vout_canPeek_9262),
       .out_peek(vout_peek_9262));
  assign v_9263 = v_9264 | v_9265;
  assign v_9264 = mux_9264(v_9250);
  assign v_9265 = mux_9265(v_9266);
  assign v_9266 = ~v_9250;
  assign v_9267 = v_9268 & 1'h1;
  assign v_9268 = v_9269 & v_9270;
  assign v_9269 = ~act_9249;
  assign v_9270 = v_9271 | v_9275;
  assign v_9271 = v_9272 | v_9273;
  assign v_9272 = mux_9272(v_9206);
  assign v_9273 = mux_9273(v_9274);
  assign v_9274 = ~v_9206;
  assign v_9275 = ~v_9246;
  assign v_9276 = v_9277 | v_9278;
  assign v_9277 = mux_9277(v_9248);
  assign v_9278 = mux_9278(v_9267);
  assign v_9279 = v_9280 & 1'h1;
  assign v_9280 = v_9281 & v_9282;
  assign v_9281 = ~act_9205;
  assign v_9282 = v_9283 | v_9287;
  assign v_9283 = v_9284 | v_9285;
  assign v_9284 = mux_9284(v_9106);
  assign v_9285 = mux_9285(v_9286);
  assign v_9286 = ~v_9106;
  assign v_9287 = ~v_9202;
  assign v_9288 = v_9289 | v_9290;
  assign v_9289 = mux_9289(v_9204);
  assign v_9290 = mux_9290(v_9279);
  assign v_9291 = v_9292 & 1'h1;
  assign v_9292 = v_9293 & v_9294;
  assign v_9293 = ~act_9105;
  assign v_9294 = v_9295 | v_9299;
  assign v_9295 = v_9296 | v_9297;
  assign v_9296 = mux_9296(v_8894);
  assign v_9297 = mux_9297(v_9298);
  assign v_9298 = ~v_8894;
  assign v_9299 = ~v_9102;
  assign v_9300 = v_9301 | v_9302;
  assign v_9301 = mux_9301(v_9104);
  assign v_9302 = mux_9302(v_9291);
  assign v_9303 = v_9304 & 1'h1;
  assign v_9304 = v_9305 & v_9306;
  assign v_9305 = ~act_8893;
  assign v_9306 = v_9307 | v_9315;
  assign v_9307 = v_9308 | v_9313;
  assign v_9308 = mux_9308(v_9309);
  assign v_9309 = v_8890 & v_9310;
  assign v_9310 = v_9311 & 1'h1;
  assign v_9311 = v_9312 | 1'h0;
  assign v_9312 = ~v_8883;
  assign v_9313 = mux_9313(v_9314);
  assign v_9314 = ~v_9309;
  assign v_9315 = ~v_8890;
  assign v_9316 = v_9317 | v_9318;
  assign v_9317 = mux_9317(v_8892);
  assign v_9318 = mux_9318(v_9303);
  assign v_9320 = v_9321 | v_9732;
  assign v_9321 = act_9322 & 1'h1;
  assign act_9322 = v_9323 | v_9521;
  assign v_9323 = v_9324 & v_9522;
  assign v_9324 = v_9325 & v_9531;
  assign v_9325 = ~v_9326;
  assign v_9327 = v_9328 | v_9515;
  assign v_9328 = act_9329 & 1'h1;
  assign act_9329 = v_9330 | v_9416;
  assign v_9330 = v_9331 & v_9417;
  assign v_9331 = v_9332 & v_9426;
  assign v_9332 = ~v_9333;
  assign v_9334 = v_9335 | v_9410;
  assign v_9335 = act_9336 & 1'h1;
  assign act_9336 = v_9337 | v_9367;
  assign v_9337 = v_9338 & v_9368;
  assign v_9338 = v_9339 & v_9377;
  assign v_9339 = ~v_9340;
  assign v_9341 = v_9342 | v_9361;
  assign v_9342 = act_9343 & 1'h1;
  assign act_9343 = v_9344 | v_9350;
  assign v_9344 = v_9345 & v_9351;
  assign v_9345 = v_9346 & vout_canPeek_9356;
  assign v_9346 = ~vout_canPeek_9347;
  pebbles_core
    pebbles_core_9347
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9348),
       .in0_consume_en(vin0_consume_en_9347),
       .out_canPeek(vout_canPeek_9347),
       .out_peek(vout_peek_9347));
  assign v_9348 = v_9349 | v_9354;
  assign v_9349 = mux_9349(v_9350);
  assign v_9350 = vout_canPeek_9347 & v_9351;
  assign v_9351 = v_9352 & 1'h1;
  assign v_9352 = v_9353 | 1'h0;
  assign v_9353 = ~v_9340;
  assign v_9354 = mux_9354(v_9355);
  assign v_9355 = ~v_9350;
  pebbles_core
    pebbles_core_9356
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9357),
       .in0_consume_en(vin0_consume_en_9356),
       .out_canPeek(vout_canPeek_9356),
       .out_peek(vout_peek_9356));
  assign v_9357 = v_9358 | v_9359;
  assign v_9358 = mux_9358(v_9344);
  assign v_9359 = mux_9359(v_9360);
  assign v_9360 = ~v_9344;
  assign v_9361 = v_9362 & 1'h1;
  assign v_9362 = v_9363 & v_9364;
  assign v_9363 = ~act_9343;
  assign v_9364 = v_9365 | v_9373;
  assign v_9365 = v_9366 | v_9371;
  assign v_9366 = mux_9366(v_9367);
  assign v_9367 = v_9340 & v_9368;
  assign v_9368 = v_9369 & 1'h1;
  assign v_9369 = v_9370 | 1'h0;
  assign v_9370 = ~v_9333;
  assign v_9371 = mux_9371(v_9372);
  assign v_9372 = ~v_9367;
  assign v_9373 = ~v_9340;
  assign v_9374 = v_9375 | v_9376;
  assign v_9375 = mux_9375(v_9342);
  assign v_9376 = mux_9376(v_9361);
  assign v_9378 = v_9379 | v_9398;
  assign v_9379 = act_9380 & 1'h1;
  assign act_9380 = v_9381 | v_9387;
  assign v_9381 = v_9382 & v_9388;
  assign v_9382 = v_9383 & vout_canPeek_9393;
  assign v_9383 = ~vout_canPeek_9384;
  pebbles_core
    pebbles_core_9384
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9385),
       .in0_consume_en(vin0_consume_en_9384),
       .out_canPeek(vout_canPeek_9384),
       .out_peek(vout_peek_9384));
  assign v_9385 = v_9386 | v_9391;
  assign v_9386 = mux_9386(v_9387);
  assign v_9387 = vout_canPeek_9384 & v_9388;
  assign v_9388 = v_9389 & 1'h1;
  assign v_9389 = v_9390 | 1'h0;
  assign v_9390 = ~v_9377;
  assign v_9391 = mux_9391(v_9392);
  assign v_9392 = ~v_9387;
  pebbles_core
    pebbles_core_9393
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9394),
       .in0_consume_en(vin0_consume_en_9393),
       .out_canPeek(vout_canPeek_9393),
       .out_peek(vout_peek_9393));
  assign v_9394 = v_9395 | v_9396;
  assign v_9395 = mux_9395(v_9381);
  assign v_9396 = mux_9396(v_9397);
  assign v_9397 = ~v_9381;
  assign v_9398 = v_9399 & 1'h1;
  assign v_9399 = v_9400 & v_9401;
  assign v_9400 = ~act_9380;
  assign v_9401 = v_9402 | v_9406;
  assign v_9402 = v_9403 | v_9404;
  assign v_9403 = mux_9403(v_9337);
  assign v_9404 = mux_9404(v_9405);
  assign v_9405 = ~v_9337;
  assign v_9406 = ~v_9377;
  assign v_9407 = v_9408 | v_9409;
  assign v_9408 = mux_9408(v_9379);
  assign v_9409 = mux_9409(v_9398);
  assign v_9410 = v_9411 & 1'h1;
  assign v_9411 = v_9412 & v_9413;
  assign v_9412 = ~act_9336;
  assign v_9413 = v_9414 | v_9422;
  assign v_9414 = v_9415 | v_9420;
  assign v_9415 = mux_9415(v_9416);
  assign v_9416 = v_9333 & v_9417;
  assign v_9417 = v_9418 & 1'h1;
  assign v_9418 = v_9419 | 1'h0;
  assign v_9419 = ~v_9326;
  assign v_9420 = mux_9420(v_9421);
  assign v_9421 = ~v_9416;
  assign v_9422 = ~v_9333;
  assign v_9423 = v_9424 | v_9425;
  assign v_9424 = mux_9424(v_9335);
  assign v_9425 = mux_9425(v_9410);
  assign v_9427 = v_9428 | v_9503;
  assign v_9428 = act_9429 & 1'h1;
  assign act_9429 = v_9430 | v_9460;
  assign v_9430 = v_9431 & v_9461;
  assign v_9431 = v_9432 & v_9470;
  assign v_9432 = ~v_9433;
  assign v_9434 = v_9435 | v_9454;
  assign v_9435 = act_9436 & 1'h1;
  assign act_9436 = v_9437 | v_9443;
  assign v_9437 = v_9438 & v_9444;
  assign v_9438 = v_9439 & vout_canPeek_9449;
  assign v_9439 = ~vout_canPeek_9440;
  pebbles_core
    pebbles_core_9440
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9441),
       .in0_consume_en(vin0_consume_en_9440),
       .out_canPeek(vout_canPeek_9440),
       .out_peek(vout_peek_9440));
  assign v_9441 = v_9442 | v_9447;
  assign v_9442 = mux_9442(v_9443);
  assign v_9443 = vout_canPeek_9440 & v_9444;
  assign v_9444 = v_9445 & 1'h1;
  assign v_9445 = v_9446 | 1'h0;
  assign v_9446 = ~v_9433;
  assign v_9447 = mux_9447(v_9448);
  assign v_9448 = ~v_9443;
  pebbles_core
    pebbles_core_9449
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9450),
       .in0_consume_en(vin0_consume_en_9449),
       .out_canPeek(vout_canPeek_9449),
       .out_peek(vout_peek_9449));
  assign v_9450 = v_9451 | v_9452;
  assign v_9451 = mux_9451(v_9437);
  assign v_9452 = mux_9452(v_9453);
  assign v_9453 = ~v_9437;
  assign v_9454 = v_9455 & 1'h1;
  assign v_9455 = v_9456 & v_9457;
  assign v_9456 = ~act_9436;
  assign v_9457 = v_9458 | v_9466;
  assign v_9458 = v_9459 | v_9464;
  assign v_9459 = mux_9459(v_9460);
  assign v_9460 = v_9433 & v_9461;
  assign v_9461 = v_9462 & 1'h1;
  assign v_9462 = v_9463 | 1'h0;
  assign v_9463 = ~v_9426;
  assign v_9464 = mux_9464(v_9465);
  assign v_9465 = ~v_9460;
  assign v_9466 = ~v_9433;
  assign v_9467 = v_9468 | v_9469;
  assign v_9468 = mux_9468(v_9435);
  assign v_9469 = mux_9469(v_9454);
  assign v_9471 = v_9472 | v_9491;
  assign v_9472 = act_9473 & 1'h1;
  assign act_9473 = v_9474 | v_9480;
  assign v_9474 = v_9475 & v_9481;
  assign v_9475 = v_9476 & vout_canPeek_9486;
  assign v_9476 = ~vout_canPeek_9477;
  pebbles_core
    pebbles_core_9477
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9478),
       .in0_consume_en(vin0_consume_en_9477),
       .out_canPeek(vout_canPeek_9477),
       .out_peek(vout_peek_9477));
  assign v_9478 = v_9479 | v_9484;
  assign v_9479 = mux_9479(v_9480);
  assign v_9480 = vout_canPeek_9477 & v_9481;
  assign v_9481 = v_9482 & 1'h1;
  assign v_9482 = v_9483 | 1'h0;
  assign v_9483 = ~v_9470;
  assign v_9484 = mux_9484(v_9485);
  assign v_9485 = ~v_9480;
  pebbles_core
    pebbles_core_9486
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9487),
       .in0_consume_en(vin0_consume_en_9486),
       .out_canPeek(vout_canPeek_9486),
       .out_peek(vout_peek_9486));
  assign v_9487 = v_9488 | v_9489;
  assign v_9488 = mux_9488(v_9474);
  assign v_9489 = mux_9489(v_9490);
  assign v_9490 = ~v_9474;
  assign v_9491 = v_9492 & 1'h1;
  assign v_9492 = v_9493 & v_9494;
  assign v_9493 = ~act_9473;
  assign v_9494 = v_9495 | v_9499;
  assign v_9495 = v_9496 | v_9497;
  assign v_9496 = mux_9496(v_9430);
  assign v_9497 = mux_9497(v_9498);
  assign v_9498 = ~v_9430;
  assign v_9499 = ~v_9470;
  assign v_9500 = v_9501 | v_9502;
  assign v_9501 = mux_9501(v_9472);
  assign v_9502 = mux_9502(v_9491);
  assign v_9503 = v_9504 & 1'h1;
  assign v_9504 = v_9505 & v_9506;
  assign v_9505 = ~act_9429;
  assign v_9506 = v_9507 | v_9511;
  assign v_9507 = v_9508 | v_9509;
  assign v_9508 = mux_9508(v_9330);
  assign v_9509 = mux_9509(v_9510);
  assign v_9510 = ~v_9330;
  assign v_9511 = ~v_9426;
  assign v_9512 = v_9513 | v_9514;
  assign v_9513 = mux_9513(v_9428);
  assign v_9514 = mux_9514(v_9503);
  assign v_9515 = v_9516 & 1'h1;
  assign v_9516 = v_9517 & v_9518;
  assign v_9517 = ~act_9329;
  assign v_9518 = v_9519 | v_9527;
  assign v_9519 = v_9520 | v_9525;
  assign v_9520 = mux_9520(v_9521);
  assign v_9521 = v_9326 & v_9522;
  assign v_9522 = v_9523 & 1'h1;
  assign v_9523 = v_9524 | 1'h0;
  assign v_9524 = ~v_9319;
  assign v_9525 = mux_9525(v_9526);
  assign v_9526 = ~v_9521;
  assign v_9527 = ~v_9326;
  assign v_9528 = v_9529 | v_9530;
  assign v_9529 = mux_9529(v_9328);
  assign v_9530 = mux_9530(v_9515);
  assign v_9532 = v_9533 | v_9720;
  assign v_9533 = act_9534 & 1'h1;
  assign act_9534 = v_9535 | v_9621;
  assign v_9535 = v_9536 & v_9622;
  assign v_9536 = v_9537 & v_9631;
  assign v_9537 = ~v_9538;
  assign v_9539 = v_9540 | v_9615;
  assign v_9540 = act_9541 & 1'h1;
  assign act_9541 = v_9542 | v_9572;
  assign v_9542 = v_9543 & v_9573;
  assign v_9543 = v_9544 & v_9582;
  assign v_9544 = ~v_9545;
  assign v_9546 = v_9547 | v_9566;
  assign v_9547 = act_9548 & 1'h1;
  assign act_9548 = v_9549 | v_9555;
  assign v_9549 = v_9550 & v_9556;
  assign v_9550 = v_9551 & vout_canPeek_9561;
  assign v_9551 = ~vout_canPeek_9552;
  pebbles_core
    pebbles_core_9552
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9553),
       .in0_consume_en(vin0_consume_en_9552),
       .out_canPeek(vout_canPeek_9552),
       .out_peek(vout_peek_9552));
  assign v_9553 = v_9554 | v_9559;
  assign v_9554 = mux_9554(v_9555);
  assign v_9555 = vout_canPeek_9552 & v_9556;
  assign v_9556 = v_9557 & 1'h1;
  assign v_9557 = v_9558 | 1'h0;
  assign v_9558 = ~v_9545;
  assign v_9559 = mux_9559(v_9560);
  assign v_9560 = ~v_9555;
  pebbles_core
    pebbles_core_9561
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9562),
       .in0_consume_en(vin0_consume_en_9561),
       .out_canPeek(vout_canPeek_9561),
       .out_peek(vout_peek_9561));
  assign v_9562 = v_9563 | v_9564;
  assign v_9563 = mux_9563(v_9549);
  assign v_9564 = mux_9564(v_9565);
  assign v_9565 = ~v_9549;
  assign v_9566 = v_9567 & 1'h1;
  assign v_9567 = v_9568 & v_9569;
  assign v_9568 = ~act_9548;
  assign v_9569 = v_9570 | v_9578;
  assign v_9570 = v_9571 | v_9576;
  assign v_9571 = mux_9571(v_9572);
  assign v_9572 = v_9545 & v_9573;
  assign v_9573 = v_9574 & 1'h1;
  assign v_9574 = v_9575 | 1'h0;
  assign v_9575 = ~v_9538;
  assign v_9576 = mux_9576(v_9577);
  assign v_9577 = ~v_9572;
  assign v_9578 = ~v_9545;
  assign v_9579 = v_9580 | v_9581;
  assign v_9580 = mux_9580(v_9547);
  assign v_9581 = mux_9581(v_9566);
  assign v_9583 = v_9584 | v_9603;
  assign v_9584 = act_9585 & 1'h1;
  assign act_9585 = v_9586 | v_9592;
  assign v_9586 = v_9587 & v_9593;
  assign v_9587 = v_9588 & vout_canPeek_9598;
  assign v_9588 = ~vout_canPeek_9589;
  pebbles_core
    pebbles_core_9589
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9590),
       .in0_consume_en(vin0_consume_en_9589),
       .out_canPeek(vout_canPeek_9589),
       .out_peek(vout_peek_9589));
  assign v_9590 = v_9591 | v_9596;
  assign v_9591 = mux_9591(v_9592);
  assign v_9592 = vout_canPeek_9589 & v_9593;
  assign v_9593 = v_9594 & 1'h1;
  assign v_9594 = v_9595 | 1'h0;
  assign v_9595 = ~v_9582;
  assign v_9596 = mux_9596(v_9597);
  assign v_9597 = ~v_9592;
  pebbles_core
    pebbles_core_9598
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9599),
       .in0_consume_en(vin0_consume_en_9598),
       .out_canPeek(vout_canPeek_9598),
       .out_peek(vout_peek_9598));
  assign v_9599 = v_9600 | v_9601;
  assign v_9600 = mux_9600(v_9586);
  assign v_9601 = mux_9601(v_9602);
  assign v_9602 = ~v_9586;
  assign v_9603 = v_9604 & 1'h1;
  assign v_9604 = v_9605 & v_9606;
  assign v_9605 = ~act_9585;
  assign v_9606 = v_9607 | v_9611;
  assign v_9607 = v_9608 | v_9609;
  assign v_9608 = mux_9608(v_9542);
  assign v_9609 = mux_9609(v_9610);
  assign v_9610 = ~v_9542;
  assign v_9611 = ~v_9582;
  assign v_9612 = v_9613 | v_9614;
  assign v_9613 = mux_9613(v_9584);
  assign v_9614 = mux_9614(v_9603);
  assign v_9615 = v_9616 & 1'h1;
  assign v_9616 = v_9617 & v_9618;
  assign v_9617 = ~act_9541;
  assign v_9618 = v_9619 | v_9627;
  assign v_9619 = v_9620 | v_9625;
  assign v_9620 = mux_9620(v_9621);
  assign v_9621 = v_9538 & v_9622;
  assign v_9622 = v_9623 & 1'h1;
  assign v_9623 = v_9624 | 1'h0;
  assign v_9624 = ~v_9531;
  assign v_9625 = mux_9625(v_9626);
  assign v_9626 = ~v_9621;
  assign v_9627 = ~v_9538;
  assign v_9628 = v_9629 | v_9630;
  assign v_9629 = mux_9629(v_9540);
  assign v_9630 = mux_9630(v_9615);
  assign v_9632 = v_9633 | v_9708;
  assign v_9633 = act_9634 & 1'h1;
  assign act_9634 = v_9635 | v_9665;
  assign v_9635 = v_9636 & v_9666;
  assign v_9636 = v_9637 & v_9675;
  assign v_9637 = ~v_9638;
  assign v_9639 = v_9640 | v_9659;
  assign v_9640 = act_9641 & 1'h1;
  assign act_9641 = v_9642 | v_9648;
  assign v_9642 = v_9643 & v_9649;
  assign v_9643 = v_9644 & vout_canPeek_9654;
  assign v_9644 = ~vout_canPeek_9645;
  pebbles_core
    pebbles_core_9645
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9646),
       .in0_consume_en(vin0_consume_en_9645),
       .out_canPeek(vout_canPeek_9645),
       .out_peek(vout_peek_9645));
  assign v_9646 = v_9647 | v_9652;
  assign v_9647 = mux_9647(v_9648);
  assign v_9648 = vout_canPeek_9645 & v_9649;
  assign v_9649 = v_9650 & 1'h1;
  assign v_9650 = v_9651 | 1'h0;
  assign v_9651 = ~v_9638;
  assign v_9652 = mux_9652(v_9653);
  assign v_9653 = ~v_9648;
  pebbles_core
    pebbles_core_9654
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9655),
       .in0_consume_en(vin0_consume_en_9654),
       .out_canPeek(vout_canPeek_9654),
       .out_peek(vout_peek_9654));
  assign v_9655 = v_9656 | v_9657;
  assign v_9656 = mux_9656(v_9642);
  assign v_9657 = mux_9657(v_9658);
  assign v_9658 = ~v_9642;
  assign v_9659 = v_9660 & 1'h1;
  assign v_9660 = v_9661 & v_9662;
  assign v_9661 = ~act_9641;
  assign v_9662 = v_9663 | v_9671;
  assign v_9663 = v_9664 | v_9669;
  assign v_9664 = mux_9664(v_9665);
  assign v_9665 = v_9638 & v_9666;
  assign v_9666 = v_9667 & 1'h1;
  assign v_9667 = v_9668 | 1'h0;
  assign v_9668 = ~v_9631;
  assign v_9669 = mux_9669(v_9670);
  assign v_9670 = ~v_9665;
  assign v_9671 = ~v_9638;
  assign v_9672 = v_9673 | v_9674;
  assign v_9673 = mux_9673(v_9640);
  assign v_9674 = mux_9674(v_9659);
  assign v_9676 = v_9677 | v_9696;
  assign v_9677 = act_9678 & 1'h1;
  assign act_9678 = v_9679 | v_9685;
  assign v_9679 = v_9680 & v_9686;
  assign v_9680 = v_9681 & vout_canPeek_9691;
  assign v_9681 = ~vout_canPeek_9682;
  pebbles_core
    pebbles_core_9682
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9683),
       .in0_consume_en(vin0_consume_en_9682),
       .out_canPeek(vout_canPeek_9682),
       .out_peek(vout_peek_9682));
  assign v_9683 = v_9684 | v_9689;
  assign v_9684 = mux_9684(v_9685);
  assign v_9685 = vout_canPeek_9682 & v_9686;
  assign v_9686 = v_9687 & 1'h1;
  assign v_9687 = v_9688 | 1'h0;
  assign v_9688 = ~v_9675;
  assign v_9689 = mux_9689(v_9690);
  assign v_9690 = ~v_9685;
  pebbles_core
    pebbles_core_9691
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9692),
       .in0_consume_en(vin0_consume_en_9691),
       .out_canPeek(vout_canPeek_9691),
       .out_peek(vout_peek_9691));
  assign v_9692 = v_9693 | v_9694;
  assign v_9693 = mux_9693(v_9679);
  assign v_9694 = mux_9694(v_9695);
  assign v_9695 = ~v_9679;
  assign v_9696 = v_9697 & 1'h1;
  assign v_9697 = v_9698 & v_9699;
  assign v_9698 = ~act_9678;
  assign v_9699 = v_9700 | v_9704;
  assign v_9700 = v_9701 | v_9702;
  assign v_9701 = mux_9701(v_9635);
  assign v_9702 = mux_9702(v_9703);
  assign v_9703 = ~v_9635;
  assign v_9704 = ~v_9675;
  assign v_9705 = v_9706 | v_9707;
  assign v_9706 = mux_9706(v_9677);
  assign v_9707 = mux_9707(v_9696);
  assign v_9708 = v_9709 & 1'h1;
  assign v_9709 = v_9710 & v_9711;
  assign v_9710 = ~act_9634;
  assign v_9711 = v_9712 | v_9716;
  assign v_9712 = v_9713 | v_9714;
  assign v_9713 = mux_9713(v_9535);
  assign v_9714 = mux_9714(v_9715);
  assign v_9715 = ~v_9535;
  assign v_9716 = ~v_9631;
  assign v_9717 = v_9718 | v_9719;
  assign v_9718 = mux_9718(v_9633);
  assign v_9719 = mux_9719(v_9708);
  assign v_9720 = v_9721 & 1'h1;
  assign v_9721 = v_9722 & v_9723;
  assign v_9722 = ~act_9534;
  assign v_9723 = v_9724 | v_9728;
  assign v_9724 = v_9725 | v_9726;
  assign v_9725 = mux_9725(v_9323);
  assign v_9726 = mux_9726(v_9727);
  assign v_9727 = ~v_9323;
  assign v_9728 = ~v_9531;
  assign v_9729 = v_9730 | v_9731;
  assign v_9730 = mux_9730(v_9533);
  assign v_9731 = mux_9731(v_9720);
  assign v_9732 = v_9733 & 1'h1;
  assign v_9733 = v_9734 & v_9735;
  assign v_9734 = ~act_9322;
  assign v_9735 = v_9736 | v_9740;
  assign v_9736 = v_9737 | v_9738;
  assign v_9737 = mux_9737(v_8887);
  assign v_9738 = mux_9738(v_9739);
  assign v_9739 = ~v_8887;
  assign v_9740 = ~v_9319;
  assign v_9741 = v_9742 | v_9743;
  assign v_9742 = mux_9742(v_9321);
  assign v_9743 = mux_9743(v_9732);
  assign v_9744 = v_9745 & 1'h1;
  assign v_9745 = v_9746 & v_9747;
  assign v_9746 = ~act_8886;
  assign v_9747 = v_9748 | v_9752;
  assign v_9748 = v_9749 | v_9750;
  assign v_9749 = mux_9749(v_8003);
  assign v_9750 = mux_9750(v_9751);
  assign v_9751 = ~v_8003;
  assign v_9752 = ~v_8883;
  assign v_9753 = v_9754 | v_9755;
  assign v_9754 = mux_9754(v_8885);
  assign v_9755 = mux_9755(v_9744);
  assign v_9756 = v_9757 & 1'h1;
  assign v_9757 = v_9758 & v_9759;
  assign v_9758 = ~act_8002;
  assign v_9759 = v_9760 | v_9768;
  assign v_9760 = v_9761 | v_9766;
  assign v_9761 = mux_9761(v_9762);
  assign v_9762 = v_7999 & v_9763;
  assign v_9763 = v_9764 & 1'h1;
  assign v_9764 = v_9765 | 1'h0;
  assign v_9765 = ~v_7992;
  assign v_9766 = mux_9766(v_9767);
  assign v_9767 = ~v_9762;
  assign v_9768 = ~v_7999;
  assign v_9769 = v_9770 | v_9771;
  assign v_9770 = mux_9770(v_8001);
  assign v_9771 = mux_9771(v_9756);
  assign v_9773 = v_9774 | v_11529;
  assign v_9774 = act_9775 & 1'h1;
  assign act_9775 = v_9776 | v_10646;
  assign v_9776 = v_9777 & v_10647;
  assign v_9777 = v_9778 & v_10656;
  assign v_9778 = ~v_9779;
  assign v_9780 = v_9781 | v_10640;
  assign v_9781 = act_9782 & 1'h1;
  assign act_9782 = v_9783 | v_10205;
  assign v_9783 = v_9784 & v_10206;
  assign v_9784 = v_9785 & v_10215;
  assign v_9785 = ~v_9786;
  assign v_9787 = v_9788 | v_10199;
  assign v_9788 = act_9789 & 1'h1;
  assign act_9789 = v_9790 | v_9988;
  assign v_9790 = v_9791 & v_9989;
  assign v_9791 = v_9792 & v_9998;
  assign v_9792 = ~v_9793;
  assign v_9794 = v_9795 | v_9982;
  assign v_9795 = act_9796 & 1'h1;
  assign act_9796 = v_9797 | v_9883;
  assign v_9797 = v_9798 & v_9884;
  assign v_9798 = v_9799 & v_9893;
  assign v_9799 = ~v_9800;
  assign v_9801 = v_9802 | v_9877;
  assign v_9802 = act_9803 & 1'h1;
  assign act_9803 = v_9804 | v_9834;
  assign v_9804 = v_9805 & v_9835;
  assign v_9805 = v_9806 & v_9844;
  assign v_9806 = ~v_9807;
  assign v_9808 = v_9809 | v_9828;
  assign v_9809 = act_9810 & 1'h1;
  assign act_9810 = v_9811 | v_9817;
  assign v_9811 = v_9812 & v_9818;
  assign v_9812 = v_9813 & vout_canPeek_9823;
  assign v_9813 = ~vout_canPeek_9814;
  pebbles_core
    pebbles_core_9814
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9815),
       .in0_consume_en(vin0_consume_en_9814),
       .out_canPeek(vout_canPeek_9814),
       .out_peek(vout_peek_9814));
  assign v_9815 = v_9816 | v_9821;
  assign v_9816 = mux_9816(v_9817);
  assign v_9817 = vout_canPeek_9814 & v_9818;
  assign v_9818 = v_9819 & 1'h1;
  assign v_9819 = v_9820 | 1'h0;
  assign v_9820 = ~v_9807;
  assign v_9821 = mux_9821(v_9822);
  assign v_9822 = ~v_9817;
  pebbles_core
    pebbles_core_9823
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9824),
       .in0_consume_en(vin0_consume_en_9823),
       .out_canPeek(vout_canPeek_9823),
       .out_peek(vout_peek_9823));
  assign v_9824 = v_9825 | v_9826;
  assign v_9825 = mux_9825(v_9811);
  assign v_9826 = mux_9826(v_9827);
  assign v_9827 = ~v_9811;
  assign v_9828 = v_9829 & 1'h1;
  assign v_9829 = v_9830 & v_9831;
  assign v_9830 = ~act_9810;
  assign v_9831 = v_9832 | v_9840;
  assign v_9832 = v_9833 | v_9838;
  assign v_9833 = mux_9833(v_9834);
  assign v_9834 = v_9807 & v_9835;
  assign v_9835 = v_9836 & 1'h1;
  assign v_9836 = v_9837 | 1'h0;
  assign v_9837 = ~v_9800;
  assign v_9838 = mux_9838(v_9839);
  assign v_9839 = ~v_9834;
  assign v_9840 = ~v_9807;
  assign v_9841 = v_9842 | v_9843;
  assign v_9842 = mux_9842(v_9809);
  assign v_9843 = mux_9843(v_9828);
  assign v_9845 = v_9846 | v_9865;
  assign v_9846 = act_9847 & 1'h1;
  assign act_9847 = v_9848 | v_9854;
  assign v_9848 = v_9849 & v_9855;
  assign v_9849 = v_9850 & vout_canPeek_9860;
  assign v_9850 = ~vout_canPeek_9851;
  pebbles_core
    pebbles_core_9851
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9852),
       .in0_consume_en(vin0_consume_en_9851),
       .out_canPeek(vout_canPeek_9851),
       .out_peek(vout_peek_9851));
  assign v_9852 = v_9853 | v_9858;
  assign v_9853 = mux_9853(v_9854);
  assign v_9854 = vout_canPeek_9851 & v_9855;
  assign v_9855 = v_9856 & 1'h1;
  assign v_9856 = v_9857 | 1'h0;
  assign v_9857 = ~v_9844;
  assign v_9858 = mux_9858(v_9859);
  assign v_9859 = ~v_9854;
  pebbles_core
    pebbles_core_9860
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9861),
       .in0_consume_en(vin0_consume_en_9860),
       .out_canPeek(vout_canPeek_9860),
       .out_peek(vout_peek_9860));
  assign v_9861 = v_9862 | v_9863;
  assign v_9862 = mux_9862(v_9848);
  assign v_9863 = mux_9863(v_9864);
  assign v_9864 = ~v_9848;
  assign v_9865 = v_9866 & 1'h1;
  assign v_9866 = v_9867 & v_9868;
  assign v_9867 = ~act_9847;
  assign v_9868 = v_9869 | v_9873;
  assign v_9869 = v_9870 | v_9871;
  assign v_9870 = mux_9870(v_9804);
  assign v_9871 = mux_9871(v_9872);
  assign v_9872 = ~v_9804;
  assign v_9873 = ~v_9844;
  assign v_9874 = v_9875 | v_9876;
  assign v_9875 = mux_9875(v_9846);
  assign v_9876 = mux_9876(v_9865);
  assign v_9877 = v_9878 & 1'h1;
  assign v_9878 = v_9879 & v_9880;
  assign v_9879 = ~act_9803;
  assign v_9880 = v_9881 | v_9889;
  assign v_9881 = v_9882 | v_9887;
  assign v_9882 = mux_9882(v_9883);
  assign v_9883 = v_9800 & v_9884;
  assign v_9884 = v_9885 & 1'h1;
  assign v_9885 = v_9886 | 1'h0;
  assign v_9886 = ~v_9793;
  assign v_9887 = mux_9887(v_9888);
  assign v_9888 = ~v_9883;
  assign v_9889 = ~v_9800;
  assign v_9890 = v_9891 | v_9892;
  assign v_9891 = mux_9891(v_9802);
  assign v_9892 = mux_9892(v_9877);
  assign v_9894 = v_9895 | v_9970;
  assign v_9895 = act_9896 & 1'h1;
  assign act_9896 = v_9897 | v_9927;
  assign v_9897 = v_9898 & v_9928;
  assign v_9898 = v_9899 & v_9937;
  assign v_9899 = ~v_9900;
  assign v_9901 = v_9902 | v_9921;
  assign v_9902 = act_9903 & 1'h1;
  assign act_9903 = v_9904 | v_9910;
  assign v_9904 = v_9905 & v_9911;
  assign v_9905 = v_9906 & vout_canPeek_9916;
  assign v_9906 = ~vout_canPeek_9907;
  pebbles_core
    pebbles_core_9907
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9908),
       .in0_consume_en(vin0_consume_en_9907),
       .out_canPeek(vout_canPeek_9907),
       .out_peek(vout_peek_9907));
  assign v_9908 = v_9909 | v_9914;
  assign v_9909 = mux_9909(v_9910);
  assign v_9910 = vout_canPeek_9907 & v_9911;
  assign v_9911 = v_9912 & 1'h1;
  assign v_9912 = v_9913 | 1'h0;
  assign v_9913 = ~v_9900;
  assign v_9914 = mux_9914(v_9915);
  assign v_9915 = ~v_9910;
  pebbles_core
    pebbles_core_9916
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9917),
       .in0_consume_en(vin0_consume_en_9916),
       .out_canPeek(vout_canPeek_9916),
       .out_peek(vout_peek_9916));
  assign v_9917 = v_9918 | v_9919;
  assign v_9918 = mux_9918(v_9904);
  assign v_9919 = mux_9919(v_9920);
  assign v_9920 = ~v_9904;
  assign v_9921 = v_9922 & 1'h1;
  assign v_9922 = v_9923 & v_9924;
  assign v_9923 = ~act_9903;
  assign v_9924 = v_9925 | v_9933;
  assign v_9925 = v_9926 | v_9931;
  assign v_9926 = mux_9926(v_9927);
  assign v_9927 = v_9900 & v_9928;
  assign v_9928 = v_9929 & 1'h1;
  assign v_9929 = v_9930 | 1'h0;
  assign v_9930 = ~v_9893;
  assign v_9931 = mux_9931(v_9932);
  assign v_9932 = ~v_9927;
  assign v_9933 = ~v_9900;
  assign v_9934 = v_9935 | v_9936;
  assign v_9935 = mux_9935(v_9902);
  assign v_9936 = mux_9936(v_9921);
  assign v_9938 = v_9939 | v_9958;
  assign v_9939 = act_9940 & 1'h1;
  assign act_9940 = v_9941 | v_9947;
  assign v_9941 = v_9942 & v_9948;
  assign v_9942 = v_9943 & vout_canPeek_9953;
  assign v_9943 = ~vout_canPeek_9944;
  pebbles_core
    pebbles_core_9944
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9945),
       .in0_consume_en(vin0_consume_en_9944),
       .out_canPeek(vout_canPeek_9944),
       .out_peek(vout_peek_9944));
  assign v_9945 = v_9946 | v_9951;
  assign v_9946 = mux_9946(v_9947);
  assign v_9947 = vout_canPeek_9944 & v_9948;
  assign v_9948 = v_9949 & 1'h1;
  assign v_9949 = v_9950 | 1'h0;
  assign v_9950 = ~v_9937;
  assign v_9951 = mux_9951(v_9952);
  assign v_9952 = ~v_9947;
  pebbles_core
    pebbles_core_9953
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_9954),
       .in0_consume_en(vin0_consume_en_9953),
       .out_canPeek(vout_canPeek_9953),
       .out_peek(vout_peek_9953));
  assign v_9954 = v_9955 | v_9956;
  assign v_9955 = mux_9955(v_9941);
  assign v_9956 = mux_9956(v_9957);
  assign v_9957 = ~v_9941;
  assign v_9958 = v_9959 & 1'h1;
  assign v_9959 = v_9960 & v_9961;
  assign v_9960 = ~act_9940;
  assign v_9961 = v_9962 | v_9966;
  assign v_9962 = v_9963 | v_9964;
  assign v_9963 = mux_9963(v_9897);
  assign v_9964 = mux_9964(v_9965);
  assign v_9965 = ~v_9897;
  assign v_9966 = ~v_9937;
  assign v_9967 = v_9968 | v_9969;
  assign v_9968 = mux_9968(v_9939);
  assign v_9969 = mux_9969(v_9958);
  assign v_9970 = v_9971 & 1'h1;
  assign v_9971 = v_9972 & v_9973;
  assign v_9972 = ~act_9896;
  assign v_9973 = v_9974 | v_9978;
  assign v_9974 = v_9975 | v_9976;
  assign v_9975 = mux_9975(v_9797);
  assign v_9976 = mux_9976(v_9977);
  assign v_9977 = ~v_9797;
  assign v_9978 = ~v_9893;
  assign v_9979 = v_9980 | v_9981;
  assign v_9980 = mux_9980(v_9895);
  assign v_9981 = mux_9981(v_9970);
  assign v_9982 = v_9983 & 1'h1;
  assign v_9983 = v_9984 & v_9985;
  assign v_9984 = ~act_9796;
  assign v_9985 = v_9986 | v_9994;
  assign v_9986 = v_9987 | v_9992;
  assign v_9987 = mux_9987(v_9988);
  assign v_9988 = v_9793 & v_9989;
  assign v_9989 = v_9990 & 1'h1;
  assign v_9990 = v_9991 | 1'h0;
  assign v_9991 = ~v_9786;
  assign v_9992 = mux_9992(v_9993);
  assign v_9993 = ~v_9988;
  assign v_9994 = ~v_9793;
  assign v_9995 = v_9996 | v_9997;
  assign v_9996 = mux_9996(v_9795);
  assign v_9997 = mux_9997(v_9982);
  assign v_9999 = v_10000 | v_10187;
  assign v_10000 = act_10001 & 1'h1;
  assign act_10001 = v_10002 | v_10088;
  assign v_10002 = v_10003 & v_10089;
  assign v_10003 = v_10004 & v_10098;
  assign v_10004 = ~v_10005;
  assign v_10006 = v_10007 | v_10082;
  assign v_10007 = act_10008 & 1'h1;
  assign act_10008 = v_10009 | v_10039;
  assign v_10009 = v_10010 & v_10040;
  assign v_10010 = v_10011 & v_10049;
  assign v_10011 = ~v_10012;
  assign v_10013 = v_10014 | v_10033;
  assign v_10014 = act_10015 & 1'h1;
  assign act_10015 = v_10016 | v_10022;
  assign v_10016 = v_10017 & v_10023;
  assign v_10017 = v_10018 & vout_canPeek_10028;
  assign v_10018 = ~vout_canPeek_10019;
  pebbles_core
    pebbles_core_10019
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10020),
       .in0_consume_en(vin0_consume_en_10019),
       .out_canPeek(vout_canPeek_10019),
       .out_peek(vout_peek_10019));
  assign v_10020 = v_10021 | v_10026;
  assign v_10021 = mux_10021(v_10022);
  assign v_10022 = vout_canPeek_10019 & v_10023;
  assign v_10023 = v_10024 & 1'h1;
  assign v_10024 = v_10025 | 1'h0;
  assign v_10025 = ~v_10012;
  assign v_10026 = mux_10026(v_10027);
  assign v_10027 = ~v_10022;
  pebbles_core
    pebbles_core_10028
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10029),
       .in0_consume_en(vin0_consume_en_10028),
       .out_canPeek(vout_canPeek_10028),
       .out_peek(vout_peek_10028));
  assign v_10029 = v_10030 | v_10031;
  assign v_10030 = mux_10030(v_10016);
  assign v_10031 = mux_10031(v_10032);
  assign v_10032 = ~v_10016;
  assign v_10033 = v_10034 & 1'h1;
  assign v_10034 = v_10035 & v_10036;
  assign v_10035 = ~act_10015;
  assign v_10036 = v_10037 | v_10045;
  assign v_10037 = v_10038 | v_10043;
  assign v_10038 = mux_10038(v_10039);
  assign v_10039 = v_10012 & v_10040;
  assign v_10040 = v_10041 & 1'h1;
  assign v_10041 = v_10042 | 1'h0;
  assign v_10042 = ~v_10005;
  assign v_10043 = mux_10043(v_10044);
  assign v_10044 = ~v_10039;
  assign v_10045 = ~v_10012;
  assign v_10046 = v_10047 | v_10048;
  assign v_10047 = mux_10047(v_10014);
  assign v_10048 = mux_10048(v_10033);
  assign v_10050 = v_10051 | v_10070;
  assign v_10051 = act_10052 & 1'h1;
  assign act_10052 = v_10053 | v_10059;
  assign v_10053 = v_10054 & v_10060;
  assign v_10054 = v_10055 & vout_canPeek_10065;
  assign v_10055 = ~vout_canPeek_10056;
  pebbles_core
    pebbles_core_10056
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10057),
       .in0_consume_en(vin0_consume_en_10056),
       .out_canPeek(vout_canPeek_10056),
       .out_peek(vout_peek_10056));
  assign v_10057 = v_10058 | v_10063;
  assign v_10058 = mux_10058(v_10059);
  assign v_10059 = vout_canPeek_10056 & v_10060;
  assign v_10060 = v_10061 & 1'h1;
  assign v_10061 = v_10062 | 1'h0;
  assign v_10062 = ~v_10049;
  assign v_10063 = mux_10063(v_10064);
  assign v_10064 = ~v_10059;
  pebbles_core
    pebbles_core_10065
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10066),
       .in0_consume_en(vin0_consume_en_10065),
       .out_canPeek(vout_canPeek_10065),
       .out_peek(vout_peek_10065));
  assign v_10066 = v_10067 | v_10068;
  assign v_10067 = mux_10067(v_10053);
  assign v_10068 = mux_10068(v_10069);
  assign v_10069 = ~v_10053;
  assign v_10070 = v_10071 & 1'h1;
  assign v_10071 = v_10072 & v_10073;
  assign v_10072 = ~act_10052;
  assign v_10073 = v_10074 | v_10078;
  assign v_10074 = v_10075 | v_10076;
  assign v_10075 = mux_10075(v_10009);
  assign v_10076 = mux_10076(v_10077);
  assign v_10077 = ~v_10009;
  assign v_10078 = ~v_10049;
  assign v_10079 = v_10080 | v_10081;
  assign v_10080 = mux_10080(v_10051);
  assign v_10081 = mux_10081(v_10070);
  assign v_10082 = v_10083 & 1'h1;
  assign v_10083 = v_10084 & v_10085;
  assign v_10084 = ~act_10008;
  assign v_10085 = v_10086 | v_10094;
  assign v_10086 = v_10087 | v_10092;
  assign v_10087 = mux_10087(v_10088);
  assign v_10088 = v_10005 & v_10089;
  assign v_10089 = v_10090 & 1'h1;
  assign v_10090 = v_10091 | 1'h0;
  assign v_10091 = ~v_9998;
  assign v_10092 = mux_10092(v_10093);
  assign v_10093 = ~v_10088;
  assign v_10094 = ~v_10005;
  assign v_10095 = v_10096 | v_10097;
  assign v_10096 = mux_10096(v_10007);
  assign v_10097 = mux_10097(v_10082);
  assign v_10099 = v_10100 | v_10175;
  assign v_10100 = act_10101 & 1'h1;
  assign act_10101 = v_10102 | v_10132;
  assign v_10102 = v_10103 & v_10133;
  assign v_10103 = v_10104 & v_10142;
  assign v_10104 = ~v_10105;
  assign v_10106 = v_10107 | v_10126;
  assign v_10107 = act_10108 & 1'h1;
  assign act_10108 = v_10109 | v_10115;
  assign v_10109 = v_10110 & v_10116;
  assign v_10110 = v_10111 & vout_canPeek_10121;
  assign v_10111 = ~vout_canPeek_10112;
  pebbles_core
    pebbles_core_10112
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10113),
       .in0_consume_en(vin0_consume_en_10112),
       .out_canPeek(vout_canPeek_10112),
       .out_peek(vout_peek_10112));
  assign v_10113 = v_10114 | v_10119;
  assign v_10114 = mux_10114(v_10115);
  assign v_10115 = vout_canPeek_10112 & v_10116;
  assign v_10116 = v_10117 & 1'h1;
  assign v_10117 = v_10118 | 1'h0;
  assign v_10118 = ~v_10105;
  assign v_10119 = mux_10119(v_10120);
  assign v_10120 = ~v_10115;
  pebbles_core
    pebbles_core_10121
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10122),
       .in0_consume_en(vin0_consume_en_10121),
       .out_canPeek(vout_canPeek_10121),
       .out_peek(vout_peek_10121));
  assign v_10122 = v_10123 | v_10124;
  assign v_10123 = mux_10123(v_10109);
  assign v_10124 = mux_10124(v_10125);
  assign v_10125 = ~v_10109;
  assign v_10126 = v_10127 & 1'h1;
  assign v_10127 = v_10128 & v_10129;
  assign v_10128 = ~act_10108;
  assign v_10129 = v_10130 | v_10138;
  assign v_10130 = v_10131 | v_10136;
  assign v_10131 = mux_10131(v_10132);
  assign v_10132 = v_10105 & v_10133;
  assign v_10133 = v_10134 & 1'h1;
  assign v_10134 = v_10135 | 1'h0;
  assign v_10135 = ~v_10098;
  assign v_10136 = mux_10136(v_10137);
  assign v_10137 = ~v_10132;
  assign v_10138 = ~v_10105;
  assign v_10139 = v_10140 | v_10141;
  assign v_10140 = mux_10140(v_10107);
  assign v_10141 = mux_10141(v_10126);
  assign v_10143 = v_10144 | v_10163;
  assign v_10144 = act_10145 & 1'h1;
  assign act_10145 = v_10146 | v_10152;
  assign v_10146 = v_10147 & v_10153;
  assign v_10147 = v_10148 & vout_canPeek_10158;
  assign v_10148 = ~vout_canPeek_10149;
  pebbles_core
    pebbles_core_10149
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10150),
       .in0_consume_en(vin0_consume_en_10149),
       .out_canPeek(vout_canPeek_10149),
       .out_peek(vout_peek_10149));
  assign v_10150 = v_10151 | v_10156;
  assign v_10151 = mux_10151(v_10152);
  assign v_10152 = vout_canPeek_10149 & v_10153;
  assign v_10153 = v_10154 & 1'h1;
  assign v_10154 = v_10155 | 1'h0;
  assign v_10155 = ~v_10142;
  assign v_10156 = mux_10156(v_10157);
  assign v_10157 = ~v_10152;
  pebbles_core
    pebbles_core_10158
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10159),
       .in0_consume_en(vin0_consume_en_10158),
       .out_canPeek(vout_canPeek_10158),
       .out_peek(vout_peek_10158));
  assign v_10159 = v_10160 | v_10161;
  assign v_10160 = mux_10160(v_10146);
  assign v_10161 = mux_10161(v_10162);
  assign v_10162 = ~v_10146;
  assign v_10163 = v_10164 & 1'h1;
  assign v_10164 = v_10165 & v_10166;
  assign v_10165 = ~act_10145;
  assign v_10166 = v_10167 | v_10171;
  assign v_10167 = v_10168 | v_10169;
  assign v_10168 = mux_10168(v_10102);
  assign v_10169 = mux_10169(v_10170);
  assign v_10170 = ~v_10102;
  assign v_10171 = ~v_10142;
  assign v_10172 = v_10173 | v_10174;
  assign v_10173 = mux_10173(v_10144);
  assign v_10174 = mux_10174(v_10163);
  assign v_10175 = v_10176 & 1'h1;
  assign v_10176 = v_10177 & v_10178;
  assign v_10177 = ~act_10101;
  assign v_10178 = v_10179 | v_10183;
  assign v_10179 = v_10180 | v_10181;
  assign v_10180 = mux_10180(v_10002);
  assign v_10181 = mux_10181(v_10182);
  assign v_10182 = ~v_10002;
  assign v_10183 = ~v_10098;
  assign v_10184 = v_10185 | v_10186;
  assign v_10185 = mux_10185(v_10100);
  assign v_10186 = mux_10186(v_10175);
  assign v_10187 = v_10188 & 1'h1;
  assign v_10188 = v_10189 & v_10190;
  assign v_10189 = ~act_10001;
  assign v_10190 = v_10191 | v_10195;
  assign v_10191 = v_10192 | v_10193;
  assign v_10192 = mux_10192(v_9790);
  assign v_10193 = mux_10193(v_10194);
  assign v_10194 = ~v_9790;
  assign v_10195 = ~v_9998;
  assign v_10196 = v_10197 | v_10198;
  assign v_10197 = mux_10197(v_10000);
  assign v_10198 = mux_10198(v_10187);
  assign v_10199 = v_10200 & 1'h1;
  assign v_10200 = v_10201 & v_10202;
  assign v_10201 = ~act_9789;
  assign v_10202 = v_10203 | v_10211;
  assign v_10203 = v_10204 | v_10209;
  assign v_10204 = mux_10204(v_10205);
  assign v_10205 = v_9786 & v_10206;
  assign v_10206 = v_10207 & 1'h1;
  assign v_10207 = v_10208 | 1'h0;
  assign v_10208 = ~v_9779;
  assign v_10209 = mux_10209(v_10210);
  assign v_10210 = ~v_10205;
  assign v_10211 = ~v_9786;
  assign v_10212 = v_10213 | v_10214;
  assign v_10213 = mux_10213(v_9788);
  assign v_10214 = mux_10214(v_10199);
  assign v_10216 = v_10217 | v_10628;
  assign v_10217 = act_10218 & 1'h1;
  assign act_10218 = v_10219 | v_10417;
  assign v_10219 = v_10220 & v_10418;
  assign v_10220 = v_10221 & v_10427;
  assign v_10221 = ~v_10222;
  assign v_10223 = v_10224 | v_10411;
  assign v_10224 = act_10225 & 1'h1;
  assign act_10225 = v_10226 | v_10312;
  assign v_10226 = v_10227 & v_10313;
  assign v_10227 = v_10228 & v_10322;
  assign v_10228 = ~v_10229;
  assign v_10230 = v_10231 | v_10306;
  assign v_10231 = act_10232 & 1'h1;
  assign act_10232 = v_10233 | v_10263;
  assign v_10233 = v_10234 & v_10264;
  assign v_10234 = v_10235 & v_10273;
  assign v_10235 = ~v_10236;
  assign v_10237 = v_10238 | v_10257;
  assign v_10238 = act_10239 & 1'h1;
  assign act_10239 = v_10240 | v_10246;
  assign v_10240 = v_10241 & v_10247;
  assign v_10241 = v_10242 & vout_canPeek_10252;
  assign v_10242 = ~vout_canPeek_10243;
  pebbles_core
    pebbles_core_10243
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10244),
       .in0_consume_en(vin0_consume_en_10243),
       .out_canPeek(vout_canPeek_10243),
       .out_peek(vout_peek_10243));
  assign v_10244 = v_10245 | v_10250;
  assign v_10245 = mux_10245(v_10246);
  assign v_10246 = vout_canPeek_10243 & v_10247;
  assign v_10247 = v_10248 & 1'h1;
  assign v_10248 = v_10249 | 1'h0;
  assign v_10249 = ~v_10236;
  assign v_10250 = mux_10250(v_10251);
  assign v_10251 = ~v_10246;
  pebbles_core
    pebbles_core_10252
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10253),
       .in0_consume_en(vin0_consume_en_10252),
       .out_canPeek(vout_canPeek_10252),
       .out_peek(vout_peek_10252));
  assign v_10253 = v_10254 | v_10255;
  assign v_10254 = mux_10254(v_10240);
  assign v_10255 = mux_10255(v_10256);
  assign v_10256 = ~v_10240;
  assign v_10257 = v_10258 & 1'h1;
  assign v_10258 = v_10259 & v_10260;
  assign v_10259 = ~act_10239;
  assign v_10260 = v_10261 | v_10269;
  assign v_10261 = v_10262 | v_10267;
  assign v_10262 = mux_10262(v_10263);
  assign v_10263 = v_10236 & v_10264;
  assign v_10264 = v_10265 & 1'h1;
  assign v_10265 = v_10266 | 1'h0;
  assign v_10266 = ~v_10229;
  assign v_10267 = mux_10267(v_10268);
  assign v_10268 = ~v_10263;
  assign v_10269 = ~v_10236;
  assign v_10270 = v_10271 | v_10272;
  assign v_10271 = mux_10271(v_10238);
  assign v_10272 = mux_10272(v_10257);
  assign v_10274 = v_10275 | v_10294;
  assign v_10275 = act_10276 & 1'h1;
  assign act_10276 = v_10277 | v_10283;
  assign v_10277 = v_10278 & v_10284;
  assign v_10278 = v_10279 & vout_canPeek_10289;
  assign v_10279 = ~vout_canPeek_10280;
  pebbles_core
    pebbles_core_10280
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10281),
       .in0_consume_en(vin0_consume_en_10280),
       .out_canPeek(vout_canPeek_10280),
       .out_peek(vout_peek_10280));
  assign v_10281 = v_10282 | v_10287;
  assign v_10282 = mux_10282(v_10283);
  assign v_10283 = vout_canPeek_10280 & v_10284;
  assign v_10284 = v_10285 & 1'h1;
  assign v_10285 = v_10286 | 1'h0;
  assign v_10286 = ~v_10273;
  assign v_10287 = mux_10287(v_10288);
  assign v_10288 = ~v_10283;
  pebbles_core
    pebbles_core_10289
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10290),
       .in0_consume_en(vin0_consume_en_10289),
       .out_canPeek(vout_canPeek_10289),
       .out_peek(vout_peek_10289));
  assign v_10290 = v_10291 | v_10292;
  assign v_10291 = mux_10291(v_10277);
  assign v_10292 = mux_10292(v_10293);
  assign v_10293 = ~v_10277;
  assign v_10294 = v_10295 & 1'h1;
  assign v_10295 = v_10296 & v_10297;
  assign v_10296 = ~act_10276;
  assign v_10297 = v_10298 | v_10302;
  assign v_10298 = v_10299 | v_10300;
  assign v_10299 = mux_10299(v_10233);
  assign v_10300 = mux_10300(v_10301);
  assign v_10301 = ~v_10233;
  assign v_10302 = ~v_10273;
  assign v_10303 = v_10304 | v_10305;
  assign v_10304 = mux_10304(v_10275);
  assign v_10305 = mux_10305(v_10294);
  assign v_10306 = v_10307 & 1'h1;
  assign v_10307 = v_10308 & v_10309;
  assign v_10308 = ~act_10232;
  assign v_10309 = v_10310 | v_10318;
  assign v_10310 = v_10311 | v_10316;
  assign v_10311 = mux_10311(v_10312);
  assign v_10312 = v_10229 & v_10313;
  assign v_10313 = v_10314 & 1'h1;
  assign v_10314 = v_10315 | 1'h0;
  assign v_10315 = ~v_10222;
  assign v_10316 = mux_10316(v_10317);
  assign v_10317 = ~v_10312;
  assign v_10318 = ~v_10229;
  assign v_10319 = v_10320 | v_10321;
  assign v_10320 = mux_10320(v_10231);
  assign v_10321 = mux_10321(v_10306);
  assign v_10323 = v_10324 | v_10399;
  assign v_10324 = act_10325 & 1'h1;
  assign act_10325 = v_10326 | v_10356;
  assign v_10326 = v_10327 & v_10357;
  assign v_10327 = v_10328 & v_10366;
  assign v_10328 = ~v_10329;
  assign v_10330 = v_10331 | v_10350;
  assign v_10331 = act_10332 & 1'h1;
  assign act_10332 = v_10333 | v_10339;
  assign v_10333 = v_10334 & v_10340;
  assign v_10334 = v_10335 & vout_canPeek_10345;
  assign v_10335 = ~vout_canPeek_10336;
  pebbles_core
    pebbles_core_10336
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10337),
       .in0_consume_en(vin0_consume_en_10336),
       .out_canPeek(vout_canPeek_10336),
       .out_peek(vout_peek_10336));
  assign v_10337 = v_10338 | v_10343;
  assign v_10338 = mux_10338(v_10339);
  assign v_10339 = vout_canPeek_10336 & v_10340;
  assign v_10340 = v_10341 & 1'h1;
  assign v_10341 = v_10342 | 1'h0;
  assign v_10342 = ~v_10329;
  assign v_10343 = mux_10343(v_10344);
  assign v_10344 = ~v_10339;
  pebbles_core
    pebbles_core_10345
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10346),
       .in0_consume_en(vin0_consume_en_10345),
       .out_canPeek(vout_canPeek_10345),
       .out_peek(vout_peek_10345));
  assign v_10346 = v_10347 | v_10348;
  assign v_10347 = mux_10347(v_10333);
  assign v_10348 = mux_10348(v_10349);
  assign v_10349 = ~v_10333;
  assign v_10350 = v_10351 & 1'h1;
  assign v_10351 = v_10352 & v_10353;
  assign v_10352 = ~act_10332;
  assign v_10353 = v_10354 | v_10362;
  assign v_10354 = v_10355 | v_10360;
  assign v_10355 = mux_10355(v_10356);
  assign v_10356 = v_10329 & v_10357;
  assign v_10357 = v_10358 & 1'h1;
  assign v_10358 = v_10359 | 1'h0;
  assign v_10359 = ~v_10322;
  assign v_10360 = mux_10360(v_10361);
  assign v_10361 = ~v_10356;
  assign v_10362 = ~v_10329;
  assign v_10363 = v_10364 | v_10365;
  assign v_10364 = mux_10364(v_10331);
  assign v_10365 = mux_10365(v_10350);
  assign v_10367 = v_10368 | v_10387;
  assign v_10368 = act_10369 & 1'h1;
  assign act_10369 = v_10370 | v_10376;
  assign v_10370 = v_10371 & v_10377;
  assign v_10371 = v_10372 & vout_canPeek_10382;
  assign v_10372 = ~vout_canPeek_10373;
  pebbles_core
    pebbles_core_10373
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10374),
       .in0_consume_en(vin0_consume_en_10373),
       .out_canPeek(vout_canPeek_10373),
       .out_peek(vout_peek_10373));
  assign v_10374 = v_10375 | v_10380;
  assign v_10375 = mux_10375(v_10376);
  assign v_10376 = vout_canPeek_10373 & v_10377;
  assign v_10377 = v_10378 & 1'h1;
  assign v_10378 = v_10379 | 1'h0;
  assign v_10379 = ~v_10366;
  assign v_10380 = mux_10380(v_10381);
  assign v_10381 = ~v_10376;
  pebbles_core
    pebbles_core_10382
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10383),
       .in0_consume_en(vin0_consume_en_10382),
       .out_canPeek(vout_canPeek_10382),
       .out_peek(vout_peek_10382));
  assign v_10383 = v_10384 | v_10385;
  assign v_10384 = mux_10384(v_10370);
  assign v_10385 = mux_10385(v_10386);
  assign v_10386 = ~v_10370;
  assign v_10387 = v_10388 & 1'h1;
  assign v_10388 = v_10389 & v_10390;
  assign v_10389 = ~act_10369;
  assign v_10390 = v_10391 | v_10395;
  assign v_10391 = v_10392 | v_10393;
  assign v_10392 = mux_10392(v_10326);
  assign v_10393 = mux_10393(v_10394);
  assign v_10394 = ~v_10326;
  assign v_10395 = ~v_10366;
  assign v_10396 = v_10397 | v_10398;
  assign v_10397 = mux_10397(v_10368);
  assign v_10398 = mux_10398(v_10387);
  assign v_10399 = v_10400 & 1'h1;
  assign v_10400 = v_10401 & v_10402;
  assign v_10401 = ~act_10325;
  assign v_10402 = v_10403 | v_10407;
  assign v_10403 = v_10404 | v_10405;
  assign v_10404 = mux_10404(v_10226);
  assign v_10405 = mux_10405(v_10406);
  assign v_10406 = ~v_10226;
  assign v_10407 = ~v_10322;
  assign v_10408 = v_10409 | v_10410;
  assign v_10409 = mux_10409(v_10324);
  assign v_10410 = mux_10410(v_10399);
  assign v_10411 = v_10412 & 1'h1;
  assign v_10412 = v_10413 & v_10414;
  assign v_10413 = ~act_10225;
  assign v_10414 = v_10415 | v_10423;
  assign v_10415 = v_10416 | v_10421;
  assign v_10416 = mux_10416(v_10417);
  assign v_10417 = v_10222 & v_10418;
  assign v_10418 = v_10419 & 1'h1;
  assign v_10419 = v_10420 | 1'h0;
  assign v_10420 = ~v_10215;
  assign v_10421 = mux_10421(v_10422);
  assign v_10422 = ~v_10417;
  assign v_10423 = ~v_10222;
  assign v_10424 = v_10425 | v_10426;
  assign v_10425 = mux_10425(v_10224);
  assign v_10426 = mux_10426(v_10411);
  assign v_10428 = v_10429 | v_10616;
  assign v_10429 = act_10430 & 1'h1;
  assign act_10430 = v_10431 | v_10517;
  assign v_10431 = v_10432 & v_10518;
  assign v_10432 = v_10433 & v_10527;
  assign v_10433 = ~v_10434;
  assign v_10435 = v_10436 | v_10511;
  assign v_10436 = act_10437 & 1'h1;
  assign act_10437 = v_10438 | v_10468;
  assign v_10438 = v_10439 & v_10469;
  assign v_10439 = v_10440 & v_10478;
  assign v_10440 = ~v_10441;
  assign v_10442 = v_10443 | v_10462;
  assign v_10443 = act_10444 & 1'h1;
  assign act_10444 = v_10445 | v_10451;
  assign v_10445 = v_10446 & v_10452;
  assign v_10446 = v_10447 & vout_canPeek_10457;
  assign v_10447 = ~vout_canPeek_10448;
  pebbles_core
    pebbles_core_10448
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10449),
       .in0_consume_en(vin0_consume_en_10448),
       .out_canPeek(vout_canPeek_10448),
       .out_peek(vout_peek_10448));
  assign v_10449 = v_10450 | v_10455;
  assign v_10450 = mux_10450(v_10451);
  assign v_10451 = vout_canPeek_10448 & v_10452;
  assign v_10452 = v_10453 & 1'h1;
  assign v_10453 = v_10454 | 1'h0;
  assign v_10454 = ~v_10441;
  assign v_10455 = mux_10455(v_10456);
  assign v_10456 = ~v_10451;
  pebbles_core
    pebbles_core_10457
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10458),
       .in0_consume_en(vin0_consume_en_10457),
       .out_canPeek(vout_canPeek_10457),
       .out_peek(vout_peek_10457));
  assign v_10458 = v_10459 | v_10460;
  assign v_10459 = mux_10459(v_10445);
  assign v_10460 = mux_10460(v_10461);
  assign v_10461 = ~v_10445;
  assign v_10462 = v_10463 & 1'h1;
  assign v_10463 = v_10464 & v_10465;
  assign v_10464 = ~act_10444;
  assign v_10465 = v_10466 | v_10474;
  assign v_10466 = v_10467 | v_10472;
  assign v_10467 = mux_10467(v_10468);
  assign v_10468 = v_10441 & v_10469;
  assign v_10469 = v_10470 & 1'h1;
  assign v_10470 = v_10471 | 1'h0;
  assign v_10471 = ~v_10434;
  assign v_10472 = mux_10472(v_10473);
  assign v_10473 = ~v_10468;
  assign v_10474 = ~v_10441;
  assign v_10475 = v_10476 | v_10477;
  assign v_10476 = mux_10476(v_10443);
  assign v_10477 = mux_10477(v_10462);
  assign v_10479 = v_10480 | v_10499;
  assign v_10480 = act_10481 & 1'h1;
  assign act_10481 = v_10482 | v_10488;
  assign v_10482 = v_10483 & v_10489;
  assign v_10483 = v_10484 & vout_canPeek_10494;
  assign v_10484 = ~vout_canPeek_10485;
  pebbles_core
    pebbles_core_10485
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10486),
       .in0_consume_en(vin0_consume_en_10485),
       .out_canPeek(vout_canPeek_10485),
       .out_peek(vout_peek_10485));
  assign v_10486 = v_10487 | v_10492;
  assign v_10487 = mux_10487(v_10488);
  assign v_10488 = vout_canPeek_10485 & v_10489;
  assign v_10489 = v_10490 & 1'h1;
  assign v_10490 = v_10491 | 1'h0;
  assign v_10491 = ~v_10478;
  assign v_10492 = mux_10492(v_10493);
  assign v_10493 = ~v_10488;
  pebbles_core
    pebbles_core_10494
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10495),
       .in0_consume_en(vin0_consume_en_10494),
       .out_canPeek(vout_canPeek_10494),
       .out_peek(vout_peek_10494));
  assign v_10495 = v_10496 | v_10497;
  assign v_10496 = mux_10496(v_10482);
  assign v_10497 = mux_10497(v_10498);
  assign v_10498 = ~v_10482;
  assign v_10499 = v_10500 & 1'h1;
  assign v_10500 = v_10501 & v_10502;
  assign v_10501 = ~act_10481;
  assign v_10502 = v_10503 | v_10507;
  assign v_10503 = v_10504 | v_10505;
  assign v_10504 = mux_10504(v_10438);
  assign v_10505 = mux_10505(v_10506);
  assign v_10506 = ~v_10438;
  assign v_10507 = ~v_10478;
  assign v_10508 = v_10509 | v_10510;
  assign v_10509 = mux_10509(v_10480);
  assign v_10510 = mux_10510(v_10499);
  assign v_10511 = v_10512 & 1'h1;
  assign v_10512 = v_10513 & v_10514;
  assign v_10513 = ~act_10437;
  assign v_10514 = v_10515 | v_10523;
  assign v_10515 = v_10516 | v_10521;
  assign v_10516 = mux_10516(v_10517);
  assign v_10517 = v_10434 & v_10518;
  assign v_10518 = v_10519 & 1'h1;
  assign v_10519 = v_10520 | 1'h0;
  assign v_10520 = ~v_10427;
  assign v_10521 = mux_10521(v_10522);
  assign v_10522 = ~v_10517;
  assign v_10523 = ~v_10434;
  assign v_10524 = v_10525 | v_10526;
  assign v_10525 = mux_10525(v_10436);
  assign v_10526 = mux_10526(v_10511);
  assign v_10528 = v_10529 | v_10604;
  assign v_10529 = act_10530 & 1'h1;
  assign act_10530 = v_10531 | v_10561;
  assign v_10531 = v_10532 & v_10562;
  assign v_10532 = v_10533 & v_10571;
  assign v_10533 = ~v_10534;
  assign v_10535 = v_10536 | v_10555;
  assign v_10536 = act_10537 & 1'h1;
  assign act_10537 = v_10538 | v_10544;
  assign v_10538 = v_10539 & v_10545;
  assign v_10539 = v_10540 & vout_canPeek_10550;
  assign v_10540 = ~vout_canPeek_10541;
  pebbles_core
    pebbles_core_10541
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10542),
       .in0_consume_en(vin0_consume_en_10541),
       .out_canPeek(vout_canPeek_10541),
       .out_peek(vout_peek_10541));
  assign v_10542 = v_10543 | v_10548;
  assign v_10543 = mux_10543(v_10544);
  assign v_10544 = vout_canPeek_10541 & v_10545;
  assign v_10545 = v_10546 & 1'h1;
  assign v_10546 = v_10547 | 1'h0;
  assign v_10547 = ~v_10534;
  assign v_10548 = mux_10548(v_10549);
  assign v_10549 = ~v_10544;
  pebbles_core
    pebbles_core_10550
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10551),
       .in0_consume_en(vin0_consume_en_10550),
       .out_canPeek(vout_canPeek_10550),
       .out_peek(vout_peek_10550));
  assign v_10551 = v_10552 | v_10553;
  assign v_10552 = mux_10552(v_10538);
  assign v_10553 = mux_10553(v_10554);
  assign v_10554 = ~v_10538;
  assign v_10555 = v_10556 & 1'h1;
  assign v_10556 = v_10557 & v_10558;
  assign v_10557 = ~act_10537;
  assign v_10558 = v_10559 | v_10567;
  assign v_10559 = v_10560 | v_10565;
  assign v_10560 = mux_10560(v_10561);
  assign v_10561 = v_10534 & v_10562;
  assign v_10562 = v_10563 & 1'h1;
  assign v_10563 = v_10564 | 1'h0;
  assign v_10564 = ~v_10527;
  assign v_10565 = mux_10565(v_10566);
  assign v_10566 = ~v_10561;
  assign v_10567 = ~v_10534;
  assign v_10568 = v_10569 | v_10570;
  assign v_10569 = mux_10569(v_10536);
  assign v_10570 = mux_10570(v_10555);
  assign v_10572 = v_10573 | v_10592;
  assign v_10573 = act_10574 & 1'h1;
  assign act_10574 = v_10575 | v_10581;
  assign v_10575 = v_10576 & v_10582;
  assign v_10576 = v_10577 & vout_canPeek_10587;
  assign v_10577 = ~vout_canPeek_10578;
  pebbles_core
    pebbles_core_10578
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10579),
       .in0_consume_en(vin0_consume_en_10578),
       .out_canPeek(vout_canPeek_10578),
       .out_peek(vout_peek_10578));
  assign v_10579 = v_10580 | v_10585;
  assign v_10580 = mux_10580(v_10581);
  assign v_10581 = vout_canPeek_10578 & v_10582;
  assign v_10582 = v_10583 & 1'h1;
  assign v_10583 = v_10584 | 1'h0;
  assign v_10584 = ~v_10571;
  assign v_10585 = mux_10585(v_10586);
  assign v_10586 = ~v_10581;
  pebbles_core
    pebbles_core_10587
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10588),
       .in0_consume_en(vin0_consume_en_10587),
       .out_canPeek(vout_canPeek_10587),
       .out_peek(vout_peek_10587));
  assign v_10588 = v_10589 | v_10590;
  assign v_10589 = mux_10589(v_10575);
  assign v_10590 = mux_10590(v_10591);
  assign v_10591 = ~v_10575;
  assign v_10592 = v_10593 & 1'h1;
  assign v_10593 = v_10594 & v_10595;
  assign v_10594 = ~act_10574;
  assign v_10595 = v_10596 | v_10600;
  assign v_10596 = v_10597 | v_10598;
  assign v_10597 = mux_10597(v_10531);
  assign v_10598 = mux_10598(v_10599);
  assign v_10599 = ~v_10531;
  assign v_10600 = ~v_10571;
  assign v_10601 = v_10602 | v_10603;
  assign v_10602 = mux_10602(v_10573);
  assign v_10603 = mux_10603(v_10592);
  assign v_10604 = v_10605 & 1'h1;
  assign v_10605 = v_10606 & v_10607;
  assign v_10606 = ~act_10530;
  assign v_10607 = v_10608 | v_10612;
  assign v_10608 = v_10609 | v_10610;
  assign v_10609 = mux_10609(v_10431);
  assign v_10610 = mux_10610(v_10611);
  assign v_10611 = ~v_10431;
  assign v_10612 = ~v_10527;
  assign v_10613 = v_10614 | v_10615;
  assign v_10614 = mux_10614(v_10529);
  assign v_10615 = mux_10615(v_10604);
  assign v_10616 = v_10617 & 1'h1;
  assign v_10617 = v_10618 & v_10619;
  assign v_10618 = ~act_10430;
  assign v_10619 = v_10620 | v_10624;
  assign v_10620 = v_10621 | v_10622;
  assign v_10621 = mux_10621(v_10219);
  assign v_10622 = mux_10622(v_10623);
  assign v_10623 = ~v_10219;
  assign v_10624 = ~v_10427;
  assign v_10625 = v_10626 | v_10627;
  assign v_10626 = mux_10626(v_10429);
  assign v_10627 = mux_10627(v_10616);
  assign v_10628 = v_10629 & 1'h1;
  assign v_10629 = v_10630 & v_10631;
  assign v_10630 = ~act_10218;
  assign v_10631 = v_10632 | v_10636;
  assign v_10632 = v_10633 | v_10634;
  assign v_10633 = mux_10633(v_9783);
  assign v_10634 = mux_10634(v_10635);
  assign v_10635 = ~v_9783;
  assign v_10636 = ~v_10215;
  assign v_10637 = v_10638 | v_10639;
  assign v_10638 = mux_10638(v_10217);
  assign v_10639 = mux_10639(v_10628);
  assign v_10640 = v_10641 & 1'h1;
  assign v_10641 = v_10642 & v_10643;
  assign v_10642 = ~act_9782;
  assign v_10643 = v_10644 | v_10652;
  assign v_10644 = v_10645 | v_10650;
  assign v_10645 = mux_10645(v_10646);
  assign v_10646 = v_9779 & v_10647;
  assign v_10647 = v_10648 & 1'h1;
  assign v_10648 = v_10649 | 1'h0;
  assign v_10649 = ~v_9772;
  assign v_10650 = mux_10650(v_10651);
  assign v_10651 = ~v_10646;
  assign v_10652 = ~v_9779;
  assign v_10653 = v_10654 | v_10655;
  assign v_10654 = mux_10654(v_9781);
  assign v_10655 = mux_10655(v_10640);
  assign v_10657 = v_10658 | v_11517;
  assign v_10658 = act_10659 & 1'h1;
  assign act_10659 = v_10660 | v_11082;
  assign v_10660 = v_10661 & v_11083;
  assign v_10661 = v_10662 & v_11092;
  assign v_10662 = ~v_10663;
  assign v_10664 = v_10665 | v_11076;
  assign v_10665 = act_10666 & 1'h1;
  assign act_10666 = v_10667 | v_10865;
  assign v_10667 = v_10668 & v_10866;
  assign v_10668 = v_10669 & v_10875;
  assign v_10669 = ~v_10670;
  assign v_10671 = v_10672 | v_10859;
  assign v_10672 = act_10673 & 1'h1;
  assign act_10673 = v_10674 | v_10760;
  assign v_10674 = v_10675 & v_10761;
  assign v_10675 = v_10676 & v_10770;
  assign v_10676 = ~v_10677;
  assign v_10678 = v_10679 | v_10754;
  assign v_10679 = act_10680 & 1'h1;
  assign act_10680 = v_10681 | v_10711;
  assign v_10681 = v_10682 & v_10712;
  assign v_10682 = v_10683 & v_10721;
  assign v_10683 = ~v_10684;
  assign v_10685 = v_10686 | v_10705;
  assign v_10686 = act_10687 & 1'h1;
  assign act_10687 = v_10688 | v_10694;
  assign v_10688 = v_10689 & v_10695;
  assign v_10689 = v_10690 & vout_canPeek_10700;
  assign v_10690 = ~vout_canPeek_10691;
  pebbles_core
    pebbles_core_10691
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10692),
       .in0_consume_en(vin0_consume_en_10691),
       .out_canPeek(vout_canPeek_10691),
       .out_peek(vout_peek_10691));
  assign v_10692 = v_10693 | v_10698;
  assign v_10693 = mux_10693(v_10694);
  assign v_10694 = vout_canPeek_10691 & v_10695;
  assign v_10695 = v_10696 & 1'h1;
  assign v_10696 = v_10697 | 1'h0;
  assign v_10697 = ~v_10684;
  assign v_10698 = mux_10698(v_10699);
  assign v_10699 = ~v_10694;
  pebbles_core
    pebbles_core_10700
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10701),
       .in0_consume_en(vin0_consume_en_10700),
       .out_canPeek(vout_canPeek_10700),
       .out_peek(vout_peek_10700));
  assign v_10701 = v_10702 | v_10703;
  assign v_10702 = mux_10702(v_10688);
  assign v_10703 = mux_10703(v_10704);
  assign v_10704 = ~v_10688;
  assign v_10705 = v_10706 & 1'h1;
  assign v_10706 = v_10707 & v_10708;
  assign v_10707 = ~act_10687;
  assign v_10708 = v_10709 | v_10717;
  assign v_10709 = v_10710 | v_10715;
  assign v_10710 = mux_10710(v_10711);
  assign v_10711 = v_10684 & v_10712;
  assign v_10712 = v_10713 & 1'h1;
  assign v_10713 = v_10714 | 1'h0;
  assign v_10714 = ~v_10677;
  assign v_10715 = mux_10715(v_10716);
  assign v_10716 = ~v_10711;
  assign v_10717 = ~v_10684;
  assign v_10718 = v_10719 | v_10720;
  assign v_10719 = mux_10719(v_10686);
  assign v_10720 = mux_10720(v_10705);
  assign v_10722 = v_10723 | v_10742;
  assign v_10723 = act_10724 & 1'h1;
  assign act_10724 = v_10725 | v_10731;
  assign v_10725 = v_10726 & v_10732;
  assign v_10726 = v_10727 & vout_canPeek_10737;
  assign v_10727 = ~vout_canPeek_10728;
  pebbles_core
    pebbles_core_10728
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10729),
       .in0_consume_en(vin0_consume_en_10728),
       .out_canPeek(vout_canPeek_10728),
       .out_peek(vout_peek_10728));
  assign v_10729 = v_10730 | v_10735;
  assign v_10730 = mux_10730(v_10731);
  assign v_10731 = vout_canPeek_10728 & v_10732;
  assign v_10732 = v_10733 & 1'h1;
  assign v_10733 = v_10734 | 1'h0;
  assign v_10734 = ~v_10721;
  assign v_10735 = mux_10735(v_10736);
  assign v_10736 = ~v_10731;
  pebbles_core
    pebbles_core_10737
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10738),
       .in0_consume_en(vin0_consume_en_10737),
       .out_canPeek(vout_canPeek_10737),
       .out_peek(vout_peek_10737));
  assign v_10738 = v_10739 | v_10740;
  assign v_10739 = mux_10739(v_10725);
  assign v_10740 = mux_10740(v_10741);
  assign v_10741 = ~v_10725;
  assign v_10742 = v_10743 & 1'h1;
  assign v_10743 = v_10744 & v_10745;
  assign v_10744 = ~act_10724;
  assign v_10745 = v_10746 | v_10750;
  assign v_10746 = v_10747 | v_10748;
  assign v_10747 = mux_10747(v_10681);
  assign v_10748 = mux_10748(v_10749);
  assign v_10749 = ~v_10681;
  assign v_10750 = ~v_10721;
  assign v_10751 = v_10752 | v_10753;
  assign v_10752 = mux_10752(v_10723);
  assign v_10753 = mux_10753(v_10742);
  assign v_10754 = v_10755 & 1'h1;
  assign v_10755 = v_10756 & v_10757;
  assign v_10756 = ~act_10680;
  assign v_10757 = v_10758 | v_10766;
  assign v_10758 = v_10759 | v_10764;
  assign v_10759 = mux_10759(v_10760);
  assign v_10760 = v_10677 & v_10761;
  assign v_10761 = v_10762 & 1'h1;
  assign v_10762 = v_10763 | 1'h0;
  assign v_10763 = ~v_10670;
  assign v_10764 = mux_10764(v_10765);
  assign v_10765 = ~v_10760;
  assign v_10766 = ~v_10677;
  assign v_10767 = v_10768 | v_10769;
  assign v_10768 = mux_10768(v_10679);
  assign v_10769 = mux_10769(v_10754);
  assign v_10771 = v_10772 | v_10847;
  assign v_10772 = act_10773 & 1'h1;
  assign act_10773 = v_10774 | v_10804;
  assign v_10774 = v_10775 & v_10805;
  assign v_10775 = v_10776 & v_10814;
  assign v_10776 = ~v_10777;
  assign v_10778 = v_10779 | v_10798;
  assign v_10779 = act_10780 & 1'h1;
  assign act_10780 = v_10781 | v_10787;
  assign v_10781 = v_10782 & v_10788;
  assign v_10782 = v_10783 & vout_canPeek_10793;
  assign v_10783 = ~vout_canPeek_10784;
  pebbles_core
    pebbles_core_10784
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10785),
       .in0_consume_en(vin0_consume_en_10784),
       .out_canPeek(vout_canPeek_10784),
       .out_peek(vout_peek_10784));
  assign v_10785 = v_10786 | v_10791;
  assign v_10786 = mux_10786(v_10787);
  assign v_10787 = vout_canPeek_10784 & v_10788;
  assign v_10788 = v_10789 & 1'h1;
  assign v_10789 = v_10790 | 1'h0;
  assign v_10790 = ~v_10777;
  assign v_10791 = mux_10791(v_10792);
  assign v_10792 = ~v_10787;
  pebbles_core
    pebbles_core_10793
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10794),
       .in0_consume_en(vin0_consume_en_10793),
       .out_canPeek(vout_canPeek_10793),
       .out_peek(vout_peek_10793));
  assign v_10794 = v_10795 | v_10796;
  assign v_10795 = mux_10795(v_10781);
  assign v_10796 = mux_10796(v_10797);
  assign v_10797 = ~v_10781;
  assign v_10798 = v_10799 & 1'h1;
  assign v_10799 = v_10800 & v_10801;
  assign v_10800 = ~act_10780;
  assign v_10801 = v_10802 | v_10810;
  assign v_10802 = v_10803 | v_10808;
  assign v_10803 = mux_10803(v_10804);
  assign v_10804 = v_10777 & v_10805;
  assign v_10805 = v_10806 & 1'h1;
  assign v_10806 = v_10807 | 1'h0;
  assign v_10807 = ~v_10770;
  assign v_10808 = mux_10808(v_10809);
  assign v_10809 = ~v_10804;
  assign v_10810 = ~v_10777;
  assign v_10811 = v_10812 | v_10813;
  assign v_10812 = mux_10812(v_10779);
  assign v_10813 = mux_10813(v_10798);
  assign v_10815 = v_10816 | v_10835;
  assign v_10816 = act_10817 & 1'h1;
  assign act_10817 = v_10818 | v_10824;
  assign v_10818 = v_10819 & v_10825;
  assign v_10819 = v_10820 & vout_canPeek_10830;
  assign v_10820 = ~vout_canPeek_10821;
  pebbles_core
    pebbles_core_10821
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10822),
       .in0_consume_en(vin0_consume_en_10821),
       .out_canPeek(vout_canPeek_10821),
       .out_peek(vout_peek_10821));
  assign v_10822 = v_10823 | v_10828;
  assign v_10823 = mux_10823(v_10824);
  assign v_10824 = vout_canPeek_10821 & v_10825;
  assign v_10825 = v_10826 & 1'h1;
  assign v_10826 = v_10827 | 1'h0;
  assign v_10827 = ~v_10814;
  assign v_10828 = mux_10828(v_10829);
  assign v_10829 = ~v_10824;
  pebbles_core
    pebbles_core_10830
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10831),
       .in0_consume_en(vin0_consume_en_10830),
       .out_canPeek(vout_canPeek_10830),
       .out_peek(vout_peek_10830));
  assign v_10831 = v_10832 | v_10833;
  assign v_10832 = mux_10832(v_10818);
  assign v_10833 = mux_10833(v_10834);
  assign v_10834 = ~v_10818;
  assign v_10835 = v_10836 & 1'h1;
  assign v_10836 = v_10837 & v_10838;
  assign v_10837 = ~act_10817;
  assign v_10838 = v_10839 | v_10843;
  assign v_10839 = v_10840 | v_10841;
  assign v_10840 = mux_10840(v_10774);
  assign v_10841 = mux_10841(v_10842);
  assign v_10842 = ~v_10774;
  assign v_10843 = ~v_10814;
  assign v_10844 = v_10845 | v_10846;
  assign v_10845 = mux_10845(v_10816);
  assign v_10846 = mux_10846(v_10835);
  assign v_10847 = v_10848 & 1'h1;
  assign v_10848 = v_10849 & v_10850;
  assign v_10849 = ~act_10773;
  assign v_10850 = v_10851 | v_10855;
  assign v_10851 = v_10852 | v_10853;
  assign v_10852 = mux_10852(v_10674);
  assign v_10853 = mux_10853(v_10854);
  assign v_10854 = ~v_10674;
  assign v_10855 = ~v_10770;
  assign v_10856 = v_10857 | v_10858;
  assign v_10857 = mux_10857(v_10772);
  assign v_10858 = mux_10858(v_10847);
  assign v_10859 = v_10860 & 1'h1;
  assign v_10860 = v_10861 & v_10862;
  assign v_10861 = ~act_10673;
  assign v_10862 = v_10863 | v_10871;
  assign v_10863 = v_10864 | v_10869;
  assign v_10864 = mux_10864(v_10865);
  assign v_10865 = v_10670 & v_10866;
  assign v_10866 = v_10867 & 1'h1;
  assign v_10867 = v_10868 | 1'h0;
  assign v_10868 = ~v_10663;
  assign v_10869 = mux_10869(v_10870);
  assign v_10870 = ~v_10865;
  assign v_10871 = ~v_10670;
  assign v_10872 = v_10873 | v_10874;
  assign v_10873 = mux_10873(v_10672);
  assign v_10874 = mux_10874(v_10859);
  assign v_10876 = v_10877 | v_11064;
  assign v_10877 = act_10878 & 1'h1;
  assign act_10878 = v_10879 | v_10965;
  assign v_10879 = v_10880 & v_10966;
  assign v_10880 = v_10881 & v_10975;
  assign v_10881 = ~v_10882;
  assign v_10883 = v_10884 | v_10959;
  assign v_10884 = act_10885 & 1'h1;
  assign act_10885 = v_10886 | v_10916;
  assign v_10886 = v_10887 & v_10917;
  assign v_10887 = v_10888 & v_10926;
  assign v_10888 = ~v_10889;
  assign v_10890 = v_10891 | v_10910;
  assign v_10891 = act_10892 & 1'h1;
  assign act_10892 = v_10893 | v_10899;
  assign v_10893 = v_10894 & v_10900;
  assign v_10894 = v_10895 & vout_canPeek_10905;
  assign v_10895 = ~vout_canPeek_10896;
  pebbles_core
    pebbles_core_10896
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10897),
       .in0_consume_en(vin0_consume_en_10896),
       .out_canPeek(vout_canPeek_10896),
       .out_peek(vout_peek_10896));
  assign v_10897 = v_10898 | v_10903;
  assign v_10898 = mux_10898(v_10899);
  assign v_10899 = vout_canPeek_10896 & v_10900;
  assign v_10900 = v_10901 & 1'h1;
  assign v_10901 = v_10902 | 1'h0;
  assign v_10902 = ~v_10889;
  assign v_10903 = mux_10903(v_10904);
  assign v_10904 = ~v_10899;
  pebbles_core
    pebbles_core_10905
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10906),
       .in0_consume_en(vin0_consume_en_10905),
       .out_canPeek(vout_canPeek_10905),
       .out_peek(vout_peek_10905));
  assign v_10906 = v_10907 | v_10908;
  assign v_10907 = mux_10907(v_10893);
  assign v_10908 = mux_10908(v_10909);
  assign v_10909 = ~v_10893;
  assign v_10910 = v_10911 & 1'h1;
  assign v_10911 = v_10912 & v_10913;
  assign v_10912 = ~act_10892;
  assign v_10913 = v_10914 | v_10922;
  assign v_10914 = v_10915 | v_10920;
  assign v_10915 = mux_10915(v_10916);
  assign v_10916 = v_10889 & v_10917;
  assign v_10917 = v_10918 & 1'h1;
  assign v_10918 = v_10919 | 1'h0;
  assign v_10919 = ~v_10882;
  assign v_10920 = mux_10920(v_10921);
  assign v_10921 = ~v_10916;
  assign v_10922 = ~v_10889;
  assign v_10923 = v_10924 | v_10925;
  assign v_10924 = mux_10924(v_10891);
  assign v_10925 = mux_10925(v_10910);
  assign v_10927 = v_10928 | v_10947;
  assign v_10928 = act_10929 & 1'h1;
  assign act_10929 = v_10930 | v_10936;
  assign v_10930 = v_10931 & v_10937;
  assign v_10931 = v_10932 & vout_canPeek_10942;
  assign v_10932 = ~vout_canPeek_10933;
  pebbles_core
    pebbles_core_10933
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10934),
       .in0_consume_en(vin0_consume_en_10933),
       .out_canPeek(vout_canPeek_10933),
       .out_peek(vout_peek_10933));
  assign v_10934 = v_10935 | v_10940;
  assign v_10935 = mux_10935(v_10936);
  assign v_10936 = vout_canPeek_10933 & v_10937;
  assign v_10937 = v_10938 & 1'h1;
  assign v_10938 = v_10939 | 1'h0;
  assign v_10939 = ~v_10926;
  assign v_10940 = mux_10940(v_10941);
  assign v_10941 = ~v_10936;
  pebbles_core
    pebbles_core_10942
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10943),
       .in0_consume_en(vin0_consume_en_10942),
       .out_canPeek(vout_canPeek_10942),
       .out_peek(vout_peek_10942));
  assign v_10943 = v_10944 | v_10945;
  assign v_10944 = mux_10944(v_10930);
  assign v_10945 = mux_10945(v_10946);
  assign v_10946 = ~v_10930;
  assign v_10947 = v_10948 & 1'h1;
  assign v_10948 = v_10949 & v_10950;
  assign v_10949 = ~act_10929;
  assign v_10950 = v_10951 | v_10955;
  assign v_10951 = v_10952 | v_10953;
  assign v_10952 = mux_10952(v_10886);
  assign v_10953 = mux_10953(v_10954);
  assign v_10954 = ~v_10886;
  assign v_10955 = ~v_10926;
  assign v_10956 = v_10957 | v_10958;
  assign v_10957 = mux_10957(v_10928);
  assign v_10958 = mux_10958(v_10947);
  assign v_10959 = v_10960 & 1'h1;
  assign v_10960 = v_10961 & v_10962;
  assign v_10961 = ~act_10885;
  assign v_10962 = v_10963 | v_10971;
  assign v_10963 = v_10964 | v_10969;
  assign v_10964 = mux_10964(v_10965);
  assign v_10965 = v_10882 & v_10966;
  assign v_10966 = v_10967 & 1'h1;
  assign v_10967 = v_10968 | 1'h0;
  assign v_10968 = ~v_10875;
  assign v_10969 = mux_10969(v_10970);
  assign v_10970 = ~v_10965;
  assign v_10971 = ~v_10882;
  assign v_10972 = v_10973 | v_10974;
  assign v_10973 = mux_10973(v_10884);
  assign v_10974 = mux_10974(v_10959);
  assign v_10976 = v_10977 | v_11052;
  assign v_10977 = act_10978 & 1'h1;
  assign act_10978 = v_10979 | v_11009;
  assign v_10979 = v_10980 & v_11010;
  assign v_10980 = v_10981 & v_11019;
  assign v_10981 = ~v_10982;
  assign v_10983 = v_10984 | v_11003;
  assign v_10984 = act_10985 & 1'h1;
  assign act_10985 = v_10986 | v_10992;
  assign v_10986 = v_10987 & v_10993;
  assign v_10987 = v_10988 & vout_canPeek_10998;
  assign v_10988 = ~vout_canPeek_10989;
  pebbles_core
    pebbles_core_10989
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10990),
       .in0_consume_en(vin0_consume_en_10989),
       .out_canPeek(vout_canPeek_10989),
       .out_peek(vout_peek_10989));
  assign v_10990 = v_10991 | v_10996;
  assign v_10991 = mux_10991(v_10992);
  assign v_10992 = vout_canPeek_10989 & v_10993;
  assign v_10993 = v_10994 & 1'h1;
  assign v_10994 = v_10995 | 1'h0;
  assign v_10995 = ~v_10982;
  assign v_10996 = mux_10996(v_10997);
  assign v_10997 = ~v_10992;
  pebbles_core
    pebbles_core_10998
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_10999),
       .in0_consume_en(vin0_consume_en_10998),
       .out_canPeek(vout_canPeek_10998),
       .out_peek(vout_peek_10998));
  assign v_10999 = v_11000 | v_11001;
  assign v_11000 = mux_11000(v_10986);
  assign v_11001 = mux_11001(v_11002);
  assign v_11002 = ~v_10986;
  assign v_11003 = v_11004 & 1'h1;
  assign v_11004 = v_11005 & v_11006;
  assign v_11005 = ~act_10985;
  assign v_11006 = v_11007 | v_11015;
  assign v_11007 = v_11008 | v_11013;
  assign v_11008 = mux_11008(v_11009);
  assign v_11009 = v_10982 & v_11010;
  assign v_11010 = v_11011 & 1'h1;
  assign v_11011 = v_11012 | 1'h0;
  assign v_11012 = ~v_10975;
  assign v_11013 = mux_11013(v_11014);
  assign v_11014 = ~v_11009;
  assign v_11015 = ~v_10982;
  assign v_11016 = v_11017 | v_11018;
  assign v_11017 = mux_11017(v_10984);
  assign v_11018 = mux_11018(v_11003);
  assign v_11020 = v_11021 | v_11040;
  assign v_11021 = act_11022 & 1'h1;
  assign act_11022 = v_11023 | v_11029;
  assign v_11023 = v_11024 & v_11030;
  assign v_11024 = v_11025 & vout_canPeek_11035;
  assign v_11025 = ~vout_canPeek_11026;
  pebbles_core
    pebbles_core_11026
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11027),
       .in0_consume_en(vin0_consume_en_11026),
       .out_canPeek(vout_canPeek_11026),
       .out_peek(vout_peek_11026));
  assign v_11027 = v_11028 | v_11033;
  assign v_11028 = mux_11028(v_11029);
  assign v_11029 = vout_canPeek_11026 & v_11030;
  assign v_11030 = v_11031 & 1'h1;
  assign v_11031 = v_11032 | 1'h0;
  assign v_11032 = ~v_11019;
  assign v_11033 = mux_11033(v_11034);
  assign v_11034 = ~v_11029;
  pebbles_core
    pebbles_core_11035
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11036),
       .in0_consume_en(vin0_consume_en_11035),
       .out_canPeek(vout_canPeek_11035),
       .out_peek(vout_peek_11035));
  assign v_11036 = v_11037 | v_11038;
  assign v_11037 = mux_11037(v_11023);
  assign v_11038 = mux_11038(v_11039);
  assign v_11039 = ~v_11023;
  assign v_11040 = v_11041 & 1'h1;
  assign v_11041 = v_11042 & v_11043;
  assign v_11042 = ~act_11022;
  assign v_11043 = v_11044 | v_11048;
  assign v_11044 = v_11045 | v_11046;
  assign v_11045 = mux_11045(v_10979);
  assign v_11046 = mux_11046(v_11047);
  assign v_11047 = ~v_10979;
  assign v_11048 = ~v_11019;
  assign v_11049 = v_11050 | v_11051;
  assign v_11050 = mux_11050(v_11021);
  assign v_11051 = mux_11051(v_11040);
  assign v_11052 = v_11053 & 1'h1;
  assign v_11053 = v_11054 & v_11055;
  assign v_11054 = ~act_10978;
  assign v_11055 = v_11056 | v_11060;
  assign v_11056 = v_11057 | v_11058;
  assign v_11057 = mux_11057(v_10879);
  assign v_11058 = mux_11058(v_11059);
  assign v_11059 = ~v_10879;
  assign v_11060 = ~v_10975;
  assign v_11061 = v_11062 | v_11063;
  assign v_11062 = mux_11062(v_10977);
  assign v_11063 = mux_11063(v_11052);
  assign v_11064 = v_11065 & 1'h1;
  assign v_11065 = v_11066 & v_11067;
  assign v_11066 = ~act_10878;
  assign v_11067 = v_11068 | v_11072;
  assign v_11068 = v_11069 | v_11070;
  assign v_11069 = mux_11069(v_10667);
  assign v_11070 = mux_11070(v_11071);
  assign v_11071 = ~v_10667;
  assign v_11072 = ~v_10875;
  assign v_11073 = v_11074 | v_11075;
  assign v_11074 = mux_11074(v_10877);
  assign v_11075 = mux_11075(v_11064);
  assign v_11076 = v_11077 & 1'h1;
  assign v_11077 = v_11078 & v_11079;
  assign v_11078 = ~act_10666;
  assign v_11079 = v_11080 | v_11088;
  assign v_11080 = v_11081 | v_11086;
  assign v_11081 = mux_11081(v_11082);
  assign v_11082 = v_10663 & v_11083;
  assign v_11083 = v_11084 & 1'h1;
  assign v_11084 = v_11085 | 1'h0;
  assign v_11085 = ~v_10656;
  assign v_11086 = mux_11086(v_11087);
  assign v_11087 = ~v_11082;
  assign v_11088 = ~v_10663;
  assign v_11089 = v_11090 | v_11091;
  assign v_11090 = mux_11090(v_10665);
  assign v_11091 = mux_11091(v_11076);
  assign v_11093 = v_11094 | v_11505;
  assign v_11094 = act_11095 & 1'h1;
  assign act_11095 = v_11096 | v_11294;
  assign v_11096 = v_11097 & v_11295;
  assign v_11097 = v_11098 & v_11304;
  assign v_11098 = ~v_11099;
  assign v_11100 = v_11101 | v_11288;
  assign v_11101 = act_11102 & 1'h1;
  assign act_11102 = v_11103 | v_11189;
  assign v_11103 = v_11104 & v_11190;
  assign v_11104 = v_11105 & v_11199;
  assign v_11105 = ~v_11106;
  assign v_11107 = v_11108 | v_11183;
  assign v_11108 = act_11109 & 1'h1;
  assign act_11109 = v_11110 | v_11140;
  assign v_11110 = v_11111 & v_11141;
  assign v_11111 = v_11112 & v_11150;
  assign v_11112 = ~v_11113;
  assign v_11114 = v_11115 | v_11134;
  assign v_11115 = act_11116 & 1'h1;
  assign act_11116 = v_11117 | v_11123;
  assign v_11117 = v_11118 & v_11124;
  assign v_11118 = v_11119 & vout_canPeek_11129;
  assign v_11119 = ~vout_canPeek_11120;
  pebbles_core
    pebbles_core_11120
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11121),
       .in0_consume_en(vin0_consume_en_11120),
       .out_canPeek(vout_canPeek_11120),
       .out_peek(vout_peek_11120));
  assign v_11121 = v_11122 | v_11127;
  assign v_11122 = mux_11122(v_11123);
  assign v_11123 = vout_canPeek_11120 & v_11124;
  assign v_11124 = v_11125 & 1'h1;
  assign v_11125 = v_11126 | 1'h0;
  assign v_11126 = ~v_11113;
  assign v_11127 = mux_11127(v_11128);
  assign v_11128 = ~v_11123;
  pebbles_core
    pebbles_core_11129
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11130),
       .in0_consume_en(vin0_consume_en_11129),
       .out_canPeek(vout_canPeek_11129),
       .out_peek(vout_peek_11129));
  assign v_11130 = v_11131 | v_11132;
  assign v_11131 = mux_11131(v_11117);
  assign v_11132 = mux_11132(v_11133);
  assign v_11133 = ~v_11117;
  assign v_11134 = v_11135 & 1'h1;
  assign v_11135 = v_11136 & v_11137;
  assign v_11136 = ~act_11116;
  assign v_11137 = v_11138 | v_11146;
  assign v_11138 = v_11139 | v_11144;
  assign v_11139 = mux_11139(v_11140);
  assign v_11140 = v_11113 & v_11141;
  assign v_11141 = v_11142 & 1'h1;
  assign v_11142 = v_11143 | 1'h0;
  assign v_11143 = ~v_11106;
  assign v_11144 = mux_11144(v_11145);
  assign v_11145 = ~v_11140;
  assign v_11146 = ~v_11113;
  assign v_11147 = v_11148 | v_11149;
  assign v_11148 = mux_11148(v_11115);
  assign v_11149 = mux_11149(v_11134);
  assign v_11151 = v_11152 | v_11171;
  assign v_11152 = act_11153 & 1'h1;
  assign act_11153 = v_11154 | v_11160;
  assign v_11154 = v_11155 & v_11161;
  assign v_11155 = v_11156 & vout_canPeek_11166;
  assign v_11156 = ~vout_canPeek_11157;
  pebbles_core
    pebbles_core_11157
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11158),
       .in0_consume_en(vin0_consume_en_11157),
       .out_canPeek(vout_canPeek_11157),
       .out_peek(vout_peek_11157));
  assign v_11158 = v_11159 | v_11164;
  assign v_11159 = mux_11159(v_11160);
  assign v_11160 = vout_canPeek_11157 & v_11161;
  assign v_11161 = v_11162 & 1'h1;
  assign v_11162 = v_11163 | 1'h0;
  assign v_11163 = ~v_11150;
  assign v_11164 = mux_11164(v_11165);
  assign v_11165 = ~v_11160;
  pebbles_core
    pebbles_core_11166
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11167),
       .in0_consume_en(vin0_consume_en_11166),
       .out_canPeek(vout_canPeek_11166),
       .out_peek(vout_peek_11166));
  assign v_11167 = v_11168 | v_11169;
  assign v_11168 = mux_11168(v_11154);
  assign v_11169 = mux_11169(v_11170);
  assign v_11170 = ~v_11154;
  assign v_11171 = v_11172 & 1'h1;
  assign v_11172 = v_11173 & v_11174;
  assign v_11173 = ~act_11153;
  assign v_11174 = v_11175 | v_11179;
  assign v_11175 = v_11176 | v_11177;
  assign v_11176 = mux_11176(v_11110);
  assign v_11177 = mux_11177(v_11178);
  assign v_11178 = ~v_11110;
  assign v_11179 = ~v_11150;
  assign v_11180 = v_11181 | v_11182;
  assign v_11181 = mux_11181(v_11152);
  assign v_11182 = mux_11182(v_11171);
  assign v_11183 = v_11184 & 1'h1;
  assign v_11184 = v_11185 & v_11186;
  assign v_11185 = ~act_11109;
  assign v_11186 = v_11187 | v_11195;
  assign v_11187 = v_11188 | v_11193;
  assign v_11188 = mux_11188(v_11189);
  assign v_11189 = v_11106 & v_11190;
  assign v_11190 = v_11191 & 1'h1;
  assign v_11191 = v_11192 | 1'h0;
  assign v_11192 = ~v_11099;
  assign v_11193 = mux_11193(v_11194);
  assign v_11194 = ~v_11189;
  assign v_11195 = ~v_11106;
  assign v_11196 = v_11197 | v_11198;
  assign v_11197 = mux_11197(v_11108);
  assign v_11198 = mux_11198(v_11183);
  assign v_11200 = v_11201 | v_11276;
  assign v_11201 = act_11202 & 1'h1;
  assign act_11202 = v_11203 | v_11233;
  assign v_11203 = v_11204 & v_11234;
  assign v_11204 = v_11205 & v_11243;
  assign v_11205 = ~v_11206;
  assign v_11207 = v_11208 | v_11227;
  assign v_11208 = act_11209 & 1'h1;
  assign act_11209 = v_11210 | v_11216;
  assign v_11210 = v_11211 & v_11217;
  assign v_11211 = v_11212 & vout_canPeek_11222;
  assign v_11212 = ~vout_canPeek_11213;
  pebbles_core
    pebbles_core_11213
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11214),
       .in0_consume_en(vin0_consume_en_11213),
       .out_canPeek(vout_canPeek_11213),
       .out_peek(vout_peek_11213));
  assign v_11214 = v_11215 | v_11220;
  assign v_11215 = mux_11215(v_11216);
  assign v_11216 = vout_canPeek_11213 & v_11217;
  assign v_11217 = v_11218 & 1'h1;
  assign v_11218 = v_11219 | 1'h0;
  assign v_11219 = ~v_11206;
  assign v_11220 = mux_11220(v_11221);
  assign v_11221 = ~v_11216;
  pebbles_core
    pebbles_core_11222
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11223),
       .in0_consume_en(vin0_consume_en_11222),
       .out_canPeek(vout_canPeek_11222),
       .out_peek(vout_peek_11222));
  assign v_11223 = v_11224 | v_11225;
  assign v_11224 = mux_11224(v_11210);
  assign v_11225 = mux_11225(v_11226);
  assign v_11226 = ~v_11210;
  assign v_11227 = v_11228 & 1'h1;
  assign v_11228 = v_11229 & v_11230;
  assign v_11229 = ~act_11209;
  assign v_11230 = v_11231 | v_11239;
  assign v_11231 = v_11232 | v_11237;
  assign v_11232 = mux_11232(v_11233);
  assign v_11233 = v_11206 & v_11234;
  assign v_11234 = v_11235 & 1'h1;
  assign v_11235 = v_11236 | 1'h0;
  assign v_11236 = ~v_11199;
  assign v_11237 = mux_11237(v_11238);
  assign v_11238 = ~v_11233;
  assign v_11239 = ~v_11206;
  assign v_11240 = v_11241 | v_11242;
  assign v_11241 = mux_11241(v_11208);
  assign v_11242 = mux_11242(v_11227);
  assign v_11244 = v_11245 | v_11264;
  assign v_11245 = act_11246 & 1'h1;
  assign act_11246 = v_11247 | v_11253;
  assign v_11247 = v_11248 & v_11254;
  assign v_11248 = v_11249 & vout_canPeek_11259;
  assign v_11249 = ~vout_canPeek_11250;
  pebbles_core
    pebbles_core_11250
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11251),
       .in0_consume_en(vin0_consume_en_11250),
       .out_canPeek(vout_canPeek_11250),
       .out_peek(vout_peek_11250));
  assign v_11251 = v_11252 | v_11257;
  assign v_11252 = mux_11252(v_11253);
  assign v_11253 = vout_canPeek_11250 & v_11254;
  assign v_11254 = v_11255 & 1'h1;
  assign v_11255 = v_11256 | 1'h0;
  assign v_11256 = ~v_11243;
  assign v_11257 = mux_11257(v_11258);
  assign v_11258 = ~v_11253;
  pebbles_core
    pebbles_core_11259
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11260),
       .in0_consume_en(vin0_consume_en_11259),
       .out_canPeek(vout_canPeek_11259),
       .out_peek(vout_peek_11259));
  assign v_11260 = v_11261 | v_11262;
  assign v_11261 = mux_11261(v_11247);
  assign v_11262 = mux_11262(v_11263);
  assign v_11263 = ~v_11247;
  assign v_11264 = v_11265 & 1'h1;
  assign v_11265 = v_11266 & v_11267;
  assign v_11266 = ~act_11246;
  assign v_11267 = v_11268 | v_11272;
  assign v_11268 = v_11269 | v_11270;
  assign v_11269 = mux_11269(v_11203);
  assign v_11270 = mux_11270(v_11271);
  assign v_11271 = ~v_11203;
  assign v_11272 = ~v_11243;
  assign v_11273 = v_11274 | v_11275;
  assign v_11274 = mux_11274(v_11245);
  assign v_11275 = mux_11275(v_11264);
  assign v_11276 = v_11277 & 1'h1;
  assign v_11277 = v_11278 & v_11279;
  assign v_11278 = ~act_11202;
  assign v_11279 = v_11280 | v_11284;
  assign v_11280 = v_11281 | v_11282;
  assign v_11281 = mux_11281(v_11103);
  assign v_11282 = mux_11282(v_11283);
  assign v_11283 = ~v_11103;
  assign v_11284 = ~v_11199;
  assign v_11285 = v_11286 | v_11287;
  assign v_11286 = mux_11286(v_11201);
  assign v_11287 = mux_11287(v_11276);
  assign v_11288 = v_11289 & 1'h1;
  assign v_11289 = v_11290 & v_11291;
  assign v_11290 = ~act_11102;
  assign v_11291 = v_11292 | v_11300;
  assign v_11292 = v_11293 | v_11298;
  assign v_11293 = mux_11293(v_11294);
  assign v_11294 = v_11099 & v_11295;
  assign v_11295 = v_11296 & 1'h1;
  assign v_11296 = v_11297 | 1'h0;
  assign v_11297 = ~v_11092;
  assign v_11298 = mux_11298(v_11299);
  assign v_11299 = ~v_11294;
  assign v_11300 = ~v_11099;
  assign v_11301 = v_11302 | v_11303;
  assign v_11302 = mux_11302(v_11101);
  assign v_11303 = mux_11303(v_11288);
  assign v_11305 = v_11306 | v_11493;
  assign v_11306 = act_11307 & 1'h1;
  assign act_11307 = v_11308 | v_11394;
  assign v_11308 = v_11309 & v_11395;
  assign v_11309 = v_11310 & v_11404;
  assign v_11310 = ~v_11311;
  assign v_11312 = v_11313 | v_11388;
  assign v_11313 = act_11314 & 1'h1;
  assign act_11314 = v_11315 | v_11345;
  assign v_11315 = v_11316 & v_11346;
  assign v_11316 = v_11317 & v_11355;
  assign v_11317 = ~v_11318;
  assign v_11319 = v_11320 | v_11339;
  assign v_11320 = act_11321 & 1'h1;
  assign act_11321 = v_11322 | v_11328;
  assign v_11322 = v_11323 & v_11329;
  assign v_11323 = v_11324 & vout_canPeek_11334;
  assign v_11324 = ~vout_canPeek_11325;
  pebbles_core
    pebbles_core_11325
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11326),
       .in0_consume_en(vin0_consume_en_11325),
       .out_canPeek(vout_canPeek_11325),
       .out_peek(vout_peek_11325));
  assign v_11326 = v_11327 | v_11332;
  assign v_11327 = mux_11327(v_11328);
  assign v_11328 = vout_canPeek_11325 & v_11329;
  assign v_11329 = v_11330 & 1'h1;
  assign v_11330 = v_11331 | 1'h0;
  assign v_11331 = ~v_11318;
  assign v_11332 = mux_11332(v_11333);
  assign v_11333 = ~v_11328;
  pebbles_core
    pebbles_core_11334
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11335),
       .in0_consume_en(vin0_consume_en_11334),
       .out_canPeek(vout_canPeek_11334),
       .out_peek(vout_peek_11334));
  assign v_11335 = v_11336 | v_11337;
  assign v_11336 = mux_11336(v_11322);
  assign v_11337 = mux_11337(v_11338);
  assign v_11338 = ~v_11322;
  assign v_11339 = v_11340 & 1'h1;
  assign v_11340 = v_11341 & v_11342;
  assign v_11341 = ~act_11321;
  assign v_11342 = v_11343 | v_11351;
  assign v_11343 = v_11344 | v_11349;
  assign v_11344 = mux_11344(v_11345);
  assign v_11345 = v_11318 & v_11346;
  assign v_11346 = v_11347 & 1'h1;
  assign v_11347 = v_11348 | 1'h0;
  assign v_11348 = ~v_11311;
  assign v_11349 = mux_11349(v_11350);
  assign v_11350 = ~v_11345;
  assign v_11351 = ~v_11318;
  assign v_11352 = v_11353 | v_11354;
  assign v_11353 = mux_11353(v_11320);
  assign v_11354 = mux_11354(v_11339);
  assign v_11356 = v_11357 | v_11376;
  assign v_11357 = act_11358 & 1'h1;
  assign act_11358 = v_11359 | v_11365;
  assign v_11359 = v_11360 & v_11366;
  assign v_11360 = v_11361 & vout_canPeek_11371;
  assign v_11361 = ~vout_canPeek_11362;
  pebbles_core
    pebbles_core_11362
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11363),
       .in0_consume_en(vin0_consume_en_11362),
       .out_canPeek(vout_canPeek_11362),
       .out_peek(vout_peek_11362));
  assign v_11363 = v_11364 | v_11369;
  assign v_11364 = mux_11364(v_11365);
  assign v_11365 = vout_canPeek_11362 & v_11366;
  assign v_11366 = v_11367 & 1'h1;
  assign v_11367 = v_11368 | 1'h0;
  assign v_11368 = ~v_11355;
  assign v_11369 = mux_11369(v_11370);
  assign v_11370 = ~v_11365;
  pebbles_core
    pebbles_core_11371
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11372),
       .in0_consume_en(vin0_consume_en_11371),
       .out_canPeek(vout_canPeek_11371),
       .out_peek(vout_peek_11371));
  assign v_11372 = v_11373 | v_11374;
  assign v_11373 = mux_11373(v_11359);
  assign v_11374 = mux_11374(v_11375);
  assign v_11375 = ~v_11359;
  assign v_11376 = v_11377 & 1'h1;
  assign v_11377 = v_11378 & v_11379;
  assign v_11378 = ~act_11358;
  assign v_11379 = v_11380 | v_11384;
  assign v_11380 = v_11381 | v_11382;
  assign v_11381 = mux_11381(v_11315);
  assign v_11382 = mux_11382(v_11383);
  assign v_11383 = ~v_11315;
  assign v_11384 = ~v_11355;
  assign v_11385 = v_11386 | v_11387;
  assign v_11386 = mux_11386(v_11357);
  assign v_11387 = mux_11387(v_11376);
  assign v_11388 = v_11389 & 1'h1;
  assign v_11389 = v_11390 & v_11391;
  assign v_11390 = ~act_11314;
  assign v_11391 = v_11392 | v_11400;
  assign v_11392 = v_11393 | v_11398;
  assign v_11393 = mux_11393(v_11394);
  assign v_11394 = v_11311 & v_11395;
  assign v_11395 = v_11396 & 1'h1;
  assign v_11396 = v_11397 | 1'h0;
  assign v_11397 = ~v_11304;
  assign v_11398 = mux_11398(v_11399);
  assign v_11399 = ~v_11394;
  assign v_11400 = ~v_11311;
  assign v_11401 = v_11402 | v_11403;
  assign v_11402 = mux_11402(v_11313);
  assign v_11403 = mux_11403(v_11388);
  assign v_11405 = v_11406 | v_11481;
  assign v_11406 = act_11407 & 1'h1;
  assign act_11407 = v_11408 | v_11438;
  assign v_11408 = v_11409 & v_11439;
  assign v_11409 = v_11410 & v_11448;
  assign v_11410 = ~v_11411;
  assign v_11412 = v_11413 | v_11432;
  assign v_11413 = act_11414 & 1'h1;
  assign act_11414 = v_11415 | v_11421;
  assign v_11415 = v_11416 & v_11422;
  assign v_11416 = v_11417 & vout_canPeek_11427;
  assign v_11417 = ~vout_canPeek_11418;
  pebbles_core
    pebbles_core_11418
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11419),
       .in0_consume_en(vin0_consume_en_11418),
       .out_canPeek(vout_canPeek_11418),
       .out_peek(vout_peek_11418));
  assign v_11419 = v_11420 | v_11425;
  assign v_11420 = mux_11420(v_11421);
  assign v_11421 = vout_canPeek_11418 & v_11422;
  assign v_11422 = v_11423 & 1'h1;
  assign v_11423 = v_11424 | 1'h0;
  assign v_11424 = ~v_11411;
  assign v_11425 = mux_11425(v_11426);
  assign v_11426 = ~v_11421;
  pebbles_core
    pebbles_core_11427
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11428),
       .in0_consume_en(vin0_consume_en_11427),
       .out_canPeek(vout_canPeek_11427),
       .out_peek(vout_peek_11427));
  assign v_11428 = v_11429 | v_11430;
  assign v_11429 = mux_11429(v_11415);
  assign v_11430 = mux_11430(v_11431);
  assign v_11431 = ~v_11415;
  assign v_11432 = v_11433 & 1'h1;
  assign v_11433 = v_11434 & v_11435;
  assign v_11434 = ~act_11414;
  assign v_11435 = v_11436 | v_11444;
  assign v_11436 = v_11437 | v_11442;
  assign v_11437 = mux_11437(v_11438);
  assign v_11438 = v_11411 & v_11439;
  assign v_11439 = v_11440 & 1'h1;
  assign v_11440 = v_11441 | 1'h0;
  assign v_11441 = ~v_11404;
  assign v_11442 = mux_11442(v_11443);
  assign v_11443 = ~v_11438;
  assign v_11444 = ~v_11411;
  assign v_11445 = v_11446 | v_11447;
  assign v_11446 = mux_11446(v_11413);
  assign v_11447 = mux_11447(v_11432);
  assign v_11449 = v_11450 | v_11469;
  assign v_11450 = act_11451 & 1'h1;
  assign act_11451 = v_11452 | v_11458;
  assign v_11452 = v_11453 & v_11459;
  assign v_11453 = v_11454 & vout_canPeek_11464;
  assign v_11454 = ~vout_canPeek_11455;
  pebbles_core
    pebbles_core_11455
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11456),
       .in0_consume_en(vin0_consume_en_11455),
       .out_canPeek(vout_canPeek_11455),
       .out_peek(vout_peek_11455));
  assign v_11456 = v_11457 | v_11462;
  assign v_11457 = mux_11457(v_11458);
  assign v_11458 = vout_canPeek_11455 & v_11459;
  assign v_11459 = v_11460 & 1'h1;
  assign v_11460 = v_11461 | 1'h0;
  assign v_11461 = ~v_11448;
  assign v_11462 = mux_11462(v_11463);
  assign v_11463 = ~v_11458;
  pebbles_core
    pebbles_core_11464
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11465),
       .in0_consume_en(vin0_consume_en_11464),
       .out_canPeek(vout_canPeek_11464),
       .out_peek(vout_peek_11464));
  assign v_11465 = v_11466 | v_11467;
  assign v_11466 = mux_11466(v_11452);
  assign v_11467 = mux_11467(v_11468);
  assign v_11468 = ~v_11452;
  assign v_11469 = v_11470 & 1'h1;
  assign v_11470 = v_11471 & v_11472;
  assign v_11471 = ~act_11451;
  assign v_11472 = v_11473 | v_11477;
  assign v_11473 = v_11474 | v_11475;
  assign v_11474 = mux_11474(v_11408);
  assign v_11475 = mux_11475(v_11476);
  assign v_11476 = ~v_11408;
  assign v_11477 = ~v_11448;
  assign v_11478 = v_11479 | v_11480;
  assign v_11479 = mux_11479(v_11450);
  assign v_11480 = mux_11480(v_11469);
  assign v_11481 = v_11482 & 1'h1;
  assign v_11482 = v_11483 & v_11484;
  assign v_11483 = ~act_11407;
  assign v_11484 = v_11485 | v_11489;
  assign v_11485 = v_11486 | v_11487;
  assign v_11486 = mux_11486(v_11308);
  assign v_11487 = mux_11487(v_11488);
  assign v_11488 = ~v_11308;
  assign v_11489 = ~v_11404;
  assign v_11490 = v_11491 | v_11492;
  assign v_11491 = mux_11491(v_11406);
  assign v_11492 = mux_11492(v_11481);
  assign v_11493 = v_11494 & 1'h1;
  assign v_11494 = v_11495 & v_11496;
  assign v_11495 = ~act_11307;
  assign v_11496 = v_11497 | v_11501;
  assign v_11497 = v_11498 | v_11499;
  assign v_11498 = mux_11498(v_11096);
  assign v_11499 = mux_11499(v_11500);
  assign v_11500 = ~v_11096;
  assign v_11501 = ~v_11304;
  assign v_11502 = v_11503 | v_11504;
  assign v_11503 = mux_11503(v_11306);
  assign v_11504 = mux_11504(v_11493);
  assign v_11505 = v_11506 & 1'h1;
  assign v_11506 = v_11507 & v_11508;
  assign v_11507 = ~act_11095;
  assign v_11508 = v_11509 | v_11513;
  assign v_11509 = v_11510 | v_11511;
  assign v_11510 = mux_11510(v_10660);
  assign v_11511 = mux_11511(v_11512);
  assign v_11512 = ~v_10660;
  assign v_11513 = ~v_11092;
  assign v_11514 = v_11515 | v_11516;
  assign v_11515 = mux_11515(v_11094);
  assign v_11516 = mux_11516(v_11505);
  assign v_11517 = v_11518 & 1'h1;
  assign v_11518 = v_11519 & v_11520;
  assign v_11519 = ~act_10659;
  assign v_11520 = v_11521 | v_11525;
  assign v_11521 = v_11522 | v_11523;
  assign v_11522 = mux_11522(v_9776);
  assign v_11523 = mux_11523(v_11524);
  assign v_11524 = ~v_9776;
  assign v_11525 = ~v_10656;
  assign v_11526 = v_11527 | v_11528;
  assign v_11527 = mux_11527(v_10658);
  assign v_11528 = mux_11528(v_11517);
  assign v_11529 = v_11530 & 1'h1;
  assign v_11530 = v_11531 & v_11532;
  assign v_11531 = ~act_9775;
  assign v_11532 = v_11533 | v_11537;
  assign v_11533 = v_11534 | v_11535;
  assign v_11534 = mux_11534(v_7996);
  assign v_11535 = mux_11535(v_11536);
  assign v_11536 = ~v_7996;
  assign v_11537 = ~v_9772;
  assign v_11538 = v_11539 | v_11540;
  assign v_11539 = mux_11539(v_9774);
  assign v_11540 = mux_11540(v_11529);
  assign v_11541 = v_11542 & 1'h1;
  assign v_11542 = v_11543 & v_11544;
  assign v_11543 = ~act_7995;
  assign v_11544 = v_11545 | v_11553;
  assign v_11545 = v_11546 | v_11551;
  assign v_11546 = mux_11546(v_11547);
  assign v_11547 = v_7992 & v_11548;
  assign v_11548 = v_11549 & 1'h1;
  assign v_11549 = v_11550 | 1'h0;
  assign v_11550 = ~v_7985;
  assign v_11551 = mux_11551(v_11552);
  assign v_11552 = ~v_11547;
  assign v_11553 = ~v_7992;
  assign v_11554 = v_11555 | v_11556;
  assign v_11555 = mux_11555(v_7994);
  assign v_11556 = mux_11556(v_11541);
  assign v_11558 = v_11559 | v_15106;
  assign v_11559 = act_11560 & 1'h1;
  assign act_11560 = v_11561 | v_13327;
  assign v_11561 = v_11562 & v_13328;
  assign v_11562 = v_11563 & v_13337;
  assign v_11563 = ~v_11564;
  assign v_11565 = v_11566 | v_13321;
  assign v_11566 = act_11567 & 1'h1;
  assign act_11567 = v_11568 | v_12438;
  assign v_11568 = v_11569 & v_12439;
  assign v_11569 = v_11570 & v_12448;
  assign v_11570 = ~v_11571;
  assign v_11572 = v_11573 | v_12432;
  assign v_11573 = act_11574 & 1'h1;
  assign act_11574 = v_11575 | v_11997;
  assign v_11575 = v_11576 & v_11998;
  assign v_11576 = v_11577 & v_12007;
  assign v_11577 = ~v_11578;
  assign v_11579 = v_11580 | v_11991;
  assign v_11580 = act_11581 & 1'h1;
  assign act_11581 = v_11582 | v_11780;
  assign v_11582 = v_11583 & v_11781;
  assign v_11583 = v_11584 & v_11790;
  assign v_11584 = ~v_11585;
  assign v_11586 = v_11587 | v_11774;
  assign v_11587 = act_11588 & 1'h1;
  assign act_11588 = v_11589 | v_11675;
  assign v_11589 = v_11590 & v_11676;
  assign v_11590 = v_11591 & v_11685;
  assign v_11591 = ~v_11592;
  assign v_11593 = v_11594 | v_11669;
  assign v_11594 = act_11595 & 1'h1;
  assign act_11595 = v_11596 | v_11626;
  assign v_11596 = v_11597 & v_11627;
  assign v_11597 = v_11598 & v_11636;
  assign v_11598 = ~v_11599;
  assign v_11600 = v_11601 | v_11620;
  assign v_11601 = act_11602 & 1'h1;
  assign act_11602 = v_11603 | v_11609;
  assign v_11603 = v_11604 & v_11610;
  assign v_11604 = v_11605 & vout_canPeek_11615;
  assign v_11605 = ~vout_canPeek_11606;
  pebbles_core
    pebbles_core_11606
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11607),
       .in0_consume_en(vin0_consume_en_11606),
       .out_canPeek(vout_canPeek_11606),
       .out_peek(vout_peek_11606));
  assign v_11607 = v_11608 | v_11613;
  assign v_11608 = mux_11608(v_11609);
  assign v_11609 = vout_canPeek_11606 & v_11610;
  assign v_11610 = v_11611 & 1'h1;
  assign v_11611 = v_11612 | 1'h0;
  assign v_11612 = ~v_11599;
  assign v_11613 = mux_11613(v_11614);
  assign v_11614 = ~v_11609;
  pebbles_core
    pebbles_core_11615
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11616),
       .in0_consume_en(vin0_consume_en_11615),
       .out_canPeek(vout_canPeek_11615),
       .out_peek(vout_peek_11615));
  assign v_11616 = v_11617 | v_11618;
  assign v_11617 = mux_11617(v_11603);
  assign v_11618 = mux_11618(v_11619);
  assign v_11619 = ~v_11603;
  assign v_11620 = v_11621 & 1'h1;
  assign v_11621 = v_11622 & v_11623;
  assign v_11622 = ~act_11602;
  assign v_11623 = v_11624 | v_11632;
  assign v_11624 = v_11625 | v_11630;
  assign v_11625 = mux_11625(v_11626);
  assign v_11626 = v_11599 & v_11627;
  assign v_11627 = v_11628 & 1'h1;
  assign v_11628 = v_11629 | 1'h0;
  assign v_11629 = ~v_11592;
  assign v_11630 = mux_11630(v_11631);
  assign v_11631 = ~v_11626;
  assign v_11632 = ~v_11599;
  assign v_11633 = v_11634 | v_11635;
  assign v_11634 = mux_11634(v_11601);
  assign v_11635 = mux_11635(v_11620);
  assign v_11637 = v_11638 | v_11657;
  assign v_11638 = act_11639 & 1'h1;
  assign act_11639 = v_11640 | v_11646;
  assign v_11640 = v_11641 & v_11647;
  assign v_11641 = v_11642 & vout_canPeek_11652;
  assign v_11642 = ~vout_canPeek_11643;
  pebbles_core
    pebbles_core_11643
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11644),
       .in0_consume_en(vin0_consume_en_11643),
       .out_canPeek(vout_canPeek_11643),
       .out_peek(vout_peek_11643));
  assign v_11644 = v_11645 | v_11650;
  assign v_11645 = mux_11645(v_11646);
  assign v_11646 = vout_canPeek_11643 & v_11647;
  assign v_11647 = v_11648 & 1'h1;
  assign v_11648 = v_11649 | 1'h0;
  assign v_11649 = ~v_11636;
  assign v_11650 = mux_11650(v_11651);
  assign v_11651 = ~v_11646;
  pebbles_core
    pebbles_core_11652
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11653),
       .in0_consume_en(vin0_consume_en_11652),
       .out_canPeek(vout_canPeek_11652),
       .out_peek(vout_peek_11652));
  assign v_11653 = v_11654 | v_11655;
  assign v_11654 = mux_11654(v_11640);
  assign v_11655 = mux_11655(v_11656);
  assign v_11656 = ~v_11640;
  assign v_11657 = v_11658 & 1'h1;
  assign v_11658 = v_11659 & v_11660;
  assign v_11659 = ~act_11639;
  assign v_11660 = v_11661 | v_11665;
  assign v_11661 = v_11662 | v_11663;
  assign v_11662 = mux_11662(v_11596);
  assign v_11663 = mux_11663(v_11664);
  assign v_11664 = ~v_11596;
  assign v_11665 = ~v_11636;
  assign v_11666 = v_11667 | v_11668;
  assign v_11667 = mux_11667(v_11638);
  assign v_11668 = mux_11668(v_11657);
  assign v_11669 = v_11670 & 1'h1;
  assign v_11670 = v_11671 & v_11672;
  assign v_11671 = ~act_11595;
  assign v_11672 = v_11673 | v_11681;
  assign v_11673 = v_11674 | v_11679;
  assign v_11674 = mux_11674(v_11675);
  assign v_11675 = v_11592 & v_11676;
  assign v_11676 = v_11677 & 1'h1;
  assign v_11677 = v_11678 | 1'h0;
  assign v_11678 = ~v_11585;
  assign v_11679 = mux_11679(v_11680);
  assign v_11680 = ~v_11675;
  assign v_11681 = ~v_11592;
  assign v_11682 = v_11683 | v_11684;
  assign v_11683 = mux_11683(v_11594);
  assign v_11684 = mux_11684(v_11669);
  assign v_11686 = v_11687 | v_11762;
  assign v_11687 = act_11688 & 1'h1;
  assign act_11688 = v_11689 | v_11719;
  assign v_11689 = v_11690 & v_11720;
  assign v_11690 = v_11691 & v_11729;
  assign v_11691 = ~v_11692;
  assign v_11693 = v_11694 | v_11713;
  assign v_11694 = act_11695 & 1'h1;
  assign act_11695 = v_11696 | v_11702;
  assign v_11696 = v_11697 & v_11703;
  assign v_11697 = v_11698 & vout_canPeek_11708;
  assign v_11698 = ~vout_canPeek_11699;
  pebbles_core
    pebbles_core_11699
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11700),
       .in0_consume_en(vin0_consume_en_11699),
       .out_canPeek(vout_canPeek_11699),
       .out_peek(vout_peek_11699));
  assign v_11700 = v_11701 | v_11706;
  assign v_11701 = mux_11701(v_11702);
  assign v_11702 = vout_canPeek_11699 & v_11703;
  assign v_11703 = v_11704 & 1'h1;
  assign v_11704 = v_11705 | 1'h0;
  assign v_11705 = ~v_11692;
  assign v_11706 = mux_11706(v_11707);
  assign v_11707 = ~v_11702;
  pebbles_core
    pebbles_core_11708
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11709),
       .in0_consume_en(vin0_consume_en_11708),
       .out_canPeek(vout_canPeek_11708),
       .out_peek(vout_peek_11708));
  assign v_11709 = v_11710 | v_11711;
  assign v_11710 = mux_11710(v_11696);
  assign v_11711 = mux_11711(v_11712);
  assign v_11712 = ~v_11696;
  assign v_11713 = v_11714 & 1'h1;
  assign v_11714 = v_11715 & v_11716;
  assign v_11715 = ~act_11695;
  assign v_11716 = v_11717 | v_11725;
  assign v_11717 = v_11718 | v_11723;
  assign v_11718 = mux_11718(v_11719);
  assign v_11719 = v_11692 & v_11720;
  assign v_11720 = v_11721 & 1'h1;
  assign v_11721 = v_11722 | 1'h0;
  assign v_11722 = ~v_11685;
  assign v_11723 = mux_11723(v_11724);
  assign v_11724 = ~v_11719;
  assign v_11725 = ~v_11692;
  assign v_11726 = v_11727 | v_11728;
  assign v_11727 = mux_11727(v_11694);
  assign v_11728 = mux_11728(v_11713);
  assign v_11730 = v_11731 | v_11750;
  assign v_11731 = act_11732 & 1'h1;
  assign act_11732 = v_11733 | v_11739;
  assign v_11733 = v_11734 & v_11740;
  assign v_11734 = v_11735 & vout_canPeek_11745;
  assign v_11735 = ~vout_canPeek_11736;
  pebbles_core
    pebbles_core_11736
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11737),
       .in0_consume_en(vin0_consume_en_11736),
       .out_canPeek(vout_canPeek_11736),
       .out_peek(vout_peek_11736));
  assign v_11737 = v_11738 | v_11743;
  assign v_11738 = mux_11738(v_11739);
  assign v_11739 = vout_canPeek_11736 & v_11740;
  assign v_11740 = v_11741 & 1'h1;
  assign v_11741 = v_11742 | 1'h0;
  assign v_11742 = ~v_11729;
  assign v_11743 = mux_11743(v_11744);
  assign v_11744 = ~v_11739;
  pebbles_core
    pebbles_core_11745
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11746),
       .in0_consume_en(vin0_consume_en_11745),
       .out_canPeek(vout_canPeek_11745),
       .out_peek(vout_peek_11745));
  assign v_11746 = v_11747 | v_11748;
  assign v_11747 = mux_11747(v_11733);
  assign v_11748 = mux_11748(v_11749);
  assign v_11749 = ~v_11733;
  assign v_11750 = v_11751 & 1'h1;
  assign v_11751 = v_11752 & v_11753;
  assign v_11752 = ~act_11732;
  assign v_11753 = v_11754 | v_11758;
  assign v_11754 = v_11755 | v_11756;
  assign v_11755 = mux_11755(v_11689);
  assign v_11756 = mux_11756(v_11757);
  assign v_11757 = ~v_11689;
  assign v_11758 = ~v_11729;
  assign v_11759 = v_11760 | v_11761;
  assign v_11760 = mux_11760(v_11731);
  assign v_11761 = mux_11761(v_11750);
  assign v_11762 = v_11763 & 1'h1;
  assign v_11763 = v_11764 & v_11765;
  assign v_11764 = ~act_11688;
  assign v_11765 = v_11766 | v_11770;
  assign v_11766 = v_11767 | v_11768;
  assign v_11767 = mux_11767(v_11589);
  assign v_11768 = mux_11768(v_11769);
  assign v_11769 = ~v_11589;
  assign v_11770 = ~v_11685;
  assign v_11771 = v_11772 | v_11773;
  assign v_11772 = mux_11772(v_11687);
  assign v_11773 = mux_11773(v_11762);
  assign v_11774 = v_11775 & 1'h1;
  assign v_11775 = v_11776 & v_11777;
  assign v_11776 = ~act_11588;
  assign v_11777 = v_11778 | v_11786;
  assign v_11778 = v_11779 | v_11784;
  assign v_11779 = mux_11779(v_11780);
  assign v_11780 = v_11585 & v_11781;
  assign v_11781 = v_11782 & 1'h1;
  assign v_11782 = v_11783 | 1'h0;
  assign v_11783 = ~v_11578;
  assign v_11784 = mux_11784(v_11785);
  assign v_11785 = ~v_11780;
  assign v_11786 = ~v_11585;
  assign v_11787 = v_11788 | v_11789;
  assign v_11788 = mux_11788(v_11587);
  assign v_11789 = mux_11789(v_11774);
  assign v_11791 = v_11792 | v_11979;
  assign v_11792 = act_11793 & 1'h1;
  assign act_11793 = v_11794 | v_11880;
  assign v_11794 = v_11795 & v_11881;
  assign v_11795 = v_11796 & v_11890;
  assign v_11796 = ~v_11797;
  assign v_11798 = v_11799 | v_11874;
  assign v_11799 = act_11800 & 1'h1;
  assign act_11800 = v_11801 | v_11831;
  assign v_11801 = v_11802 & v_11832;
  assign v_11802 = v_11803 & v_11841;
  assign v_11803 = ~v_11804;
  assign v_11805 = v_11806 | v_11825;
  assign v_11806 = act_11807 & 1'h1;
  assign act_11807 = v_11808 | v_11814;
  assign v_11808 = v_11809 & v_11815;
  assign v_11809 = v_11810 & vout_canPeek_11820;
  assign v_11810 = ~vout_canPeek_11811;
  pebbles_core
    pebbles_core_11811
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11812),
       .in0_consume_en(vin0_consume_en_11811),
       .out_canPeek(vout_canPeek_11811),
       .out_peek(vout_peek_11811));
  assign v_11812 = v_11813 | v_11818;
  assign v_11813 = mux_11813(v_11814);
  assign v_11814 = vout_canPeek_11811 & v_11815;
  assign v_11815 = v_11816 & 1'h1;
  assign v_11816 = v_11817 | 1'h0;
  assign v_11817 = ~v_11804;
  assign v_11818 = mux_11818(v_11819);
  assign v_11819 = ~v_11814;
  pebbles_core
    pebbles_core_11820
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11821),
       .in0_consume_en(vin0_consume_en_11820),
       .out_canPeek(vout_canPeek_11820),
       .out_peek(vout_peek_11820));
  assign v_11821 = v_11822 | v_11823;
  assign v_11822 = mux_11822(v_11808);
  assign v_11823 = mux_11823(v_11824);
  assign v_11824 = ~v_11808;
  assign v_11825 = v_11826 & 1'h1;
  assign v_11826 = v_11827 & v_11828;
  assign v_11827 = ~act_11807;
  assign v_11828 = v_11829 | v_11837;
  assign v_11829 = v_11830 | v_11835;
  assign v_11830 = mux_11830(v_11831);
  assign v_11831 = v_11804 & v_11832;
  assign v_11832 = v_11833 & 1'h1;
  assign v_11833 = v_11834 | 1'h0;
  assign v_11834 = ~v_11797;
  assign v_11835 = mux_11835(v_11836);
  assign v_11836 = ~v_11831;
  assign v_11837 = ~v_11804;
  assign v_11838 = v_11839 | v_11840;
  assign v_11839 = mux_11839(v_11806);
  assign v_11840 = mux_11840(v_11825);
  assign v_11842 = v_11843 | v_11862;
  assign v_11843 = act_11844 & 1'h1;
  assign act_11844 = v_11845 | v_11851;
  assign v_11845 = v_11846 & v_11852;
  assign v_11846 = v_11847 & vout_canPeek_11857;
  assign v_11847 = ~vout_canPeek_11848;
  pebbles_core
    pebbles_core_11848
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11849),
       .in0_consume_en(vin0_consume_en_11848),
       .out_canPeek(vout_canPeek_11848),
       .out_peek(vout_peek_11848));
  assign v_11849 = v_11850 | v_11855;
  assign v_11850 = mux_11850(v_11851);
  assign v_11851 = vout_canPeek_11848 & v_11852;
  assign v_11852 = v_11853 & 1'h1;
  assign v_11853 = v_11854 | 1'h0;
  assign v_11854 = ~v_11841;
  assign v_11855 = mux_11855(v_11856);
  assign v_11856 = ~v_11851;
  pebbles_core
    pebbles_core_11857
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11858),
       .in0_consume_en(vin0_consume_en_11857),
       .out_canPeek(vout_canPeek_11857),
       .out_peek(vout_peek_11857));
  assign v_11858 = v_11859 | v_11860;
  assign v_11859 = mux_11859(v_11845);
  assign v_11860 = mux_11860(v_11861);
  assign v_11861 = ~v_11845;
  assign v_11862 = v_11863 & 1'h1;
  assign v_11863 = v_11864 & v_11865;
  assign v_11864 = ~act_11844;
  assign v_11865 = v_11866 | v_11870;
  assign v_11866 = v_11867 | v_11868;
  assign v_11867 = mux_11867(v_11801);
  assign v_11868 = mux_11868(v_11869);
  assign v_11869 = ~v_11801;
  assign v_11870 = ~v_11841;
  assign v_11871 = v_11872 | v_11873;
  assign v_11872 = mux_11872(v_11843);
  assign v_11873 = mux_11873(v_11862);
  assign v_11874 = v_11875 & 1'h1;
  assign v_11875 = v_11876 & v_11877;
  assign v_11876 = ~act_11800;
  assign v_11877 = v_11878 | v_11886;
  assign v_11878 = v_11879 | v_11884;
  assign v_11879 = mux_11879(v_11880);
  assign v_11880 = v_11797 & v_11881;
  assign v_11881 = v_11882 & 1'h1;
  assign v_11882 = v_11883 | 1'h0;
  assign v_11883 = ~v_11790;
  assign v_11884 = mux_11884(v_11885);
  assign v_11885 = ~v_11880;
  assign v_11886 = ~v_11797;
  assign v_11887 = v_11888 | v_11889;
  assign v_11888 = mux_11888(v_11799);
  assign v_11889 = mux_11889(v_11874);
  assign v_11891 = v_11892 | v_11967;
  assign v_11892 = act_11893 & 1'h1;
  assign act_11893 = v_11894 | v_11924;
  assign v_11894 = v_11895 & v_11925;
  assign v_11895 = v_11896 & v_11934;
  assign v_11896 = ~v_11897;
  assign v_11898 = v_11899 | v_11918;
  assign v_11899 = act_11900 & 1'h1;
  assign act_11900 = v_11901 | v_11907;
  assign v_11901 = v_11902 & v_11908;
  assign v_11902 = v_11903 & vout_canPeek_11913;
  assign v_11903 = ~vout_canPeek_11904;
  pebbles_core
    pebbles_core_11904
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11905),
       .in0_consume_en(vin0_consume_en_11904),
       .out_canPeek(vout_canPeek_11904),
       .out_peek(vout_peek_11904));
  assign v_11905 = v_11906 | v_11911;
  assign v_11906 = mux_11906(v_11907);
  assign v_11907 = vout_canPeek_11904 & v_11908;
  assign v_11908 = v_11909 & 1'h1;
  assign v_11909 = v_11910 | 1'h0;
  assign v_11910 = ~v_11897;
  assign v_11911 = mux_11911(v_11912);
  assign v_11912 = ~v_11907;
  pebbles_core
    pebbles_core_11913
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11914),
       .in0_consume_en(vin0_consume_en_11913),
       .out_canPeek(vout_canPeek_11913),
       .out_peek(vout_peek_11913));
  assign v_11914 = v_11915 | v_11916;
  assign v_11915 = mux_11915(v_11901);
  assign v_11916 = mux_11916(v_11917);
  assign v_11917 = ~v_11901;
  assign v_11918 = v_11919 & 1'h1;
  assign v_11919 = v_11920 & v_11921;
  assign v_11920 = ~act_11900;
  assign v_11921 = v_11922 | v_11930;
  assign v_11922 = v_11923 | v_11928;
  assign v_11923 = mux_11923(v_11924);
  assign v_11924 = v_11897 & v_11925;
  assign v_11925 = v_11926 & 1'h1;
  assign v_11926 = v_11927 | 1'h0;
  assign v_11927 = ~v_11890;
  assign v_11928 = mux_11928(v_11929);
  assign v_11929 = ~v_11924;
  assign v_11930 = ~v_11897;
  assign v_11931 = v_11932 | v_11933;
  assign v_11932 = mux_11932(v_11899);
  assign v_11933 = mux_11933(v_11918);
  assign v_11935 = v_11936 | v_11955;
  assign v_11936 = act_11937 & 1'h1;
  assign act_11937 = v_11938 | v_11944;
  assign v_11938 = v_11939 & v_11945;
  assign v_11939 = v_11940 & vout_canPeek_11950;
  assign v_11940 = ~vout_canPeek_11941;
  pebbles_core
    pebbles_core_11941
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11942),
       .in0_consume_en(vin0_consume_en_11941),
       .out_canPeek(vout_canPeek_11941),
       .out_peek(vout_peek_11941));
  assign v_11942 = v_11943 | v_11948;
  assign v_11943 = mux_11943(v_11944);
  assign v_11944 = vout_canPeek_11941 & v_11945;
  assign v_11945 = v_11946 & 1'h1;
  assign v_11946 = v_11947 | 1'h0;
  assign v_11947 = ~v_11934;
  assign v_11948 = mux_11948(v_11949);
  assign v_11949 = ~v_11944;
  pebbles_core
    pebbles_core_11950
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_11951),
       .in0_consume_en(vin0_consume_en_11950),
       .out_canPeek(vout_canPeek_11950),
       .out_peek(vout_peek_11950));
  assign v_11951 = v_11952 | v_11953;
  assign v_11952 = mux_11952(v_11938);
  assign v_11953 = mux_11953(v_11954);
  assign v_11954 = ~v_11938;
  assign v_11955 = v_11956 & 1'h1;
  assign v_11956 = v_11957 & v_11958;
  assign v_11957 = ~act_11937;
  assign v_11958 = v_11959 | v_11963;
  assign v_11959 = v_11960 | v_11961;
  assign v_11960 = mux_11960(v_11894);
  assign v_11961 = mux_11961(v_11962);
  assign v_11962 = ~v_11894;
  assign v_11963 = ~v_11934;
  assign v_11964 = v_11965 | v_11966;
  assign v_11965 = mux_11965(v_11936);
  assign v_11966 = mux_11966(v_11955);
  assign v_11967 = v_11968 & 1'h1;
  assign v_11968 = v_11969 & v_11970;
  assign v_11969 = ~act_11893;
  assign v_11970 = v_11971 | v_11975;
  assign v_11971 = v_11972 | v_11973;
  assign v_11972 = mux_11972(v_11794);
  assign v_11973 = mux_11973(v_11974);
  assign v_11974 = ~v_11794;
  assign v_11975 = ~v_11890;
  assign v_11976 = v_11977 | v_11978;
  assign v_11977 = mux_11977(v_11892);
  assign v_11978 = mux_11978(v_11967);
  assign v_11979 = v_11980 & 1'h1;
  assign v_11980 = v_11981 & v_11982;
  assign v_11981 = ~act_11793;
  assign v_11982 = v_11983 | v_11987;
  assign v_11983 = v_11984 | v_11985;
  assign v_11984 = mux_11984(v_11582);
  assign v_11985 = mux_11985(v_11986);
  assign v_11986 = ~v_11582;
  assign v_11987 = ~v_11790;
  assign v_11988 = v_11989 | v_11990;
  assign v_11989 = mux_11989(v_11792);
  assign v_11990 = mux_11990(v_11979);
  assign v_11991 = v_11992 & 1'h1;
  assign v_11992 = v_11993 & v_11994;
  assign v_11993 = ~act_11581;
  assign v_11994 = v_11995 | v_12003;
  assign v_11995 = v_11996 | v_12001;
  assign v_11996 = mux_11996(v_11997);
  assign v_11997 = v_11578 & v_11998;
  assign v_11998 = v_11999 & 1'h1;
  assign v_11999 = v_12000 | 1'h0;
  assign v_12000 = ~v_11571;
  assign v_12001 = mux_12001(v_12002);
  assign v_12002 = ~v_11997;
  assign v_12003 = ~v_11578;
  assign v_12004 = v_12005 | v_12006;
  assign v_12005 = mux_12005(v_11580);
  assign v_12006 = mux_12006(v_11991);
  assign v_12008 = v_12009 | v_12420;
  assign v_12009 = act_12010 & 1'h1;
  assign act_12010 = v_12011 | v_12209;
  assign v_12011 = v_12012 & v_12210;
  assign v_12012 = v_12013 & v_12219;
  assign v_12013 = ~v_12014;
  assign v_12015 = v_12016 | v_12203;
  assign v_12016 = act_12017 & 1'h1;
  assign act_12017 = v_12018 | v_12104;
  assign v_12018 = v_12019 & v_12105;
  assign v_12019 = v_12020 & v_12114;
  assign v_12020 = ~v_12021;
  assign v_12022 = v_12023 | v_12098;
  assign v_12023 = act_12024 & 1'h1;
  assign act_12024 = v_12025 | v_12055;
  assign v_12025 = v_12026 & v_12056;
  assign v_12026 = v_12027 & v_12065;
  assign v_12027 = ~v_12028;
  assign v_12029 = v_12030 | v_12049;
  assign v_12030 = act_12031 & 1'h1;
  assign act_12031 = v_12032 | v_12038;
  assign v_12032 = v_12033 & v_12039;
  assign v_12033 = v_12034 & vout_canPeek_12044;
  assign v_12034 = ~vout_canPeek_12035;
  pebbles_core
    pebbles_core_12035
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12036),
       .in0_consume_en(vin0_consume_en_12035),
       .out_canPeek(vout_canPeek_12035),
       .out_peek(vout_peek_12035));
  assign v_12036 = v_12037 | v_12042;
  assign v_12037 = mux_12037(v_12038);
  assign v_12038 = vout_canPeek_12035 & v_12039;
  assign v_12039 = v_12040 & 1'h1;
  assign v_12040 = v_12041 | 1'h0;
  assign v_12041 = ~v_12028;
  assign v_12042 = mux_12042(v_12043);
  assign v_12043 = ~v_12038;
  pebbles_core
    pebbles_core_12044
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12045),
       .in0_consume_en(vin0_consume_en_12044),
       .out_canPeek(vout_canPeek_12044),
       .out_peek(vout_peek_12044));
  assign v_12045 = v_12046 | v_12047;
  assign v_12046 = mux_12046(v_12032);
  assign v_12047 = mux_12047(v_12048);
  assign v_12048 = ~v_12032;
  assign v_12049 = v_12050 & 1'h1;
  assign v_12050 = v_12051 & v_12052;
  assign v_12051 = ~act_12031;
  assign v_12052 = v_12053 | v_12061;
  assign v_12053 = v_12054 | v_12059;
  assign v_12054 = mux_12054(v_12055);
  assign v_12055 = v_12028 & v_12056;
  assign v_12056 = v_12057 & 1'h1;
  assign v_12057 = v_12058 | 1'h0;
  assign v_12058 = ~v_12021;
  assign v_12059 = mux_12059(v_12060);
  assign v_12060 = ~v_12055;
  assign v_12061 = ~v_12028;
  assign v_12062 = v_12063 | v_12064;
  assign v_12063 = mux_12063(v_12030);
  assign v_12064 = mux_12064(v_12049);
  assign v_12066 = v_12067 | v_12086;
  assign v_12067 = act_12068 & 1'h1;
  assign act_12068 = v_12069 | v_12075;
  assign v_12069 = v_12070 & v_12076;
  assign v_12070 = v_12071 & vout_canPeek_12081;
  assign v_12071 = ~vout_canPeek_12072;
  pebbles_core
    pebbles_core_12072
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12073),
       .in0_consume_en(vin0_consume_en_12072),
       .out_canPeek(vout_canPeek_12072),
       .out_peek(vout_peek_12072));
  assign v_12073 = v_12074 | v_12079;
  assign v_12074 = mux_12074(v_12075);
  assign v_12075 = vout_canPeek_12072 & v_12076;
  assign v_12076 = v_12077 & 1'h1;
  assign v_12077 = v_12078 | 1'h0;
  assign v_12078 = ~v_12065;
  assign v_12079 = mux_12079(v_12080);
  assign v_12080 = ~v_12075;
  pebbles_core
    pebbles_core_12081
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12082),
       .in0_consume_en(vin0_consume_en_12081),
       .out_canPeek(vout_canPeek_12081),
       .out_peek(vout_peek_12081));
  assign v_12082 = v_12083 | v_12084;
  assign v_12083 = mux_12083(v_12069);
  assign v_12084 = mux_12084(v_12085);
  assign v_12085 = ~v_12069;
  assign v_12086 = v_12087 & 1'h1;
  assign v_12087 = v_12088 & v_12089;
  assign v_12088 = ~act_12068;
  assign v_12089 = v_12090 | v_12094;
  assign v_12090 = v_12091 | v_12092;
  assign v_12091 = mux_12091(v_12025);
  assign v_12092 = mux_12092(v_12093);
  assign v_12093 = ~v_12025;
  assign v_12094 = ~v_12065;
  assign v_12095 = v_12096 | v_12097;
  assign v_12096 = mux_12096(v_12067);
  assign v_12097 = mux_12097(v_12086);
  assign v_12098 = v_12099 & 1'h1;
  assign v_12099 = v_12100 & v_12101;
  assign v_12100 = ~act_12024;
  assign v_12101 = v_12102 | v_12110;
  assign v_12102 = v_12103 | v_12108;
  assign v_12103 = mux_12103(v_12104);
  assign v_12104 = v_12021 & v_12105;
  assign v_12105 = v_12106 & 1'h1;
  assign v_12106 = v_12107 | 1'h0;
  assign v_12107 = ~v_12014;
  assign v_12108 = mux_12108(v_12109);
  assign v_12109 = ~v_12104;
  assign v_12110 = ~v_12021;
  assign v_12111 = v_12112 | v_12113;
  assign v_12112 = mux_12112(v_12023);
  assign v_12113 = mux_12113(v_12098);
  assign v_12115 = v_12116 | v_12191;
  assign v_12116 = act_12117 & 1'h1;
  assign act_12117 = v_12118 | v_12148;
  assign v_12118 = v_12119 & v_12149;
  assign v_12119 = v_12120 & v_12158;
  assign v_12120 = ~v_12121;
  assign v_12122 = v_12123 | v_12142;
  assign v_12123 = act_12124 & 1'h1;
  assign act_12124 = v_12125 | v_12131;
  assign v_12125 = v_12126 & v_12132;
  assign v_12126 = v_12127 & vout_canPeek_12137;
  assign v_12127 = ~vout_canPeek_12128;
  pebbles_core
    pebbles_core_12128
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12129),
       .in0_consume_en(vin0_consume_en_12128),
       .out_canPeek(vout_canPeek_12128),
       .out_peek(vout_peek_12128));
  assign v_12129 = v_12130 | v_12135;
  assign v_12130 = mux_12130(v_12131);
  assign v_12131 = vout_canPeek_12128 & v_12132;
  assign v_12132 = v_12133 & 1'h1;
  assign v_12133 = v_12134 | 1'h0;
  assign v_12134 = ~v_12121;
  assign v_12135 = mux_12135(v_12136);
  assign v_12136 = ~v_12131;
  pebbles_core
    pebbles_core_12137
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12138),
       .in0_consume_en(vin0_consume_en_12137),
       .out_canPeek(vout_canPeek_12137),
       .out_peek(vout_peek_12137));
  assign v_12138 = v_12139 | v_12140;
  assign v_12139 = mux_12139(v_12125);
  assign v_12140 = mux_12140(v_12141);
  assign v_12141 = ~v_12125;
  assign v_12142 = v_12143 & 1'h1;
  assign v_12143 = v_12144 & v_12145;
  assign v_12144 = ~act_12124;
  assign v_12145 = v_12146 | v_12154;
  assign v_12146 = v_12147 | v_12152;
  assign v_12147 = mux_12147(v_12148);
  assign v_12148 = v_12121 & v_12149;
  assign v_12149 = v_12150 & 1'h1;
  assign v_12150 = v_12151 | 1'h0;
  assign v_12151 = ~v_12114;
  assign v_12152 = mux_12152(v_12153);
  assign v_12153 = ~v_12148;
  assign v_12154 = ~v_12121;
  assign v_12155 = v_12156 | v_12157;
  assign v_12156 = mux_12156(v_12123);
  assign v_12157 = mux_12157(v_12142);
  assign v_12159 = v_12160 | v_12179;
  assign v_12160 = act_12161 & 1'h1;
  assign act_12161 = v_12162 | v_12168;
  assign v_12162 = v_12163 & v_12169;
  assign v_12163 = v_12164 & vout_canPeek_12174;
  assign v_12164 = ~vout_canPeek_12165;
  pebbles_core
    pebbles_core_12165
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12166),
       .in0_consume_en(vin0_consume_en_12165),
       .out_canPeek(vout_canPeek_12165),
       .out_peek(vout_peek_12165));
  assign v_12166 = v_12167 | v_12172;
  assign v_12167 = mux_12167(v_12168);
  assign v_12168 = vout_canPeek_12165 & v_12169;
  assign v_12169 = v_12170 & 1'h1;
  assign v_12170 = v_12171 | 1'h0;
  assign v_12171 = ~v_12158;
  assign v_12172 = mux_12172(v_12173);
  assign v_12173 = ~v_12168;
  pebbles_core
    pebbles_core_12174
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12175),
       .in0_consume_en(vin0_consume_en_12174),
       .out_canPeek(vout_canPeek_12174),
       .out_peek(vout_peek_12174));
  assign v_12175 = v_12176 | v_12177;
  assign v_12176 = mux_12176(v_12162);
  assign v_12177 = mux_12177(v_12178);
  assign v_12178 = ~v_12162;
  assign v_12179 = v_12180 & 1'h1;
  assign v_12180 = v_12181 & v_12182;
  assign v_12181 = ~act_12161;
  assign v_12182 = v_12183 | v_12187;
  assign v_12183 = v_12184 | v_12185;
  assign v_12184 = mux_12184(v_12118);
  assign v_12185 = mux_12185(v_12186);
  assign v_12186 = ~v_12118;
  assign v_12187 = ~v_12158;
  assign v_12188 = v_12189 | v_12190;
  assign v_12189 = mux_12189(v_12160);
  assign v_12190 = mux_12190(v_12179);
  assign v_12191 = v_12192 & 1'h1;
  assign v_12192 = v_12193 & v_12194;
  assign v_12193 = ~act_12117;
  assign v_12194 = v_12195 | v_12199;
  assign v_12195 = v_12196 | v_12197;
  assign v_12196 = mux_12196(v_12018);
  assign v_12197 = mux_12197(v_12198);
  assign v_12198 = ~v_12018;
  assign v_12199 = ~v_12114;
  assign v_12200 = v_12201 | v_12202;
  assign v_12201 = mux_12201(v_12116);
  assign v_12202 = mux_12202(v_12191);
  assign v_12203 = v_12204 & 1'h1;
  assign v_12204 = v_12205 & v_12206;
  assign v_12205 = ~act_12017;
  assign v_12206 = v_12207 | v_12215;
  assign v_12207 = v_12208 | v_12213;
  assign v_12208 = mux_12208(v_12209);
  assign v_12209 = v_12014 & v_12210;
  assign v_12210 = v_12211 & 1'h1;
  assign v_12211 = v_12212 | 1'h0;
  assign v_12212 = ~v_12007;
  assign v_12213 = mux_12213(v_12214);
  assign v_12214 = ~v_12209;
  assign v_12215 = ~v_12014;
  assign v_12216 = v_12217 | v_12218;
  assign v_12217 = mux_12217(v_12016);
  assign v_12218 = mux_12218(v_12203);
  assign v_12220 = v_12221 | v_12408;
  assign v_12221 = act_12222 & 1'h1;
  assign act_12222 = v_12223 | v_12309;
  assign v_12223 = v_12224 & v_12310;
  assign v_12224 = v_12225 & v_12319;
  assign v_12225 = ~v_12226;
  assign v_12227 = v_12228 | v_12303;
  assign v_12228 = act_12229 & 1'h1;
  assign act_12229 = v_12230 | v_12260;
  assign v_12230 = v_12231 & v_12261;
  assign v_12231 = v_12232 & v_12270;
  assign v_12232 = ~v_12233;
  assign v_12234 = v_12235 | v_12254;
  assign v_12235 = act_12236 & 1'h1;
  assign act_12236 = v_12237 | v_12243;
  assign v_12237 = v_12238 & v_12244;
  assign v_12238 = v_12239 & vout_canPeek_12249;
  assign v_12239 = ~vout_canPeek_12240;
  pebbles_core
    pebbles_core_12240
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12241),
       .in0_consume_en(vin0_consume_en_12240),
       .out_canPeek(vout_canPeek_12240),
       .out_peek(vout_peek_12240));
  assign v_12241 = v_12242 | v_12247;
  assign v_12242 = mux_12242(v_12243);
  assign v_12243 = vout_canPeek_12240 & v_12244;
  assign v_12244 = v_12245 & 1'h1;
  assign v_12245 = v_12246 | 1'h0;
  assign v_12246 = ~v_12233;
  assign v_12247 = mux_12247(v_12248);
  assign v_12248 = ~v_12243;
  pebbles_core
    pebbles_core_12249
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12250),
       .in0_consume_en(vin0_consume_en_12249),
       .out_canPeek(vout_canPeek_12249),
       .out_peek(vout_peek_12249));
  assign v_12250 = v_12251 | v_12252;
  assign v_12251 = mux_12251(v_12237);
  assign v_12252 = mux_12252(v_12253);
  assign v_12253 = ~v_12237;
  assign v_12254 = v_12255 & 1'h1;
  assign v_12255 = v_12256 & v_12257;
  assign v_12256 = ~act_12236;
  assign v_12257 = v_12258 | v_12266;
  assign v_12258 = v_12259 | v_12264;
  assign v_12259 = mux_12259(v_12260);
  assign v_12260 = v_12233 & v_12261;
  assign v_12261 = v_12262 & 1'h1;
  assign v_12262 = v_12263 | 1'h0;
  assign v_12263 = ~v_12226;
  assign v_12264 = mux_12264(v_12265);
  assign v_12265 = ~v_12260;
  assign v_12266 = ~v_12233;
  assign v_12267 = v_12268 | v_12269;
  assign v_12268 = mux_12268(v_12235);
  assign v_12269 = mux_12269(v_12254);
  assign v_12271 = v_12272 | v_12291;
  assign v_12272 = act_12273 & 1'h1;
  assign act_12273 = v_12274 | v_12280;
  assign v_12274 = v_12275 & v_12281;
  assign v_12275 = v_12276 & vout_canPeek_12286;
  assign v_12276 = ~vout_canPeek_12277;
  pebbles_core
    pebbles_core_12277
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12278),
       .in0_consume_en(vin0_consume_en_12277),
       .out_canPeek(vout_canPeek_12277),
       .out_peek(vout_peek_12277));
  assign v_12278 = v_12279 | v_12284;
  assign v_12279 = mux_12279(v_12280);
  assign v_12280 = vout_canPeek_12277 & v_12281;
  assign v_12281 = v_12282 & 1'h1;
  assign v_12282 = v_12283 | 1'h0;
  assign v_12283 = ~v_12270;
  assign v_12284 = mux_12284(v_12285);
  assign v_12285 = ~v_12280;
  pebbles_core
    pebbles_core_12286
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12287),
       .in0_consume_en(vin0_consume_en_12286),
       .out_canPeek(vout_canPeek_12286),
       .out_peek(vout_peek_12286));
  assign v_12287 = v_12288 | v_12289;
  assign v_12288 = mux_12288(v_12274);
  assign v_12289 = mux_12289(v_12290);
  assign v_12290 = ~v_12274;
  assign v_12291 = v_12292 & 1'h1;
  assign v_12292 = v_12293 & v_12294;
  assign v_12293 = ~act_12273;
  assign v_12294 = v_12295 | v_12299;
  assign v_12295 = v_12296 | v_12297;
  assign v_12296 = mux_12296(v_12230);
  assign v_12297 = mux_12297(v_12298);
  assign v_12298 = ~v_12230;
  assign v_12299 = ~v_12270;
  assign v_12300 = v_12301 | v_12302;
  assign v_12301 = mux_12301(v_12272);
  assign v_12302 = mux_12302(v_12291);
  assign v_12303 = v_12304 & 1'h1;
  assign v_12304 = v_12305 & v_12306;
  assign v_12305 = ~act_12229;
  assign v_12306 = v_12307 | v_12315;
  assign v_12307 = v_12308 | v_12313;
  assign v_12308 = mux_12308(v_12309);
  assign v_12309 = v_12226 & v_12310;
  assign v_12310 = v_12311 & 1'h1;
  assign v_12311 = v_12312 | 1'h0;
  assign v_12312 = ~v_12219;
  assign v_12313 = mux_12313(v_12314);
  assign v_12314 = ~v_12309;
  assign v_12315 = ~v_12226;
  assign v_12316 = v_12317 | v_12318;
  assign v_12317 = mux_12317(v_12228);
  assign v_12318 = mux_12318(v_12303);
  assign v_12320 = v_12321 | v_12396;
  assign v_12321 = act_12322 & 1'h1;
  assign act_12322 = v_12323 | v_12353;
  assign v_12323 = v_12324 & v_12354;
  assign v_12324 = v_12325 & v_12363;
  assign v_12325 = ~v_12326;
  assign v_12327 = v_12328 | v_12347;
  assign v_12328 = act_12329 & 1'h1;
  assign act_12329 = v_12330 | v_12336;
  assign v_12330 = v_12331 & v_12337;
  assign v_12331 = v_12332 & vout_canPeek_12342;
  assign v_12332 = ~vout_canPeek_12333;
  pebbles_core
    pebbles_core_12333
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12334),
       .in0_consume_en(vin0_consume_en_12333),
       .out_canPeek(vout_canPeek_12333),
       .out_peek(vout_peek_12333));
  assign v_12334 = v_12335 | v_12340;
  assign v_12335 = mux_12335(v_12336);
  assign v_12336 = vout_canPeek_12333 & v_12337;
  assign v_12337 = v_12338 & 1'h1;
  assign v_12338 = v_12339 | 1'h0;
  assign v_12339 = ~v_12326;
  assign v_12340 = mux_12340(v_12341);
  assign v_12341 = ~v_12336;
  pebbles_core
    pebbles_core_12342
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12343),
       .in0_consume_en(vin0_consume_en_12342),
       .out_canPeek(vout_canPeek_12342),
       .out_peek(vout_peek_12342));
  assign v_12343 = v_12344 | v_12345;
  assign v_12344 = mux_12344(v_12330);
  assign v_12345 = mux_12345(v_12346);
  assign v_12346 = ~v_12330;
  assign v_12347 = v_12348 & 1'h1;
  assign v_12348 = v_12349 & v_12350;
  assign v_12349 = ~act_12329;
  assign v_12350 = v_12351 | v_12359;
  assign v_12351 = v_12352 | v_12357;
  assign v_12352 = mux_12352(v_12353);
  assign v_12353 = v_12326 & v_12354;
  assign v_12354 = v_12355 & 1'h1;
  assign v_12355 = v_12356 | 1'h0;
  assign v_12356 = ~v_12319;
  assign v_12357 = mux_12357(v_12358);
  assign v_12358 = ~v_12353;
  assign v_12359 = ~v_12326;
  assign v_12360 = v_12361 | v_12362;
  assign v_12361 = mux_12361(v_12328);
  assign v_12362 = mux_12362(v_12347);
  assign v_12364 = v_12365 | v_12384;
  assign v_12365 = act_12366 & 1'h1;
  assign act_12366 = v_12367 | v_12373;
  assign v_12367 = v_12368 & v_12374;
  assign v_12368 = v_12369 & vout_canPeek_12379;
  assign v_12369 = ~vout_canPeek_12370;
  pebbles_core
    pebbles_core_12370
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12371),
       .in0_consume_en(vin0_consume_en_12370),
       .out_canPeek(vout_canPeek_12370),
       .out_peek(vout_peek_12370));
  assign v_12371 = v_12372 | v_12377;
  assign v_12372 = mux_12372(v_12373);
  assign v_12373 = vout_canPeek_12370 & v_12374;
  assign v_12374 = v_12375 & 1'h1;
  assign v_12375 = v_12376 | 1'h0;
  assign v_12376 = ~v_12363;
  assign v_12377 = mux_12377(v_12378);
  assign v_12378 = ~v_12373;
  pebbles_core
    pebbles_core_12379
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12380),
       .in0_consume_en(vin0_consume_en_12379),
       .out_canPeek(vout_canPeek_12379),
       .out_peek(vout_peek_12379));
  assign v_12380 = v_12381 | v_12382;
  assign v_12381 = mux_12381(v_12367);
  assign v_12382 = mux_12382(v_12383);
  assign v_12383 = ~v_12367;
  assign v_12384 = v_12385 & 1'h1;
  assign v_12385 = v_12386 & v_12387;
  assign v_12386 = ~act_12366;
  assign v_12387 = v_12388 | v_12392;
  assign v_12388 = v_12389 | v_12390;
  assign v_12389 = mux_12389(v_12323);
  assign v_12390 = mux_12390(v_12391);
  assign v_12391 = ~v_12323;
  assign v_12392 = ~v_12363;
  assign v_12393 = v_12394 | v_12395;
  assign v_12394 = mux_12394(v_12365);
  assign v_12395 = mux_12395(v_12384);
  assign v_12396 = v_12397 & 1'h1;
  assign v_12397 = v_12398 & v_12399;
  assign v_12398 = ~act_12322;
  assign v_12399 = v_12400 | v_12404;
  assign v_12400 = v_12401 | v_12402;
  assign v_12401 = mux_12401(v_12223);
  assign v_12402 = mux_12402(v_12403);
  assign v_12403 = ~v_12223;
  assign v_12404 = ~v_12319;
  assign v_12405 = v_12406 | v_12407;
  assign v_12406 = mux_12406(v_12321);
  assign v_12407 = mux_12407(v_12396);
  assign v_12408 = v_12409 & 1'h1;
  assign v_12409 = v_12410 & v_12411;
  assign v_12410 = ~act_12222;
  assign v_12411 = v_12412 | v_12416;
  assign v_12412 = v_12413 | v_12414;
  assign v_12413 = mux_12413(v_12011);
  assign v_12414 = mux_12414(v_12415);
  assign v_12415 = ~v_12011;
  assign v_12416 = ~v_12219;
  assign v_12417 = v_12418 | v_12419;
  assign v_12418 = mux_12418(v_12221);
  assign v_12419 = mux_12419(v_12408);
  assign v_12420 = v_12421 & 1'h1;
  assign v_12421 = v_12422 & v_12423;
  assign v_12422 = ~act_12010;
  assign v_12423 = v_12424 | v_12428;
  assign v_12424 = v_12425 | v_12426;
  assign v_12425 = mux_12425(v_11575);
  assign v_12426 = mux_12426(v_12427);
  assign v_12427 = ~v_11575;
  assign v_12428 = ~v_12007;
  assign v_12429 = v_12430 | v_12431;
  assign v_12430 = mux_12430(v_12009);
  assign v_12431 = mux_12431(v_12420);
  assign v_12432 = v_12433 & 1'h1;
  assign v_12433 = v_12434 & v_12435;
  assign v_12434 = ~act_11574;
  assign v_12435 = v_12436 | v_12444;
  assign v_12436 = v_12437 | v_12442;
  assign v_12437 = mux_12437(v_12438);
  assign v_12438 = v_11571 & v_12439;
  assign v_12439 = v_12440 & 1'h1;
  assign v_12440 = v_12441 | 1'h0;
  assign v_12441 = ~v_11564;
  assign v_12442 = mux_12442(v_12443);
  assign v_12443 = ~v_12438;
  assign v_12444 = ~v_11571;
  assign v_12445 = v_12446 | v_12447;
  assign v_12446 = mux_12446(v_11573);
  assign v_12447 = mux_12447(v_12432);
  assign v_12449 = v_12450 | v_13309;
  assign v_12450 = act_12451 & 1'h1;
  assign act_12451 = v_12452 | v_12874;
  assign v_12452 = v_12453 & v_12875;
  assign v_12453 = v_12454 & v_12884;
  assign v_12454 = ~v_12455;
  assign v_12456 = v_12457 | v_12868;
  assign v_12457 = act_12458 & 1'h1;
  assign act_12458 = v_12459 | v_12657;
  assign v_12459 = v_12460 & v_12658;
  assign v_12460 = v_12461 & v_12667;
  assign v_12461 = ~v_12462;
  assign v_12463 = v_12464 | v_12651;
  assign v_12464 = act_12465 & 1'h1;
  assign act_12465 = v_12466 | v_12552;
  assign v_12466 = v_12467 & v_12553;
  assign v_12467 = v_12468 & v_12562;
  assign v_12468 = ~v_12469;
  assign v_12470 = v_12471 | v_12546;
  assign v_12471 = act_12472 & 1'h1;
  assign act_12472 = v_12473 | v_12503;
  assign v_12473 = v_12474 & v_12504;
  assign v_12474 = v_12475 & v_12513;
  assign v_12475 = ~v_12476;
  assign v_12477 = v_12478 | v_12497;
  assign v_12478 = act_12479 & 1'h1;
  assign act_12479 = v_12480 | v_12486;
  assign v_12480 = v_12481 & v_12487;
  assign v_12481 = v_12482 & vout_canPeek_12492;
  assign v_12482 = ~vout_canPeek_12483;
  pebbles_core
    pebbles_core_12483
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12484),
       .in0_consume_en(vin0_consume_en_12483),
       .out_canPeek(vout_canPeek_12483),
       .out_peek(vout_peek_12483));
  assign v_12484 = v_12485 | v_12490;
  assign v_12485 = mux_12485(v_12486);
  assign v_12486 = vout_canPeek_12483 & v_12487;
  assign v_12487 = v_12488 & 1'h1;
  assign v_12488 = v_12489 | 1'h0;
  assign v_12489 = ~v_12476;
  assign v_12490 = mux_12490(v_12491);
  assign v_12491 = ~v_12486;
  pebbles_core
    pebbles_core_12492
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12493),
       .in0_consume_en(vin0_consume_en_12492),
       .out_canPeek(vout_canPeek_12492),
       .out_peek(vout_peek_12492));
  assign v_12493 = v_12494 | v_12495;
  assign v_12494 = mux_12494(v_12480);
  assign v_12495 = mux_12495(v_12496);
  assign v_12496 = ~v_12480;
  assign v_12497 = v_12498 & 1'h1;
  assign v_12498 = v_12499 & v_12500;
  assign v_12499 = ~act_12479;
  assign v_12500 = v_12501 | v_12509;
  assign v_12501 = v_12502 | v_12507;
  assign v_12502 = mux_12502(v_12503);
  assign v_12503 = v_12476 & v_12504;
  assign v_12504 = v_12505 & 1'h1;
  assign v_12505 = v_12506 | 1'h0;
  assign v_12506 = ~v_12469;
  assign v_12507 = mux_12507(v_12508);
  assign v_12508 = ~v_12503;
  assign v_12509 = ~v_12476;
  assign v_12510 = v_12511 | v_12512;
  assign v_12511 = mux_12511(v_12478);
  assign v_12512 = mux_12512(v_12497);
  assign v_12514 = v_12515 | v_12534;
  assign v_12515 = act_12516 & 1'h1;
  assign act_12516 = v_12517 | v_12523;
  assign v_12517 = v_12518 & v_12524;
  assign v_12518 = v_12519 & vout_canPeek_12529;
  assign v_12519 = ~vout_canPeek_12520;
  pebbles_core
    pebbles_core_12520
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12521),
       .in0_consume_en(vin0_consume_en_12520),
       .out_canPeek(vout_canPeek_12520),
       .out_peek(vout_peek_12520));
  assign v_12521 = v_12522 | v_12527;
  assign v_12522 = mux_12522(v_12523);
  assign v_12523 = vout_canPeek_12520 & v_12524;
  assign v_12524 = v_12525 & 1'h1;
  assign v_12525 = v_12526 | 1'h0;
  assign v_12526 = ~v_12513;
  assign v_12527 = mux_12527(v_12528);
  assign v_12528 = ~v_12523;
  pebbles_core
    pebbles_core_12529
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12530),
       .in0_consume_en(vin0_consume_en_12529),
       .out_canPeek(vout_canPeek_12529),
       .out_peek(vout_peek_12529));
  assign v_12530 = v_12531 | v_12532;
  assign v_12531 = mux_12531(v_12517);
  assign v_12532 = mux_12532(v_12533);
  assign v_12533 = ~v_12517;
  assign v_12534 = v_12535 & 1'h1;
  assign v_12535 = v_12536 & v_12537;
  assign v_12536 = ~act_12516;
  assign v_12537 = v_12538 | v_12542;
  assign v_12538 = v_12539 | v_12540;
  assign v_12539 = mux_12539(v_12473);
  assign v_12540 = mux_12540(v_12541);
  assign v_12541 = ~v_12473;
  assign v_12542 = ~v_12513;
  assign v_12543 = v_12544 | v_12545;
  assign v_12544 = mux_12544(v_12515);
  assign v_12545 = mux_12545(v_12534);
  assign v_12546 = v_12547 & 1'h1;
  assign v_12547 = v_12548 & v_12549;
  assign v_12548 = ~act_12472;
  assign v_12549 = v_12550 | v_12558;
  assign v_12550 = v_12551 | v_12556;
  assign v_12551 = mux_12551(v_12552);
  assign v_12552 = v_12469 & v_12553;
  assign v_12553 = v_12554 & 1'h1;
  assign v_12554 = v_12555 | 1'h0;
  assign v_12555 = ~v_12462;
  assign v_12556 = mux_12556(v_12557);
  assign v_12557 = ~v_12552;
  assign v_12558 = ~v_12469;
  assign v_12559 = v_12560 | v_12561;
  assign v_12560 = mux_12560(v_12471);
  assign v_12561 = mux_12561(v_12546);
  assign v_12563 = v_12564 | v_12639;
  assign v_12564 = act_12565 & 1'h1;
  assign act_12565 = v_12566 | v_12596;
  assign v_12566 = v_12567 & v_12597;
  assign v_12567 = v_12568 & v_12606;
  assign v_12568 = ~v_12569;
  assign v_12570 = v_12571 | v_12590;
  assign v_12571 = act_12572 & 1'h1;
  assign act_12572 = v_12573 | v_12579;
  assign v_12573 = v_12574 & v_12580;
  assign v_12574 = v_12575 & vout_canPeek_12585;
  assign v_12575 = ~vout_canPeek_12576;
  pebbles_core
    pebbles_core_12576
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12577),
       .in0_consume_en(vin0_consume_en_12576),
       .out_canPeek(vout_canPeek_12576),
       .out_peek(vout_peek_12576));
  assign v_12577 = v_12578 | v_12583;
  assign v_12578 = mux_12578(v_12579);
  assign v_12579 = vout_canPeek_12576 & v_12580;
  assign v_12580 = v_12581 & 1'h1;
  assign v_12581 = v_12582 | 1'h0;
  assign v_12582 = ~v_12569;
  assign v_12583 = mux_12583(v_12584);
  assign v_12584 = ~v_12579;
  pebbles_core
    pebbles_core_12585
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12586),
       .in0_consume_en(vin0_consume_en_12585),
       .out_canPeek(vout_canPeek_12585),
       .out_peek(vout_peek_12585));
  assign v_12586 = v_12587 | v_12588;
  assign v_12587 = mux_12587(v_12573);
  assign v_12588 = mux_12588(v_12589);
  assign v_12589 = ~v_12573;
  assign v_12590 = v_12591 & 1'h1;
  assign v_12591 = v_12592 & v_12593;
  assign v_12592 = ~act_12572;
  assign v_12593 = v_12594 | v_12602;
  assign v_12594 = v_12595 | v_12600;
  assign v_12595 = mux_12595(v_12596);
  assign v_12596 = v_12569 & v_12597;
  assign v_12597 = v_12598 & 1'h1;
  assign v_12598 = v_12599 | 1'h0;
  assign v_12599 = ~v_12562;
  assign v_12600 = mux_12600(v_12601);
  assign v_12601 = ~v_12596;
  assign v_12602 = ~v_12569;
  assign v_12603 = v_12604 | v_12605;
  assign v_12604 = mux_12604(v_12571);
  assign v_12605 = mux_12605(v_12590);
  assign v_12607 = v_12608 | v_12627;
  assign v_12608 = act_12609 & 1'h1;
  assign act_12609 = v_12610 | v_12616;
  assign v_12610 = v_12611 & v_12617;
  assign v_12611 = v_12612 & vout_canPeek_12622;
  assign v_12612 = ~vout_canPeek_12613;
  pebbles_core
    pebbles_core_12613
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12614),
       .in0_consume_en(vin0_consume_en_12613),
       .out_canPeek(vout_canPeek_12613),
       .out_peek(vout_peek_12613));
  assign v_12614 = v_12615 | v_12620;
  assign v_12615 = mux_12615(v_12616);
  assign v_12616 = vout_canPeek_12613 & v_12617;
  assign v_12617 = v_12618 & 1'h1;
  assign v_12618 = v_12619 | 1'h0;
  assign v_12619 = ~v_12606;
  assign v_12620 = mux_12620(v_12621);
  assign v_12621 = ~v_12616;
  pebbles_core
    pebbles_core_12622
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12623),
       .in0_consume_en(vin0_consume_en_12622),
       .out_canPeek(vout_canPeek_12622),
       .out_peek(vout_peek_12622));
  assign v_12623 = v_12624 | v_12625;
  assign v_12624 = mux_12624(v_12610);
  assign v_12625 = mux_12625(v_12626);
  assign v_12626 = ~v_12610;
  assign v_12627 = v_12628 & 1'h1;
  assign v_12628 = v_12629 & v_12630;
  assign v_12629 = ~act_12609;
  assign v_12630 = v_12631 | v_12635;
  assign v_12631 = v_12632 | v_12633;
  assign v_12632 = mux_12632(v_12566);
  assign v_12633 = mux_12633(v_12634);
  assign v_12634 = ~v_12566;
  assign v_12635 = ~v_12606;
  assign v_12636 = v_12637 | v_12638;
  assign v_12637 = mux_12637(v_12608);
  assign v_12638 = mux_12638(v_12627);
  assign v_12639 = v_12640 & 1'h1;
  assign v_12640 = v_12641 & v_12642;
  assign v_12641 = ~act_12565;
  assign v_12642 = v_12643 | v_12647;
  assign v_12643 = v_12644 | v_12645;
  assign v_12644 = mux_12644(v_12466);
  assign v_12645 = mux_12645(v_12646);
  assign v_12646 = ~v_12466;
  assign v_12647 = ~v_12562;
  assign v_12648 = v_12649 | v_12650;
  assign v_12649 = mux_12649(v_12564);
  assign v_12650 = mux_12650(v_12639);
  assign v_12651 = v_12652 & 1'h1;
  assign v_12652 = v_12653 & v_12654;
  assign v_12653 = ~act_12465;
  assign v_12654 = v_12655 | v_12663;
  assign v_12655 = v_12656 | v_12661;
  assign v_12656 = mux_12656(v_12657);
  assign v_12657 = v_12462 & v_12658;
  assign v_12658 = v_12659 & 1'h1;
  assign v_12659 = v_12660 | 1'h0;
  assign v_12660 = ~v_12455;
  assign v_12661 = mux_12661(v_12662);
  assign v_12662 = ~v_12657;
  assign v_12663 = ~v_12462;
  assign v_12664 = v_12665 | v_12666;
  assign v_12665 = mux_12665(v_12464);
  assign v_12666 = mux_12666(v_12651);
  assign v_12668 = v_12669 | v_12856;
  assign v_12669 = act_12670 & 1'h1;
  assign act_12670 = v_12671 | v_12757;
  assign v_12671 = v_12672 & v_12758;
  assign v_12672 = v_12673 & v_12767;
  assign v_12673 = ~v_12674;
  assign v_12675 = v_12676 | v_12751;
  assign v_12676 = act_12677 & 1'h1;
  assign act_12677 = v_12678 | v_12708;
  assign v_12678 = v_12679 & v_12709;
  assign v_12679 = v_12680 & v_12718;
  assign v_12680 = ~v_12681;
  assign v_12682 = v_12683 | v_12702;
  assign v_12683 = act_12684 & 1'h1;
  assign act_12684 = v_12685 | v_12691;
  assign v_12685 = v_12686 & v_12692;
  assign v_12686 = v_12687 & vout_canPeek_12697;
  assign v_12687 = ~vout_canPeek_12688;
  pebbles_core
    pebbles_core_12688
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12689),
       .in0_consume_en(vin0_consume_en_12688),
       .out_canPeek(vout_canPeek_12688),
       .out_peek(vout_peek_12688));
  assign v_12689 = v_12690 | v_12695;
  assign v_12690 = mux_12690(v_12691);
  assign v_12691 = vout_canPeek_12688 & v_12692;
  assign v_12692 = v_12693 & 1'h1;
  assign v_12693 = v_12694 | 1'h0;
  assign v_12694 = ~v_12681;
  assign v_12695 = mux_12695(v_12696);
  assign v_12696 = ~v_12691;
  pebbles_core
    pebbles_core_12697
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12698),
       .in0_consume_en(vin0_consume_en_12697),
       .out_canPeek(vout_canPeek_12697),
       .out_peek(vout_peek_12697));
  assign v_12698 = v_12699 | v_12700;
  assign v_12699 = mux_12699(v_12685);
  assign v_12700 = mux_12700(v_12701);
  assign v_12701 = ~v_12685;
  assign v_12702 = v_12703 & 1'h1;
  assign v_12703 = v_12704 & v_12705;
  assign v_12704 = ~act_12684;
  assign v_12705 = v_12706 | v_12714;
  assign v_12706 = v_12707 | v_12712;
  assign v_12707 = mux_12707(v_12708);
  assign v_12708 = v_12681 & v_12709;
  assign v_12709 = v_12710 & 1'h1;
  assign v_12710 = v_12711 | 1'h0;
  assign v_12711 = ~v_12674;
  assign v_12712 = mux_12712(v_12713);
  assign v_12713 = ~v_12708;
  assign v_12714 = ~v_12681;
  assign v_12715 = v_12716 | v_12717;
  assign v_12716 = mux_12716(v_12683);
  assign v_12717 = mux_12717(v_12702);
  assign v_12719 = v_12720 | v_12739;
  assign v_12720 = act_12721 & 1'h1;
  assign act_12721 = v_12722 | v_12728;
  assign v_12722 = v_12723 & v_12729;
  assign v_12723 = v_12724 & vout_canPeek_12734;
  assign v_12724 = ~vout_canPeek_12725;
  pebbles_core
    pebbles_core_12725
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12726),
       .in0_consume_en(vin0_consume_en_12725),
       .out_canPeek(vout_canPeek_12725),
       .out_peek(vout_peek_12725));
  assign v_12726 = v_12727 | v_12732;
  assign v_12727 = mux_12727(v_12728);
  assign v_12728 = vout_canPeek_12725 & v_12729;
  assign v_12729 = v_12730 & 1'h1;
  assign v_12730 = v_12731 | 1'h0;
  assign v_12731 = ~v_12718;
  assign v_12732 = mux_12732(v_12733);
  assign v_12733 = ~v_12728;
  pebbles_core
    pebbles_core_12734
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12735),
       .in0_consume_en(vin0_consume_en_12734),
       .out_canPeek(vout_canPeek_12734),
       .out_peek(vout_peek_12734));
  assign v_12735 = v_12736 | v_12737;
  assign v_12736 = mux_12736(v_12722);
  assign v_12737 = mux_12737(v_12738);
  assign v_12738 = ~v_12722;
  assign v_12739 = v_12740 & 1'h1;
  assign v_12740 = v_12741 & v_12742;
  assign v_12741 = ~act_12721;
  assign v_12742 = v_12743 | v_12747;
  assign v_12743 = v_12744 | v_12745;
  assign v_12744 = mux_12744(v_12678);
  assign v_12745 = mux_12745(v_12746);
  assign v_12746 = ~v_12678;
  assign v_12747 = ~v_12718;
  assign v_12748 = v_12749 | v_12750;
  assign v_12749 = mux_12749(v_12720);
  assign v_12750 = mux_12750(v_12739);
  assign v_12751 = v_12752 & 1'h1;
  assign v_12752 = v_12753 & v_12754;
  assign v_12753 = ~act_12677;
  assign v_12754 = v_12755 | v_12763;
  assign v_12755 = v_12756 | v_12761;
  assign v_12756 = mux_12756(v_12757);
  assign v_12757 = v_12674 & v_12758;
  assign v_12758 = v_12759 & 1'h1;
  assign v_12759 = v_12760 | 1'h0;
  assign v_12760 = ~v_12667;
  assign v_12761 = mux_12761(v_12762);
  assign v_12762 = ~v_12757;
  assign v_12763 = ~v_12674;
  assign v_12764 = v_12765 | v_12766;
  assign v_12765 = mux_12765(v_12676);
  assign v_12766 = mux_12766(v_12751);
  assign v_12768 = v_12769 | v_12844;
  assign v_12769 = act_12770 & 1'h1;
  assign act_12770 = v_12771 | v_12801;
  assign v_12771 = v_12772 & v_12802;
  assign v_12772 = v_12773 & v_12811;
  assign v_12773 = ~v_12774;
  assign v_12775 = v_12776 | v_12795;
  assign v_12776 = act_12777 & 1'h1;
  assign act_12777 = v_12778 | v_12784;
  assign v_12778 = v_12779 & v_12785;
  assign v_12779 = v_12780 & vout_canPeek_12790;
  assign v_12780 = ~vout_canPeek_12781;
  pebbles_core
    pebbles_core_12781
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12782),
       .in0_consume_en(vin0_consume_en_12781),
       .out_canPeek(vout_canPeek_12781),
       .out_peek(vout_peek_12781));
  assign v_12782 = v_12783 | v_12788;
  assign v_12783 = mux_12783(v_12784);
  assign v_12784 = vout_canPeek_12781 & v_12785;
  assign v_12785 = v_12786 & 1'h1;
  assign v_12786 = v_12787 | 1'h0;
  assign v_12787 = ~v_12774;
  assign v_12788 = mux_12788(v_12789);
  assign v_12789 = ~v_12784;
  pebbles_core
    pebbles_core_12790
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12791),
       .in0_consume_en(vin0_consume_en_12790),
       .out_canPeek(vout_canPeek_12790),
       .out_peek(vout_peek_12790));
  assign v_12791 = v_12792 | v_12793;
  assign v_12792 = mux_12792(v_12778);
  assign v_12793 = mux_12793(v_12794);
  assign v_12794 = ~v_12778;
  assign v_12795 = v_12796 & 1'h1;
  assign v_12796 = v_12797 & v_12798;
  assign v_12797 = ~act_12777;
  assign v_12798 = v_12799 | v_12807;
  assign v_12799 = v_12800 | v_12805;
  assign v_12800 = mux_12800(v_12801);
  assign v_12801 = v_12774 & v_12802;
  assign v_12802 = v_12803 & 1'h1;
  assign v_12803 = v_12804 | 1'h0;
  assign v_12804 = ~v_12767;
  assign v_12805 = mux_12805(v_12806);
  assign v_12806 = ~v_12801;
  assign v_12807 = ~v_12774;
  assign v_12808 = v_12809 | v_12810;
  assign v_12809 = mux_12809(v_12776);
  assign v_12810 = mux_12810(v_12795);
  assign v_12812 = v_12813 | v_12832;
  assign v_12813 = act_12814 & 1'h1;
  assign act_12814 = v_12815 | v_12821;
  assign v_12815 = v_12816 & v_12822;
  assign v_12816 = v_12817 & vout_canPeek_12827;
  assign v_12817 = ~vout_canPeek_12818;
  pebbles_core
    pebbles_core_12818
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12819),
       .in0_consume_en(vin0_consume_en_12818),
       .out_canPeek(vout_canPeek_12818),
       .out_peek(vout_peek_12818));
  assign v_12819 = v_12820 | v_12825;
  assign v_12820 = mux_12820(v_12821);
  assign v_12821 = vout_canPeek_12818 & v_12822;
  assign v_12822 = v_12823 & 1'h1;
  assign v_12823 = v_12824 | 1'h0;
  assign v_12824 = ~v_12811;
  assign v_12825 = mux_12825(v_12826);
  assign v_12826 = ~v_12821;
  pebbles_core
    pebbles_core_12827
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12828),
       .in0_consume_en(vin0_consume_en_12827),
       .out_canPeek(vout_canPeek_12827),
       .out_peek(vout_peek_12827));
  assign v_12828 = v_12829 | v_12830;
  assign v_12829 = mux_12829(v_12815);
  assign v_12830 = mux_12830(v_12831);
  assign v_12831 = ~v_12815;
  assign v_12832 = v_12833 & 1'h1;
  assign v_12833 = v_12834 & v_12835;
  assign v_12834 = ~act_12814;
  assign v_12835 = v_12836 | v_12840;
  assign v_12836 = v_12837 | v_12838;
  assign v_12837 = mux_12837(v_12771);
  assign v_12838 = mux_12838(v_12839);
  assign v_12839 = ~v_12771;
  assign v_12840 = ~v_12811;
  assign v_12841 = v_12842 | v_12843;
  assign v_12842 = mux_12842(v_12813);
  assign v_12843 = mux_12843(v_12832);
  assign v_12844 = v_12845 & 1'h1;
  assign v_12845 = v_12846 & v_12847;
  assign v_12846 = ~act_12770;
  assign v_12847 = v_12848 | v_12852;
  assign v_12848 = v_12849 | v_12850;
  assign v_12849 = mux_12849(v_12671);
  assign v_12850 = mux_12850(v_12851);
  assign v_12851 = ~v_12671;
  assign v_12852 = ~v_12767;
  assign v_12853 = v_12854 | v_12855;
  assign v_12854 = mux_12854(v_12769);
  assign v_12855 = mux_12855(v_12844);
  assign v_12856 = v_12857 & 1'h1;
  assign v_12857 = v_12858 & v_12859;
  assign v_12858 = ~act_12670;
  assign v_12859 = v_12860 | v_12864;
  assign v_12860 = v_12861 | v_12862;
  assign v_12861 = mux_12861(v_12459);
  assign v_12862 = mux_12862(v_12863);
  assign v_12863 = ~v_12459;
  assign v_12864 = ~v_12667;
  assign v_12865 = v_12866 | v_12867;
  assign v_12866 = mux_12866(v_12669);
  assign v_12867 = mux_12867(v_12856);
  assign v_12868 = v_12869 & 1'h1;
  assign v_12869 = v_12870 & v_12871;
  assign v_12870 = ~act_12458;
  assign v_12871 = v_12872 | v_12880;
  assign v_12872 = v_12873 | v_12878;
  assign v_12873 = mux_12873(v_12874);
  assign v_12874 = v_12455 & v_12875;
  assign v_12875 = v_12876 & 1'h1;
  assign v_12876 = v_12877 | 1'h0;
  assign v_12877 = ~v_12448;
  assign v_12878 = mux_12878(v_12879);
  assign v_12879 = ~v_12874;
  assign v_12880 = ~v_12455;
  assign v_12881 = v_12882 | v_12883;
  assign v_12882 = mux_12882(v_12457);
  assign v_12883 = mux_12883(v_12868);
  assign v_12885 = v_12886 | v_13297;
  assign v_12886 = act_12887 & 1'h1;
  assign act_12887 = v_12888 | v_13086;
  assign v_12888 = v_12889 & v_13087;
  assign v_12889 = v_12890 & v_13096;
  assign v_12890 = ~v_12891;
  assign v_12892 = v_12893 | v_13080;
  assign v_12893 = act_12894 & 1'h1;
  assign act_12894 = v_12895 | v_12981;
  assign v_12895 = v_12896 & v_12982;
  assign v_12896 = v_12897 & v_12991;
  assign v_12897 = ~v_12898;
  assign v_12899 = v_12900 | v_12975;
  assign v_12900 = act_12901 & 1'h1;
  assign act_12901 = v_12902 | v_12932;
  assign v_12902 = v_12903 & v_12933;
  assign v_12903 = v_12904 & v_12942;
  assign v_12904 = ~v_12905;
  assign v_12906 = v_12907 | v_12926;
  assign v_12907 = act_12908 & 1'h1;
  assign act_12908 = v_12909 | v_12915;
  assign v_12909 = v_12910 & v_12916;
  assign v_12910 = v_12911 & vout_canPeek_12921;
  assign v_12911 = ~vout_canPeek_12912;
  pebbles_core
    pebbles_core_12912
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12913),
       .in0_consume_en(vin0_consume_en_12912),
       .out_canPeek(vout_canPeek_12912),
       .out_peek(vout_peek_12912));
  assign v_12913 = v_12914 | v_12919;
  assign v_12914 = mux_12914(v_12915);
  assign v_12915 = vout_canPeek_12912 & v_12916;
  assign v_12916 = v_12917 & 1'h1;
  assign v_12917 = v_12918 | 1'h0;
  assign v_12918 = ~v_12905;
  assign v_12919 = mux_12919(v_12920);
  assign v_12920 = ~v_12915;
  pebbles_core
    pebbles_core_12921
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12922),
       .in0_consume_en(vin0_consume_en_12921),
       .out_canPeek(vout_canPeek_12921),
       .out_peek(vout_peek_12921));
  assign v_12922 = v_12923 | v_12924;
  assign v_12923 = mux_12923(v_12909);
  assign v_12924 = mux_12924(v_12925);
  assign v_12925 = ~v_12909;
  assign v_12926 = v_12927 & 1'h1;
  assign v_12927 = v_12928 & v_12929;
  assign v_12928 = ~act_12908;
  assign v_12929 = v_12930 | v_12938;
  assign v_12930 = v_12931 | v_12936;
  assign v_12931 = mux_12931(v_12932);
  assign v_12932 = v_12905 & v_12933;
  assign v_12933 = v_12934 & 1'h1;
  assign v_12934 = v_12935 | 1'h0;
  assign v_12935 = ~v_12898;
  assign v_12936 = mux_12936(v_12937);
  assign v_12937 = ~v_12932;
  assign v_12938 = ~v_12905;
  assign v_12939 = v_12940 | v_12941;
  assign v_12940 = mux_12940(v_12907);
  assign v_12941 = mux_12941(v_12926);
  assign v_12943 = v_12944 | v_12963;
  assign v_12944 = act_12945 & 1'h1;
  assign act_12945 = v_12946 | v_12952;
  assign v_12946 = v_12947 & v_12953;
  assign v_12947 = v_12948 & vout_canPeek_12958;
  assign v_12948 = ~vout_canPeek_12949;
  pebbles_core
    pebbles_core_12949
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12950),
       .in0_consume_en(vin0_consume_en_12949),
       .out_canPeek(vout_canPeek_12949),
       .out_peek(vout_peek_12949));
  assign v_12950 = v_12951 | v_12956;
  assign v_12951 = mux_12951(v_12952);
  assign v_12952 = vout_canPeek_12949 & v_12953;
  assign v_12953 = v_12954 & 1'h1;
  assign v_12954 = v_12955 | 1'h0;
  assign v_12955 = ~v_12942;
  assign v_12956 = mux_12956(v_12957);
  assign v_12957 = ~v_12952;
  pebbles_core
    pebbles_core_12958
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_12959),
       .in0_consume_en(vin0_consume_en_12958),
       .out_canPeek(vout_canPeek_12958),
       .out_peek(vout_peek_12958));
  assign v_12959 = v_12960 | v_12961;
  assign v_12960 = mux_12960(v_12946);
  assign v_12961 = mux_12961(v_12962);
  assign v_12962 = ~v_12946;
  assign v_12963 = v_12964 & 1'h1;
  assign v_12964 = v_12965 & v_12966;
  assign v_12965 = ~act_12945;
  assign v_12966 = v_12967 | v_12971;
  assign v_12967 = v_12968 | v_12969;
  assign v_12968 = mux_12968(v_12902);
  assign v_12969 = mux_12969(v_12970);
  assign v_12970 = ~v_12902;
  assign v_12971 = ~v_12942;
  assign v_12972 = v_12973 | v_12974;
  assign v_12973 = mux_12973(v_12944);
  assign v_12974 = mux_12974(v_12963);
  assign v_12975 = v_12976 & 1'h1;
  assign v_12976 = v_12977 & v_12978;
  assign v_12977 = ~act_12901;
  assign v_12978 = v_12979 | v_12987;
  assign v_12979 = v_12980 | v_12985;
  assign v_12980 = mux_12980(v_12981);
  assign v_12981 = v_12898 & v_12982;
  assign v_12982 = v_12983 & 1'h1;
  assign v_12983 = v_12984 | 1'h0;
  assign v_12984 = ~v_12891;
  assign v_12985 = mux_12985(v_12986);
  assign v_12986 = ~v_12981;
  assign v_12987 = ~v_12898;
  assign v_12988 = v_12989 | v_12990;
  assign v_12989 = mux_12989(v_12900);
  assign v_12990 = mux_12990(v_12975);
  assign v_12992 = v_12993 | v_13068;
  assign v_12993 = act_12994 & 1'h1;
  assign act_12994 = v_12995 | v_13025;
  assign v_12995 = v_12996 & v_13026;
  assign v_12996 = v_12997 & v_13035;
  assign v_12997 = ~v_12998;
  assign v_12999 = v_13000 | v_13019;
  assign v_13000 = act_13001 & 1'h1;
  assign act_13001 = v_13002 | v_13008;
  assign v_13002 = v_13003 & v_13009;
  assign v_13003 = v_13004 & vout_canPeek_13014;
  assign v_13004 = ~vout_canPeek_13005;
  pebbles_core
    pebbles_core_13005
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13006),
       .in0_consume_en(vin0_consume_en_13005),
       .out_canPeek(vout_canPeek_13005),
       .out_peek(vout_peek_13005));
  assign v_13006 = v_13007 | v_13012;
  assign v_13007 = mux_13007(v_13008);
  assign v_13008 = vout_canPeek_13005 & v_13009;
  assign v_13009 = v_13010 & 1'h1;
  assign v_13010 = v_13011 | 1'h0;
  assign v_13011 = ~v_12998;
  assign v_13012 = mux_13012(v_13013);
  assign v_13013 = ~v_13008;
  pebbles_core
    pebbles_core_13014
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13015),
       .in0_consume_en(vin0_consume_en_13014),
       .out_canPeek(vout_canPeek_13014),
       .out_peek(vout_peek_13014));
  assign v_13015 = v_13016 | v_13017;
  assign v_13016 = mux_13016(v_13002);
  assign v_13017 = mux_13017(v_13018);
  assign v_13018 = ~v_13002;
  assign v_13019 = v_13020 & 1'h1;
  assign v_13020 = v_13021 & v_13022;
  assign v_13021 = ~act_13001;
  assign v_13022 = v_13023 | v_13031;
  assign v_13023 = v_13024 | v_13029;
  assign v_13024 = mux_13024(v_13025);
  assign v_13025 = v_12998 & v_13026;
  assign v_13026 = v_13027 & 1'h1;
  assign v_13027 = v_13028 | 1'h0;
  assign v_13028 = ~v_12991;
  assign v_13029 = mux_13029(v_13030);
  assign v_13030 = ~v_13025;
  assign v_13031 = ~v_12998;
  assign v_13032 = v_13033 | v_13034;
  assign v_13033 = mux_13033(v_13000);
  assign v_13034 = mux_13034(v_13019);
  assign v_13036 = v_13037 | v_13056;
  assign v_13037 = act_13038 & 1'h1;
  assign act_13038 = v_13039 | v_13045;
  assign v_13039 = v_13040 & v_13046;
  assign v_13040 = v_13041 & vout_canPeek_13051;
  assign v_13041 = ~vout_canPeek_13042;
  pebbles_core
    pebbles_core_13042
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13043),
       .in0_consume_en(vin0_consume_en_13042),
       .out_canPeek(vout_canPeek_13042),
       .out_peek(vout_peek_13042));
  assign v_13043 = v_13044 | v_13049;
  assign v_13044 = mux_13044(v_13045);
  assign v_13045 = vout_canPeek_13042 & v_13046;
  assign v_13046 = v_13047 & 1'h1;
  assign v_13047 = v_13048 | 1'h0;
  assign v_13048 = ~v_13035;
  assign v_13049 = mux_13049(v_13050);
  assign v_13050 = ~v_13045;
  pebbles_core
    pebbles_core_13051
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13052),
       .in0_consume_en(vin0_consume_en_13051),
       .out_canPeek(vout_canPeek_13051),
       .out_peek(vout_peek_13051));
  assign v_13052 = v_13053 | v_13054;
  assign v_13053 = mux_13053(v_13039);
  assign v_13054 = mux_13054(v_13055);
  assign v_13055 = ~v_13039;
  assign v_13056 = v_13057 & 1'h1;
  assign v_13057 = v_13058 & v_13059;
  assign v_13058 = ~act_13038;
  assign v_13059 = v_13060 | v_13064;
  assign v_13060 = v_13061 | v_13062;
  assign v_13061 = mux_13061(v_12995);
  assign v_13062 = mux_13062(v_13063);
  assign v_13063 = ~v_12995;
  assign v_13064 = ~v_13035;
  assign v_13065 = v_13066 | v_13067;
  assign v_13066 = mux_13066(v_13037);
  assign v_13067 = mux_13067(v_13056);
  assign v_13068 = v_13069 & 1'h1;
  assign v_13069 = v_13070 & v_13071;
  assign v_13070 = ~act_12994;
  assign v_13071 = v_13072 | v_13076;
  assign v_13072 = v_13073 | v_13074;
  assign v_13073 = mux_13073(v_12895);
  assign v_13074 = mux_13074(v_13075);
  assign v_13075 = ~v_12895;
  assign v_13076 = ~v_12991;
  assign v_13077 = v_13078 | v_13079;
  assign v_13078 = mux_13078(v_12993);
  assign v_13079 = mux_13079(v_13068);
  assign v_13080 = v_13081 & 1'h1;
  assign v_13081 = v_13082 & v_13083;
  assign v_13082 = ~act_12894;
  assign v_13083 = v_13084 | v_13092;
  assign v_13084 = v_13085 | v_13090;
  assign v_13085 = mux_13085(v_13086);
  assign v_13086 = v_12891 & v_13087;
  assign v_13087 = v_13088 & 1'h1;
  assign v_13088 = v_13089 | 1'h0;
  assign v_13089 = ~v_12884;
  assign v_13090 = mux_13090(v_13091);
  assign v_13091 = ~v_13086;
  assign v_13092 = ~v_12891;
  assign v_13093 = v_13094 | v_13095;
  assign v_13094 = mux_13094(v_12893);
  assign v_13095 = mux_13095(v_13080);
  assign v_13097 = v_13098 | v_13285;
  assign v_13098 = act_13099 & 1'h1;
  assign act_13099 = v_13100 | v_13186;
  assign v_13100 = v_13101 & v_13187;
  assign v_13101 = v_13102 & v_13196;
  assign v_13102 = ~v_13103;
  assign v_13104 = v_13105 | v_13180;
  assign v_13105 = act_13106 & 1'h1;
  assign act_13106 = v_13107 | v_13137;
  assign v_13107 = v_13108 & v_13138;
  assign v_13108 = v_13109 & v_13147;
  assign v_13109 = ~v_13110;
  assign v_13111 = v_13112 | v_13131;
  assign v_13112 = act_13113 & 1'h1;
  assign act_13113 = v_13114 | v_13120;
  assign v_13114 = v_13115 & v_13121;
  assign v_13115 = v_13116 & vout_canPeek_13126;
  assign v_13116 = ~vout_canPeek_13117;
  pebbles_core
    pebbles_core_13117
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13118),
       .in0_consume_en(vin0_consume_en_13117),
       .out_canPeek(vout_canPeek_13117),
       .out_peek(vout_peek_13117));
  assign v_13118 = v_13119 | v_13124;
  assign v_13119 = mux_13119(v_13120);
  assign v_13120 = vout_canPeek_13117 & v_13121;
  assign v_13121 = v_13122 & 1'h1;
  assign v_13122 = v_13123 | 1'h0;
  assign v_13123 = ~v_13110;
  assign v_13124 = mux_13124(v_13125);
  assign v_13125 = ~v_13120;
  pebbles_core
    pebbles_core_13126
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13127),
       .in0_consume_en(vin0_consume_en_13126),
       .out_canPeek(vout_canPeek_13126),
       .out_peek(vout_peek_13126));
  assign v_13127 = v_13128 | v_13129;
  assign v_13128 = mux_13128(v_13114);
  assign v_13129 = mux_13129(v_13130);
  assign v_13130 = ~v_13114;
  assign v_13131 = v_13132 & 1'h1;
  assign v_13132 = v_13133 & v_13134;
  assign v_13133 = ~act_13113;
  assign v_13134 = v_13135 | v_13143;
  assign v_13135 = v_13136 | v_13141;
  assign v_13136 = mux_13136(v_13137);
  assign v_13137 = v_13110 & v_13138;
  assign v_13138 = v_13139 & 1'h1;
  assign v_13139 = v_13140 | 1'h0;
  assign v_13140 = ~v_13103;
  assign v_13141 = mux_13141(v_13142);
  assign v_13142 = ~v_13137;
  assign v_13143 = ~v_13110;
  assign v_13144 = v_13145 | v_13146;
  assign v_13145 = mux_13145(v_13112);
  assign v_13146 = mux_13146(v_13131);
  assign v_13148 = v_13149 | v_13168;
  assign v_13149 = act_13150 & 1'h1;
  assign act_13150 = v_13151 | v_13157;
  assign v_13151 = v_13152 & v_13158;
  assign v_13152 = v_13153 & vout_canPeek_13163;
  assign v_13153 = ~vout_canPeek_13154;
  pebbles_core
    pebbles_core_13154
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13155),
       .in0_consume_en(vin0_consume_en_13154),
       .out_canPeek(vout_canPeek_13154),
       .out_peek(vout_peek_13154));
  assign v_13155 = v_13156 | v_13161;
  assign v_13156 = mux_13156(v_13157);
  assign v_13157 = vout_canPeek_13154 & v_13158;
  assign v_13158 = v_13159 & 1'h1;
  assign v_13159 = v_13160 | 1'h0;
  assign v_13160 = ~v_13147;
  assign v_13161 = mux_13161(v_13162);
  assign v_13162 = ~v_13157;
  pebbles_core
    pebbles_core_13163
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13164),
       .in0_consume_en(vin0_consume_en_13163),
       .out_canPeek(vout_canPeek_13163),
       .out_peek(vout_peek_13163));
  assign v_13164 = v_13165 | v_13166;
  assign v_13165 = mux_13165(v_13151);
  assign v_13166 = mux_13166(v_13167);
  assign v_13167 = ~v_13151;
  assign v_13168 = v_13169 & 1'h1;
  assign v_13169 = v_13170 & v_13171;
  assign v_13170 = ~act_13150;
  assign v_13171 = v_13172 | v_13176;
  assign v_13172 = v_13173 | v_13174;
  assign v_13173 = mux_13173(v_13107);
  assign v_13174 = mux_13174(v_13175);
  assign v_13175 = ~v_13107;
  assign v_13176 = ~v_13147;
  assign v_13177 = v_13178 | v_13179;
  assign v_13178 = mux_13178(v_13149);
  assign v_13179 = mux_13179(v_13168);
  assign v_13180 = v_13181 & 1'h1;
  assign v_13181 = v_13182 & v_13183;
  assign v_13182 = ~act_13106;
  assign v_13183 = v_13184 | v_13192;
  assign v_13184 = v_13185 | v_13190;
  assign v_13185 = mux_13185(v_13186);
  assign v_13186 = v_13103 & v_13187;
  assign v_13187 = v_13188 & 1'h1;
  assign v_13188 = v_13189 | 1'h0;
  assign v_13189 = ~v_13096;
  assign v_13190 = mux_13190(v_13191);
  assign v_13191 = ~v_13186;
  assign v_13192 = ~v_13103;
  assign v_13193 = v_13194 | v_13195;
  assign v_13194 = mux_13194(v_13105);
  assign v_13195 = mux_13195(v_13180);
  assign v_13197 = v_13198 | v_13273;
  assign v_13198 = act_13199 & 1'h1;
  assign act_13199 = v_13200 | v_13230;
  assign v_13200 = v_13201 & v_13231;
  assign v_13201 = v_13202 & v_13240;
  assign v_13202 = ~v_13203;
  assign v_13204 = v_13205 | v_13224;
  assign v_13205 = act_13206 & 1'h1;
  assign act_13206 = v_13207 | v_13213;
  assign v_13207 = v_13208 & v_13214;
  assign v_13208 = v_13209 & vout_canPeek_13219;
  assign v_13209 = ~vout_canPeek_13210;
  pebbles_core
    pebbles_core_13210
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13211),
       .in0_consume_en(vin0_consume_en_13210),
       .out_canPeek(vout_canPeek_13210),
       .out_peek(vout_peek_13210));
  assign v_13211 = v_13212 | v_13217;
  assign v_13212 = mux_13212(v_13213);
  assign v_13213 = vout_canPeek_13210 & v_13214;
  assign v_13214 = v_13215 & 1'h1;
  assign v_13215 = v_13216 | 1'h0;
  assign v_13216 = ~v_13203;
  assign v_13217 = mux_13217(v_13218);
  assign v_13218 = ~v_13213;
  pebbles_core
    pebbles_core_13219
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13220),
       .in0_consume_en(vin0_consume_en_13219),
       .out_canPeek(vout_canPeek_13219),
       .out_peek(vout_peek_13219));
  assign v_13220 = v_13221 | v_13222;
  assign v_13221 = mux_13221(v_13207);
  assign v_13222 = mux_13222(v_13223);
  assign v_13223 = ~v_13207;
  assign v_13224 = v_13225 & 1'h1;
  assign v_13225 = v_13226 & v_13227;
  assign v_13226 = ~act_13206;
  assign v_13227 = v_13228 | v_13236;
  assign v_13228 = v_13229 | v_13234;
  assign v_13229 = mux_13229(v_13230);
  assign v_13230 = v_13203 & v_13231;
  assign v_13231 = v_13232 & 1'h1;
  assign v_13232 = v_13233 | 1'h0;
  assign v_13233 = ~v_13196;
  assign v_13234 = mux_13234(v_13235);
  assign v_13235 = ~v_13230;
  assign v_13236 = ~v_13203;
  assign v_13237 = v_13238 | v_13239;
  assign v_13238 = mux_13238(v_13205);
  assign v_13239 = mux_13239(v_13224);
  assign v_13241 = v_13242 | v_13261;
  assign v_13242 = act_13243 & 1'h1;
  assign act_13243 = v_13244 | v_13250;
  assign v_13244 = v_13245 & v_13251;
  assign v_13245 = v_13246 & vout_canPeek_13256;
  assign v_13246 = ~vout_canPeek_13247;
  pebbles_core
    pebbles_core_13247
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13248),
       .in0_consume_en(vin0_consume_en_13247),
       .out_canPeek(vout_canPeek_13247),
       .out_peek(vout_peek_13247));
  assign v_13248 = v_13249 | v_13254;
  assign v_13249 = mux_13249(v_13250);
  assign v_13250 = vout_canPeek_13247 & v_13251;
  assign v_13251 = v_13252 & 1'h1;
  assign v_13252 = v_13253 | 1'h0;
  assign v_13253 = ~v_13240;
  assign v_13254 = mux_13254(v_13255);
  assign v_13255 = ~v_13250;
  pebbles_core
    pebbles_core_13256
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13257),
       .in0_consume_en(vin0_consume_en_13256),
       .out_canPeek(vout_canPeek_13256),
       .out_peek(vout_peek_13256));
  assign v_13257 = v_13258 | v_13259;
  assign v_13258 = mux_13258(v_13244);
  assign v_13259 = mux_13259(v_13260);
  assign v_13260 = ~v_13244;
  assign v_13261 = v_13262 & 1'h1;
  assign v_13262 = v_13263 & v_13264;
  assign v_13263 = ~act_13243;
  assign v_13264 = v_13265 | v_13269;
  assign v_13265 = v_13266 | v_13267;
  assign v_13266 = mux_13266(v_13200);
  assign v_13267 = mux_13267(v_13268);
  assign v_13268 = ~v_13200;
  assign v_13269 = ~v_13240;
  assign v_13270 = v_13271 | v_13272;
  assign v_13271 = mux_13271(v_13242);
  assign v_13272 = mux_13272(v_13261);
  assign v_13273 = v_13274 & 1'h1;
  assign v_13274 = v_13275 & v_13276;
  assign v_13275 = ~act_13199;
  assign v_13276 = v_13277 | v_13281;
  assign v_13277 = v_13278 | v_13279;
  assign v_13278 = mux_13278(v_13100);
  assign v_13279 = mux_13279(v_13280);
  assign v_13280 = ~v_13100;
  assign v_13281 = ~v_13196;
  assign v_13282 = v_13283 | v_13284;
  assign v_13283 = mux_13283(v_13198);
  assign v_13284 = mux_13284(v_13273);
  assign v_13285 = v_13286 & 1'h1;
  assign v_13286 = v_13287 & v_13288;
  assign v_13287 = ~act_13099;
  assign v_13288 = v_13289 | v_13293;
  assign v_13289 = v_13290 | v_13291;
  assign v_13290 = mux_13290(v_12888);
  assign v_13291 = mux_13291(v_13292);
  assign v_13292 = ~v_12888;
  assign v_13293 = ~v_13096;
  assign v_13294 = v_13295 | v_13296;
  assign v_13295 = mux_13295(v_13098);
  assign v_13296 = mux_13296(v_13285);
  assign v_13297 = v_13298 & 1'h1;
  assign v_13298 = v_13299 & v_13300;
  assign v_13299 = ~act_12887;
  assign v_13300 = v_13301 | v_13305;
  assign v_13301 = v_13302 | v_13303;
  assign v_13302 = mux_13302(v_12452);
  assign v_13303 = mux_13303(v_13304);
  assign v_13304 = ~v_12452;
  assign v_13305 = ~v_12884;
  assign v_13306 = v_13307 | v_13308;
  assign v_13307 = mux_13307(v_12886);
  assign v_13308 = mux_13308(v_13297);
  assign v_13309 = v_13310 & 1'h1;
  assign v_13310 = v_13311 & v_13312;
  assign v_13311 = ~act_12451;
  assign v_13312 = v_13313 | v_13317;
  assign v_13313 = v_13314 | v_13315;
  assign v_13314 = mux_13314(v_11568);
  assign v_13315 = mux_13315(v_13316);
  assign v_13316 = ~v_11568;
  assign v_13317 = ~v_12448;
  assign v_13318 = v_13319 | v_13320;
  assign v_13319 = mux_13319(v_12450);
  assign v_13320 = mux_13320(v_13309);
  assign v_13321 = v_13322 & 1'h1;
  assign v_13322 = v_13323 & v_13324;
  assign v_13323 = ~act_11567;
  assign v_13324 = v_13325 | v_13333;
  assign v_13325 = v_13326 | v_13331;
  assign v_13326 = mux_13326(v_13327);
  assign v_13327 = v_11564 & v_13328;
  assign v_13328 = v_13329 & 1'h1;
  assign v_13329 = v_13330 | 1'h0;
  assign v_13330 = ~v_11557;
  assign v_13331 = mux_13331(v_13332);
  assign v_13332 = ~v_13327;
  assign v_13333 = ~v_11564;
  assign v_13334 = v_13335 | v_13336;
  assign v_13335 = mux_13335(v_11566);
  assign v_13336 = mux_13336(v_13321);
  assign v_13338 = v_13339 | v_15094;
  assign v_13339 = act_13340 & 1'h1;
  assign act_13340 = v_13341 | v_14211;
  assign v_13341 = v_13342 & v_14212;
  assign v_13342 = v_13343 & v_14221;
  assign v_13343 = ~v_13344;
  assign v_13345 = v_13346 | v_14205;
  assign v_13346 = act_13347 & 1'h1;
  assign act_13347 = v_13348 | v_13770;
  assign v_13348 = v_13349 & v_13771;
  assign v_13349 = v_13350 & v_13780;
  assign v_13350 = ~v_13351;
  assign v_13352 = v_13353 | v_13764;
  assign v_13353 = act_13354 & 1'h1;
  assign act_13354 = v_13355 | v_13553;
  assign v_13355 = v_13356 & v_13554;
  assign v_13356 = v_13357 & v_13563;
  assign v_13357 = ~v_13358;
  assign v_13359 = v_13360 | v_13547;
  assign v_13360 = act_13361 & 1'h1;
  assign act_13361 = v_13362 | v_13448;
  assign v_13362 = v_13363 & v_13449;
  assign v_13363 = v_13364 & v_13458;
  assign v_13364 = ~v_13365;
  assign v_13366 = v_13367 | v_13442;
  assign v_13367 = act_13368 & 1'h1;
  assign act_13368 = v_13369 | v_13399;
  assign v_13369 = v_13370 & v_13400;
  assign v_13370 = v_13371 & v_13409;
  assign v_13371 = ~v_13372;
  assign v_13373 = v_13374 | v_13393;
  assign v_13374 = act_13375 & 1'h1;
  assign act_13375 = v_13376 | v_13382;
  assign v_13376 = v_13377 & v_13383;
  assign v_13377 = v_13378 & vout_canPeek_13388;
  assign v_13378 = ~vout_canPeek_13379;
  pebbles_core
    pebbles_core_13379
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13380),
       .in0_consume_en(vin0_consume_en_13379),
       .out_canPeek(vout_canPeek_13379),
       .out_peek(vout_peek_13379));
  assign v_13380 = v_13381 | v_13386;
  assign v_13381 = mux_13381(v_13382);
  assign v_13382 = vout_canPeek_13379 & v_13383;
  assign v_13383 = v_13384 & 1'h1;
  assign v_13384 = v_13385 | 1'h0;
  assign v_13385 = ~v_13372;
  assign v_13386 = mux_13386(v_13387);
  assign v_13387 = ~v_13382;
  pebbles_core
    pebbles_core_13388
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13389),
       .in0_consume_en(vin0_consume_en_13388),
       .out_canPeek(vout_canPeek_13388),
       .out_peek(vout_peek_13388));
  assign v_13389 = v_13390 | v_13391;
  assign v_13390 = mux_13390(v_13376);
  assign v_13391 = mux_13391(v_13392);
  assign v_13392 = ~v_13376;
  assign v_13393 = v_13394 & 1'h1;
  assign v_13394 = v_13395 & v_13396;
  assign v_13395 = ~act_13375;
  assign v_13396 = v_13397 | v_13405;
  assign v_13397 = v_13398 | v_13403;
  assign v_13398 = mux_13398(v_13399);
  assign v_13399 = v_13372 & v_13400;
  assign v_13400 = v_13401 & 1'h1;
  assign v_13401 = v_13402 | 1'h0;
  assign v_13402 = ~v_13365;
  assign v_13403 = mux_13403(v_13404);
  assign v_13404 = ~v_13399;
  assign v_13405 = ~v_13372;
  assign v_13406 = v_13407 | v_13408;
  assign v_13407 = mux_13407(v_13374);
  assign v_13408 = mux_13408(v_13393);
  assign v_13410 = v_13411 | v_13430;
  assign v_13411 = act_13412 & 1'h1;
  assign act_13412 = v_13413 | v_13419;
  assign v_13413 = v_13414 & v_13420;
  assign v_13414 = v_13415 & vout_canPeek_13425;
  assign v_13415 = ~vout_canPeek_13416;
  pebbles_core
    pebbles_core_13416
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13417),
       .in0_consume_en(vin0_consume_en_13416),
       .out_canPeek(vout_canPeek_13416),
       .out_peek(vout_peek_13416));
  assign v_13417 = v_13418 | v_13423;
  assign v_13418 = mux_13418(v_13419);
  assign v_13419 = vout_canPeek_13416 & v_13420;
  assign v_13420 = v_13421 & 1'h1;
  assign v_13421 = v_13422 | 1'h0;
  assign v_13422 = ~v_13409;
  assign v_13423 = mux_13423(v_13424);
  assign v_13424 = ~v_13419;
  pebbles_core
    pebbles_core_13425
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13426),
       .in0_consume_en(vin0_consume_en_13425),
       .out_canPeek(vout_canPeek_13425),
       .out_peek(vout_peek_13425));
  assign v_13426 = v_13427 | v_13428;
  assign v_13427 = mux_13427(v_13413);
  assign v_13428 = mux_13428(v_13429);
  assign v_13429 = ~v_13413;
  assign v_13430 = v_13431 & 1'h1;
  assign v_13431 = v_13432 & v_13433;
  assign v_13432 = ~act_13412;
  assign v_13433 = v_13434 | v_13438;
  assign v_13434 = v_13435 | v_13436;
  assign v_13435 = mux_13435(v_13369);
  assign v_13436 = mux_13436(v_13437);
  assign v_13437 = ~v_13369;
  assign v_13438 = ~v_13409;
  assign v_13439 = v_13440 | v_13441;
  assign v_13440 = mux_13440(v_13411);
  assign v_13441 = mux_13441(v_13430);
  assign v_13442 = v_13443 & 1'h1;
  assign v_13443 = v_13444 & v_13445;
  assign v_13444 = ~act_13368;
  assign v_13445 = v_13446 | v_13454;
  assign v_13446 = v_13447 | v_13452;
  assign v_13447 = mux_13447(v_13448);
  assign v_13448 = v_13365 & v_13449;
  assign v_13449 = v_13450 & 1'h1;
  assign v_13450 = v_13451 | 1'h0;
  assign v_13451 = ~v_13358;
  assign v_13452 = mux_13452(v_13453);
  assign v_13453 = ~v_13448;
  assign v_13454 = ~v_13365;
  assign v_13455 = v_13456 | v_13457;
  assign v_13456 = mux_13456(v_13367);
  assign v_13457 = mux_13457(v_13442);
  assign v_13459 = v_13460 | v_13535;
  assign v_13460 = act_13461 & 1'h1;
  assign act_13461 = v_13462 | v_13492;
  assign v_13462 = v_13463 & v_13493;
  assign v_13463 = v_13464 & v_13502;
  assign v_13464 = ~v_13465;
  assign v_13466 = v_13467 | v_13486;
  assign v_13467 = act_13468 & 1'h1;
  assign act_13468 = v_13469 | v_13475;
  assign v_13469 = v_13470 & v_13476;
  assign v_13470 = v_13471 & vout_canPeek_13481;
  assign v_13471 = ~vout_canPeek_13472;
  pebbles_core
    pebbles_core_13472
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13473),
       .in0_consume_en(vin0_consume_en_13472),
       .out_canPeek(vout_canPeek_13472),
       .out_peek(vout_peek_13472));
  assign v_13473 = v_13474 | v_13479;
  assign v_13474 = mux_13474(v_13475);
  assign v_13475 = vout_canPeek_13472 & v_13476;
  assign v_13476 = v_13477 & 1'h1;
  assign v_13477 = v_13478 | 1'h0;
  assign v_13478 = ~v_13465;
  assign v_13479 = mux_13479(v_13480);
  assign v_13480 = ~v_13475;
  pebbles_core
    pebbles_core_13481
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13482),
       .in0_consume_en(vin0_consume_en_13481),
       .out_canPeek(vout_canPeek_13481),
       .out_peek(vout_peek_13481));
  assign v_13482 = v_13483 | v_13484;
  assign v_13483 = mux_13483(v_13469);
  assign v_13484 = mux_13484(v_13485);
  assign v_13485 = ~v_13469;
  assign v_13486 = v_13487 & 1'h1;
  assign v_13487 = v_13488 & v_13489;
  assign v_13488 = ~act_13468;
  assign v_13489 = v_13490 | v_13498;
  assign v_13490 = v_13491 | v_13496;
  assign v_13491 = mux_13491(v_13492);
  assign v_13492 = v_13465 & v_13493;
  assign v_13493 = v_13494 & 1'h1;
  assign v_13494 = v_13495 | 1'h0;
  assign v_13495 = ~v_13458;
  assign v_13496 = mux_13496(v_13497);
  assign v_13497 = ~v_13492;
  assign v_13498 = ~v_13465;
  assign v_13499 = v_13500 | v_13501;
  assign v_13500 = mux_13500(v_13467);
  assign v_13501 = mux_13501(v_13486);
  assign v_13503 = v_13504 | v_13523;
  assign v_13504 = act_13505 & 1'h1;
  assign act_13505 = v_13506 | v_13512;
  assign v_13506 = v_13507 & v_13513;
  assign v_13507 = v_13508 & vout_canPeek_13518;
  assign v_13508 = ~vout_canPeek_13509;
  pebbles_core
    pebbles_core_13509
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13510),
       .in0_consume_en(vin0_consume_en_13509),
       .out_canPeek(vout_canPeek_13509),
       .out_peek(vout_peek_13509));
  assign v_13510 = v_13511 | v_13516;
  assign v_13511 = mux_13511(v_13512);
  assign v_13512 = vout_canPeek_13509 & v_13513;
  assign v_13513 = v_13514 & 1'h1;
  assign v_13514 = v_13515 | 1'h0;
  assign v_13515 = ~v_13502;
  assign v_13516 = mux_13516(v_13517);
  assign v_13517 = ~v_13512;
  pebbles_core
    pebbles_core_13518
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13519),
       .in0_consume_en(vin0_consume_en_13518),
       .out_canPeek(vout_canPeek_13518),
       .out_peek(vout_peek_13518));
  assign v_13519 = v_13520 | v_13521;
  assign v_13520 = mux_13520(v_13506);
  assign v_13521 = mux_13521(v_13522);
  assign v_13522 = ~v_13506;
  assign v_13523 = v_13524 & 1'h1;
  assign v_13524 = v_13525 & v_13526;
  assign v_13525 = ~act_13505;
  assign v_13526 = v_13527 | v_13531;
  assign v_13527 = v_13528 | v_13529;
  assign v_13528 = mux_13528(v_13462);
  assign v_13529 = mux_13529(v_13530);
  assign v_13530 = ~v_13462;
  assign v_13531 = ~v_13502;
  assign v_13532 = v_13533 | v_13534;
  assign v_13533 = mux_13533(v_13504);
  assign v_13534 = mux_13534(v_13523);
  assign v_13535 = v_13536 & 1'h1;
  assign v_13536 = v_13537 & v_13538;
  assign v_13537 = ~act_13461;
  assign v_13538 = v_13539 | v_13543;
  assign v_13539 = v_13540 | v_13541;
  assign v_13540 = mux_13540(v_13362);
  assign v_13541 = mux_13541(v_13542);
  assign v_13542 = ~v_13362;
  assign v_13543 = ~v_13458;
  assign v_13544 = v_13545 | v_13546;
  assign v_13545 = mux_13545(v_13460);
  assign v_13546 = mux_13546(v_13535);
  assign v_13547 = v_13548 & 1'h1;
  assign v_13548 = v_13549 & v_13550;
  assign v_13549 = ~act_13361;
  assign v_13550 = v_13551 | v_13559;
  assign v_13551 = v_13552 | v_13557;
  assign v_13552 = mux_13552(v_13553);
  assign v_13553 = v_13358 & v_13554;
  assign v_13554 = v_13555 & 1'h1;
  assign v_13555 = v_13556 | 1'h0;
  assign v_13556 = ~v_13351;
  assign v_13557 = mux_13557(v_13558);
  assign v_13558 = ~v_13553;
  assign v_13559 = ~v_13358;
  assign v_13560 = v_13561 | v_13562;
  assign v_13561 = mux_13561(v_13360);
  assign v_13562 = mux_13562(v_13547);
  assign v_13564 = v_13565 | v_13752;
  assign v_13565 = act_13566 & 1'h1;
  assign act_13566 = v_13567 | v_13653;
  assign v_13567 = v_13568 & v_13654;
  assign v_13568 = v_13569 & v_13663;
  assign v_13569 = ~v_13570;
  assign v_13571 = v_13572 | v_13647;
  assign v_13572 = act_13573 & 1'h1;
  assign act_13573 = v_13574 | v_13604;
  assign v_13574 = v_13575 & v_13605;
  assign v_13575 = v_13576 & v_13614;
  assign v_13576 = ~v_13577;
  assign v_13578 = v_13579 | v_13598;
  assign v_13579 = act_13580 & 1'h1;
  assign act_13580 = v_13581 | v_13587;
  assign v_13581 = v_13582 & v_13588;
  assign v_13582 = v_13583 & vout_canPeek_13593;
  assign v_13583 = ~vout_canPeek_13584;
  pebbles_core
    pebbles_core_13584
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13585),
       .in0_consume_en(vin0_consume_en_13584),
       .out_canPeek(vout_canPeek_13584),
       .out_peek(vout_peek_13584));
  assign v_13585 = v_13586 | v_13591;
  assign v_13586 = mux_13586(v_13587);
  assign v_13587 = vout_canPeek_13584 & v_13588;
  assign v_13588 = v_13589 & 1'h1;
  assign v_13589 = v_13590 | 1'h0;
  assign v_13590 = ~v_13577;
  assign v_13591 = mux_13591(v_13592);
  assign v_13592 = ~v_13587;
  pebbles_core
    pebbles_core_13593
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13594),
       .in0_consume_en(vin0_consume_en_13593),
       .out_canPeek(vout_canPeek_13593),
       .out_peek(vout_peek_13593));
  assign v_13594 = v_13595 | v_13596;
  assign v_13595 = mux_13595(v_13581);
  assign v_13596 = mux_13596(v_13597);
  assign v_13597 = ~v_13581;
  assign v_13598 = v_13599 & 1'h1;
  assign v_13599 = v_13600 & v_13601;
  assign v_13600 = ~act_13580;
  assign v_13601 = v_13602 | v_13610;
  assign v_13602 = v_13603 | v_13608;
  assign v_13603 = mux_13603(v_13604);
  assign v_13604 = v_13577 & v_13605;
  assign v_13605 = v_13606 & 1'h1;
  assign v_13606 = v_13607 | 1'h0;
  assign v_13607 = ~v_13570;
  assign v_13608 = mux_13608(v_13609);
  assign v_13609 = ~v_13604;
  assign v_13610 = ~v_13577;
  assign v_13611 = v_13612 | v_13613;
  assign v_13612 = mux_13612(v_13579);
  assign v_13613 = mux_13613(v_13598);
  assign v_13615 = v_13616 | v_13635;
  assign v_13616 = act_13617 & 1'h1;
  assign act_13617 = v_13618 | v_13624;
  assign v_13618 = v_13619 & v_13625;
  assign v_13619 = v_13620 & vout_canPeek_13630;
  assign v_13620 = ~vout_canPeek_13621;
  pebbles_core
    pebbles_core_13621
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13622),
       .in0_consume_en(vin0_consume_en_13621),
       .out_canPeek(vout_canPeek_13621),
       .out_peek(vout_peek_13621));
  assign v_13622 = v_13623 | v_13628;
  assign v_13623 = mux_13623(v_13624);
  assign v_13624 = vout_canPeek_13621 & v_13625;
  assign v_13625 = v_13626 & 1'h1;
  assign v_13626 = v_13627 | 1'h0;
  assign v_13627 = ~v_13614;
  assign v_13628 = mux_13628(v_13629);
  assign v_13629 = ~v_13624;
  pebbles_core
    pebbles_core_13630
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13631),
       .in0_consume_en(vin0_consume_en_13630),
       .out_canPeek(vout_canPeek_13630),
       .out_peek(vout_peek_13630));
  assign v_13631 = v_13632 | v_13633;
  assign v_13632 = mux_13632(v_13618);
  assign v_13633 = mux_13633(v_13634);
  assign v_13634 = ~v_13618;
  assign v_13635 = v_13636 & 1'h1;
  assign v_13636 = v_13637 & v_13638;
  assign v_13637 = ~act_13617;
  assign v_13638 = v_13639 | v_13643;
  assign v_13639 = v_13640 | v_13641;
  assign v_13640 = mux_13640(v_13574);
  assign v_13641 = mux_13641(v_13642);
  assign v_13642 = ~v_13574;
  assign v_13643 = ~v_13614;
  assign v_13644 = v_13645 | v_13646;
  assign v_13645 = mux_13645(v_13616);
  assign v_13646 = mux_13646(v_13635);
  assign v_13647 = v_13648 & 1'h1;
  assign v_13648 = v_13649 & v_13650;
  assign v_13649 = ~act_13573;
  assign v_13650 = v_13651 | v_13659;
  assign v_13651 = v_13652 | v_13657;
  assign v_13652 = mux_13652(v_13653);
  assign v_13653 = v_13570 & v_13654;
  assign v_13654 = v_13655 & 1'h1;
  assign v_13655 = v_13656 | 1'h0;
  assign v_13656 = ~v_13563;
  assign v_13657 = mux_13657(v_13658);
  assign v_13658 = ~v_13653;
  assign v_13659 = ~v_13570;
  assign v_13660 = v_13661 | v_13662;
  assign v_13661 = mux_13661(v_13572);
  assign v_13662 = mux_13662(v_13647);
  assign v_13664 = v_13665 | v_13740;
  assign v_13665 = act_13666 & 1'h1;
  assign act_13666 = v_13667 | v_13697;
  assign v_13667 = v_13668 & v_13698;
  assign v_13668 = v_13669 & v_13707;
  assign v_13669 = ~v_13670;
  assign v_13671 = v_13672 | v_13691;
  assign v_13672 = act_13673 & 1'h1;
  assign act_13673 = v_13674 | v_13680;
  assign v_13674 = v_13675 & v_13681;
  assign v_13675 = v_13676 & vout_canPeek_13686;
  assign v_13676 = ~vout_canPeek_13677;
  pebbles_core
    pebbles_core_13677
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13678),
       .in0_consume_en(vin0_consume_en_13677),
       .out_canPeek(vout_canPeek_13677),
       .out_peek(vout_peek_13677));
  assign v_13678 = v_13679 | v_13684;
  assign v_13679 = mux_13679(v_13680);
  assign v_13680 = vout_canPeek_13677 & v_13681;
  assign v_13681 = v_13682 & 1'h1;
  assign v_13682 = v_13683 | 1'h0;
  assign v_13683 = ~v_13670;
  assign v_13684 = mux_13684(v_13685);
  assign v_13685 = ~v_13680;
  pebbles_core
    pebbles_core_13686
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13687),
       .in0_consume_en(vin0_consume_en_13686),
       .out_canPeek(vout_canPeek_13686),
       .out_peek(vout_peek_13686));
  assign v_13687 = v_13688 | v_13689;
  assign v_13688 = mux_13688(v_13674);
  assign v_13689 = mux_13689(v_13690);
  assign v_13690 = ~v_13674;
  assign v_13691 = v_13692 & 1'h1;
  assign v_13692 = v_13693 & v_13694;
  assign v_13693 = ~act_13673;
  assign v_13694 = v_13695 | v_13703;
  assign v_13695 = v_13696 | v_13701;
  assign v_13696 = mux_13696(v_13697);
  assign v_13697 = v_13670 & v_13698;
  assign v_13698 = v_13699 & 1'h1;
  assign v_13699 = v_13700 | 1'h0;
  assign v_13700 = ~v_13663;
  assign v_13701 = mux_13701(v_13702);
  assign v_13702 = ~v_13697;
  assign v_13703 = ~v_13670;
  assign v_13704 = v_13705 | v_13706;
  assign v_13705 = mux_13705(v_13672);
  assign v_13706 = mux_13706(v_13691);
  assign v_13708 = v_13709 | v_13728;
  assign v_13709 = act_13710 & 1'h1;
  assign act_13710 = v_13711 | v_13717;
  assign v_13711 = v_13712 & v_13718;
  assign v_13712 = v_13713 & vout_canPeek_13723;
  assign v_13713 = ~vout_canPeek_13714;
  pebbles_core
    pebbles_core_13714
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13715),
       .in0_consume_en(vin0_consume_en_13714),
       .out_canPeek(vout_canPeek_13714),
       .out_peek(vout_peek_13714));
  assign v_13715 = v_13716 | v_13721;
  assign v_13716 = mux_13716(v_13717);
  assign v_13717 = vout_canPeek_13714 & v_13718;
  assign v_13718 = v_13719 & 1'h1;
  assign v_13719 = v_13720 | 1'h0;
  assign v_13720 = ~v_13707;
  assign v_13721 = mux_13721(v_13722);
  assign v_13722 = ~v_13717;
  pebbles_core
    pebbles_core_13723
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13724),
       .in0_consume_en(vin0_consume_en_13723),
       .out_canPeek(vout_canPeek_13723),
       .out_peek(vout_peek_13723));
  assign v_13724 = v_13725 | v_13726;
  assign v_13725 = mux_13725(v_13711);
  assign v_13726 = mux_13726(v_13727);
  assign v_13727 = ~v_13711;
  assign v_13728 = v_13729 & 1'h1;
  assign v_13729 = v_13730 & v_13731;
  assign v_13730 = ~act_13710;
  assign v_13731 = v_13732 | v_13736;
  assign v_13732 = v_13733 | v_13734;
  assign v_13733 = mux_13733(v_13667);
  assign v_13734 = mux_13734(v_13735);
  assign v_13735 = ~v_13667;
  assign v_13736 = ~v_13707;
  assign v_13737 = v_13738 | v_13739;
  assign v_13738 = mux_13738(v_13709);
  assign v_13739 = mux_13739(v_13728);
  assign v_13740 = v_13741 & 1'h1;
  assign v_13741 = v_13742 & v_13743;
  assign v_13742 = ~act_13666;
  assign v_13743 = v_13744 | v_13748;
  assign v_13744 = v_13745 | v_13746;
  assign v_13745 = mux_13745(v_13567);
  assign v_13746 = mux_13746(v_13747);
  assign v_13747 = ~v_13567;
  assign v_13748 = ~v_13663;
  assign v_13749 = v_13750 | v_13751;
  assign v_13750 = mux_13750(v_13665);
  assign v_13751 = mux_13751(v_13740);
  assign v_13752 = v_13753 & 1'h1;
  assign v_13753 = v_13754 & v_13755;
  assign v_13754 = ~act_13566;
  assign v_13755 = v_13756 | v_13760;
  assign v_13756 = v_13757 | v_13758;
  assign v_13757 = mux_13757(v_13355);
  assign v_13758 = mux_13758(v_13759);
  assign v_13759 = ~v_13355;
  assign v_13760 = ~v_13563;
  assign v_13761 = v_13762 | v_13763;
  assign v_13762 = mux_13762(v_13565);
  assign v_13763 = mux_13763(v_13752);
  assign v_13764 = v_13765 & 1'h1;
  assign v_13765 = v_13766 & v_13767;
  assign v_13766 = ~act_13354;
  assign v_13767 = v_13768 | v_13776;
  assign v_13768 = v_13769 | v_13774;
  assign v_13769 = mux_13769(v_13770);
  assign v_13770 = v_13351 & v_13771;
  assign v_13771 = v_13772 & 1'h1;
  assign v_13772 = v_13773 | 1'h0;
  assign v_13773 = ~v_13344;
  assign v_13774 = mux_13774(v_13775);
  assign v_13775 = ~v_13770;
  assign v_13776 = ~v_13351;
  assign v_13777 = v_13778 | v_13779;
  assign v_13778 = mux_13778(v_13353);
  assign v_13779 = mux_13779(v_13764);
  assign v_13781 = v_13782 | v_14193;
  assign v_13782 = act_13783 & 1'h1;
  assign act_13783 = v_13784 | v_13982;
  assign v_13784 = v_13785 & v_13983;
  assign v_13785 = v_13786 & v_13992;
  assign v_13786 = ~v_13787;
  assign v_13788 = v_13789 | v_13976;
  assign v_13789 = act_13790 & 1'h1;
  assign act_13790 = v_13791 | v_13877;
  assign v_13791 = v_13792 & v_13878;
  assign v_13792 = v_13793 & v_13887;
  assign v_13793 = ~v_13794;
  assign v_13795 = v_13796 | v_13871;
  assign v_13796 = act_13797 & 1'h1;
  assign act_13797 = v_13798 | v_13828;
  assign v_13798 = v_13799 & v_13829;
  assign v_13799 = v_13800 & v_13838;
  assign v_13800 = ~v_13801;
  assign v_13802 = v_13803 | v_13822;
  assign v_13803 = act_13804 & 1'h1;
  assign act_13804 = v_13805 | v_13811;
  assign v_13805 = v_13806 & v_13812;
  assign v_13806 = v_13807 & vout_canPeek_13817;
  assign v_13807 = ~vout_canPeek_13808;
  pebbles_core
    pebbles_core_13808
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13809),
       .in0_consume_en(vin0_consume_en_13808),
       .out_canPeek(vout_canPeek_13808),
       .out_peek(vout_peek_13808));
  assign v_13809 = v_13810 | v_13815;
  assign v_13810 = mux_13810(v_13811);
  assign v_13811 = vout_canPeek_13808 & v_13812;
  assign v_13812 = v_13813 & 1'h1;
  assign v_13813 = v_13814 | 1'h0;
  assign v_13814 = ~v_13801;
  assign v_13815 = mux_13815(v_13816);
  assign v_13816 = ~v_13811;
  pebbles_core
    pebbles_core_13817
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13818),
       .in0_consume_en(vin0_consume_en_13817),
       .out_canPeek(vout_canPeek_13817),
       .out_peek(vout_peek_13817));
  assign v_13818 = v_13819 | v_13820;
  assign v_13819 = mux_13819(v_13805);
  assign v_13820 = mux_13820(v_13821);
  assign v_13821 = ~v_13805;
  assign v_13822 = v_13823 & 1'h1;
  assign v_13823 = v_13824 & v_13825;
  assign v_13824 = ~act_13804;
  assign v_13825 = v_13826 | v_13834;
  assign v_13826 = v_13827 | v_13832;
  assign v_13827 = mux_13827(v_13828);
  assign v_13828 = v_13801 & v_13829;
  assign v_13829 = v_13830 & 1'h1;
  assign v_13830 = v_13831 | 1'h0;
  assign v_13831 = ~v_13794;
  assign v_13832 = mux_13832(v_13833);
  assign v_13833 = ~v_13828;
  assign v_13834 = ~v_13801;
  assign v_13835 = v_13836 | v_13837;
  assign v_13836 = mux_13836(v_13803);
  assign v_13837 = mux_13837(v_13822);
  assign v_13839 = v_13840 | v_13859;
  assign v_13840 = act_13841 & 1'h1;
  assign act_13841 = v_13842 | v_13848;
  assign v_13842 = v_13843 & v_13849;
  assign v_13843 = v_13844 & vout_canPeek_13854;
  assign v_13844 = ~vout_canPeek_13845;
  pebbles_core
    pebbles_core_13845
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13846),
       .in0_consume_en(vin0_consume_en_13845),
       .out_canPeek(vout_canPeek_13845),
       .out_peek(vout_peek_13845));
  assign v_13846 = v_13847 | v_13852;
  assign v_13847 = mux_13847(v_13848);
  assign v_13848 = vout_canPeek_13845 & v_13849;
  assign v_13849 = v_13850 & 1'h1;
  assign v_13850 = v_13851 | 1'h0;
  assign v_13851 = ~v_13838;
  assign v_13852 = mux_13852(v_13853);
  assign v_13853 = ~v_13848;
  pebbles_core
    pebbles_core_13854
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13855),
       .in0_consume_en(vin0_consume_en_13854),
       .out_canPeek(vout_canPeek_13854),
       .out_peek(vout_peek_13854));
  assign v_13855 = v_13856 | v_13857;
  assign v_13856 = mux_13856(v_13842);
  assign v_13857 = mux_13857(v_13858);
  assign v_13858 = ~v_13842;
  assign v_13859 = v_13860 & 1'h1;
  assign v_13860 = v_13861 & v_13862;
  assign v_13861 = ~act_13841;
  assign v_13862 = v_13863 | v_13867;
  assign v_13863 = v_13864 | v_13865;
  assign v_13864 = mux_13864(v_13798);
  assign v_13865 = mux_13865(v_13866);
  assign v_13866 = ~v_13798;
  assign v_13867 = ~v_13838;
  assign v_13868 = v_13869 | v_13870;
  assign v_13869 = mux_13869(v_13840);
  assign v_13870 = mux_13870(v_13859);
  assign v_13871 = v_13872 & 1'h1;
  assign v_13872 = v_13873 & v_13874;
  assign v_13873 = ~act_13797;
  assign v_13874 = v_13875 | v_13883;
  assign v_13875 = v_13876 | v_13881;
  assign v_13876 = mux_13876(v_13877);
  assign v_13877 = v_13794 & v_13878;
  assign v_13878 = v_13879 & 1'h1;
  assign v_13879 = v_13880 | 1'h0;
  assign v_13880 = ~v_13787;
  assign v_13881 = mux_13881(v_13882);
  assign v_13882 = ~v_13877;
  assign v_13883 = ~v_13794;
  assign v_13884 = v_13885 | v_13886;
  assign v_13885 = mux_13885(v_13796);
  assign v_13886 = mux_13886(v_13871);
  assign v_13888 = v_13889 | v_13964;
  assign v_13889 = act_13890 & 1'h1;
  assign act_13890 = v_13891 | v_13921;
  assign v_13891 = v_13892 & v_13922;
  assign v_13892 = v_13893 & v_13931;
  assign v_13893 = ~v_13894;
  assign v_13895 = v_13896 | v_13915;
  assign v_13896 = act_13897 & 1'h1;
  assign act_13897 = v_13898 | v_13904;
  assign v_13898 = v_13899 & v_13905;
  assign v_13899 = v_13900 & vout_canPeek_13910;
  assign v_13900 = ~vout_canPeek_13901;
  pebbles_core
    pebbles_core_13901
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13902),
       .in0_consume_en(vin0_consume_en_13901),
       .out_canPeek(vout_canPeek_13901),
       .out_peek(vout_peek_13901));
  assign v_13902 = v_13903 | v_13908;
  assign v_13903 = mux_13903(v_13904);
  assign v_13904 = vout_canPeek_13901 & v_13905;
  assign v_13905 = v_13906 & 1'h1;
  assign v_13906 = v_13907 | 1'h0;
  assign v_13907 = ~v_13894;
  assign v_13908 = mux_13908(v_13909);
  assign v_13909 = ~v_13904;
  pebbles_core
    pebbles_core_13910
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13911),
       .in0_consume_en(vin0_consume_en_13910),
       .out_canPeek(vout_canPeek_13910),
       .out_peek(vout_peek_13910));
  assign v_13911 = v_13912 | v_13913;
  assign v_13912 = mux_13912(v_13898);
  assign v_13913 = mux_13913(v_13914);
  assign v_13914 = ~v_13898;
  assign v_13915 = v_13916 & 1'h1;
  assign v_13916 = v_13917 & v_13918;
  assign v_13917 = ~act_13897;
  assign v_13918 = v_13919 | v_13927;
  assign v_13919 = v_13920 | v_13925;
  assign v_13920 = mux_13920(v_13921);
  assign v_13921 = v_13894 & v_13922;
  assign v_13922 = v_13923 & 1'h1;
  assign v_13923 = v_13924 | 1'h0;
  assign v_13924 = ~v_13887;
  assign v_13925 = mux_13925(v_13926);
  assign v_13926 = ~v_13921;
  assign v_13927 = ~v_13894;
  assign v_13928 = v_13929 | v_13930;
  assign v_13929 = mux_13929(v_13896);
  assign v_13930 = mux_13930(v_13915);
  assign v_13932 = v_13933 | v_13952;
  assign v_13933 = act_13934 & 1'h1;
  assign act_13934 = v_13935 | v_13941;
  assign v_13935 = v_13936 & v_13942;
  assign v_13936 = v_13937 & vout_canPeek_13947;
  assign v_13937 = ~vout_canPeek_13938;
  pebbles_core
    pebbles_core_13938
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13939),
       .in0_consume_en(vin0_consume_en_13938),
       .out_canPeek(vout_canPeek_13938),
       .out_peek(vout_peek_13938));
  assign v_13939 = v_13940 | v_13945;
  assign v_13940 = mux_13940(v_13941);
  assign v_13941 = vout_canPeek_13938 & v_13942;
  assign v_13942 = v_13943 & 1'h1;
  assign v_13943 = v_13944 | 1'h0;
  assign v_13944 = ~v_13931;
  assign v_13945 = mux_13945(v_13946);
  assign v_13946 = ~v_13941;
  pebbles_core
    pebbles_core_13947
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_13948),
       .in0_consume_en(vin0_consume_en_13947),
       .out_canPeek(vout_canPeek_13947),
       .out_peek(vout_peek_13947));
  assign v_13948 = v_13949 | v_13950;
  assign v_13949 = mux_13949(v_13935);
  assign v_13950 = mux_13950(v_13951);
  assign v_13951 = ~v_13935;
  assign v_13952 = v_13953 & 1'h1;
  assign v_13953 = v_13954 & v_13955;
  assign v_13954 = ~act_13934;
  assign v_13955 = v_13956 | v_13960;
  assign v_13956 = v_13957 | v_13958;
  assign v_13957 = mux_13957(v_13891);
  assign v_13958 = mux_13958(v_13959);
  assign v_13959 = ~v_13891;
  assign v_13960 = ~v_13931;
  assign v_13961 = v_13962 | v_13963;
  assign v_13962 = mux_13962(v_13933);
  assign v_13963 = mux_13963(v_13952);
  assign v_13964 = v_13965 & 1'h1;
  assign v_13965 = v_13966 & v_13967;
  assign v_13966 = ~act_13890;
  assign v_13967 = v_13968 | v_13972;
  assign v_13968 = v_13969 | v_13970;
  assign v_13969 = mux_13969(v_13791);
  assign v_13970 = mux_13970(v_13971);
  assign v_13971 = ~v_13791;
  assign v_13972 = ~v_13887;
  assign v_13973 = v_13974 | v_13975;
  assign v_13974 = mux_13974(v_13889);
  assign v_13975 = mux_13975(v_13964);
  assign v_13976 = v_13977 & 1'h1;
  assign v_13977 = v_13978 & v_13979;
  assign v_13978 = ~act_13790;
  assign v_13979 = v_13980 | v_13988;
  assign v_13980 = v_13981 | v_13986;
  assign v_13981 = mux_13981(v_13982);
  assign v_13982 = v_13787 & v_13983;
  assign v_13983 = v_13984 & 1'h1;
  assign v_13984 = v_13985 | 1'h0;
  assign v_13985 = ~v_13780;
  assign v_13986 = mux_13986(v_13987);
  assign v_13987 = ~v_13982;
  assign v_13988 = ~v_13787;
  assign v_13989 = v_13990 | v_13991;
  assign v_13990 = mux_13990(v_13789);
  assign v_13991 = mux_13991(v_13976);
  assign v_13993 = v_13994 | v_14181;
  assign v_13994 = act_13995 & 1'h1;
  assign act_13995 = v_13996 | v_14082;
  assign v_13996 = v_13997 & v_14083;
  assign v_13997 = v_13998 & v_14092;
  assign v_13998 = ~v_13999;
  assign v_14000 = v_14001 | v_14076;
  assign v_14001 = act_14002 & 1'h1;
  assign act_14002 = v_14003 | v_14033;
  assign v_14003 = v_14004 & v_14034;
  assign v_14004 = v_14005 & v_14043;
  assign v_14005 = ~v_14006;
  assign v_14007 = v_14008 | v_14027;
  assign v_14008 = act_14009 & 1'h1;
  assign act_14009 = v_14010 | v_14016;
  assign v_14010 = v_14011 & v_14017;
  assign v_14011 = v_14012 & vout_canPeek_14022;
  assign v_14012 = ~vout_canPeek_14013;
  pebbles_core
    pebbles_core_14013
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14014),
       .in0_consume_en(vin0_consume_en_14013),
       .out_canPeek(vout_canPeek_14013),
       .out_peek(vout_peek_14013));
  assign v_14014 = v_14015 | v_14020;
  assign v_14015 = mux_14015(v_14016);
  assign v_14016 = vout_canPeek_14013 & v_14017;
  assign v_14017 = v_14018 & 1'h1;
  assign v_14018 = v_14019 | 1'h0;
  assign v_14019 = ~v_14006;
  assign v_14020 = mux_14020(v_14021);
  assign v_14021 = ~v_14016;
  pebbles_core
    pebbles_core_14022
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14023),
       .in0_consume_en(vin0_consume_en_14022),
       .out_canPeek(vout_canPeek_14022),
       .out_peek(vout_peek_14022));
  assign v_14023 = v_14024 | v_14025;
  assign v_14024 = mux_14024(v_14010);
  assign v_14025 = mux_14025(v_14026);
  assign v_14026 = ~v_14010;
  assign v_14027 = v_14028 & 1'h1;
  assign v_14028 = v_14029 & v_14030;
  assign v_14029 = ~act_14009;
  assign v_14030 = v_14031 | v_14039;
  assign v_14031 = v_14032 | v_14037;
  assign v_14032 = mux_14032(v_14033);
  assign v_14033 = v_14006 & v_14034;
  assign v_14034 = v_14035 & 1'h1;
  assign v_14035 = v_14036 | 1'h0;
  assign v_14036 = ~v_13999;
  assign v_14037 = mux_14037(v_14038);
  assign v_14038 = ~v_14033;
  assign v_14039 = ~v_14006;
  assign v_14040 = v_14041 | v_14042;
  assign v_14041 = mux_14041(v_14008);
  assign v_14042 = mux_14042(v_14027);
  assign v_14044 = v_14045 | v_14064;
  assign v_14045 = act_14046 & 1'h1;
  assign act_14046 = v_14047 | v_14053;
  assign v_14047 = v_14048 & v_14054;
  assign v_14048 = v_14049 & vout_canPeek_14059;
  assign v_14049 = ~vout_canPeek_14050;
  pebbles_core
    pebbles_core_14050
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14051),
       .in0_consume_en(vin0_consume_en_14050),
       .out_canPeek(vout_canPeek_14050),
       .out_peek(vout_peek_14050));
  assign v_14051 = v_14052 | v_14057;
  assign v_14052 = mux_14052(v_14053);
  assign v_14053 = vout_canPeek_14050 & v_14054;
  assign v_14054 = v_14055 & 1'h1;
  assign v_14055 = v_14056 | 1'h0;
  assign v_14056 = ~v_14043;
  assign v_14057 = mux_14057(v_14058);
  assign v_14058 = ~v_14053;
  pebbles_core
    pebbles_core_14059
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14060),
       .in0_consume_en(vin0_consume_en_14059),
       .out_canPeek(vout_canPeek_14059),
       .out_peek(vout_peek_14059));
  assign v_14060 = v_14061 | v_14062;
  assign v_14061 = mux_14061(v_14047);
  assign v_14062 = mux_14062(v_14063);
  assign v_14063 = ~v_14047;
  assign v_14064 = v_14065 & 1'h1;
  assign v_14065 = v_14066 & v_14067;
  assign v_14066 = ~act_14046;
  assign v_14067 = v_14068 | v_14072;
  assign v_14068 = v_14069 | v_14070;
  assign v_14069 = mux_14069(v_14003);
  assign v_14070 = mux_14070(v_14071);
  assign v_14071 = ~v_14003;
  assign v_14072 = ~v_14043;
  assign v_14073 = v_14074 | v_14075;
  assign v_14074 = mux_14074(v_14045);
  assign v_14075 = mux_14075(v_14064);
  assign v_14076 = v_14077 & 1'h1;
  assign v_14077 = v_14078 & v_14079;
  assign v_14078 = ~act_14002;
  assign v_14079 = v_14080 | v_14088;
  assign v_14080 = v_14081 | v_14086;
  assign v_14081 = mux_14081(v_14082);
  assign v_14082 = v_13999 & v_14083;
  assign v_14083 = v_14084 & 1'h1;
  assign v_14084 = v_14085 | 1'h0;
  assign v_14085 = ~v_13992;
  assign v_14086 = mux_14086(v_14087);
  assign v_14087 = ~v_14082;
  assign v_14088 = ~v_13999;
  assign v_14089 = v_14090 | v_14091;
  assign v_14090 = mux_14090(v_14001);
  assign v_14091 = mux_14091(v_14076);
  assign v_14093 = v_14094 | v_14169;
  assign v_14094 = act_14095 & 1'h1;
  assign act_14095 = v_14096 | v_14126;
  assign v_14096 = v_14097 & v_14127;
  assign v_14097 = v_14098 & v_14136;
  assign v_14098 = ~v_14099;
  assign v_14100 = v_14101 | v_14120;
  assign v_14101 = act_14102 & 1'h1;
  assign act_14102 = v_14103 | v_14109;
  assign v_14103 = v_14104 & v_14110;
  assign v_14104 = v_14105 & vout_canPeek_14115;
  assign v_14105 = ~vout_canPeek_14106;
  pebbles_core
    pebbles_core_14106
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14107),
       .in0_consume_en(vin0_consume_en_14106),
       .out_canPeek(vout_canPeek_14106),
       .out_peek(vout_peek_14106));
  assign v_14107 = v_14108 | v_14113;
  assign v_14108 = mux_14108(v_14109);
  assign v_14109 = vout_canPeek_14106 & v_14110;
  assign v_14110 = v_14111 & 1'h1;
  assign v_14111 = v_14112 | 1'h0;
  assign v_14112 = ~v_14099;
  assign v_14113 = mux_14113(v_14114);
  assign v_14114 = ~v_14109;
  pebbles_core
    pebbles_core_14115
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14116),
       .in0_consume_en(vin0_consume_en_14115),
       .out_canPeek(vout_canPeek_14115),
       .out_peek(vout_peek_14115));
  assign v_14116 = v_14117 | v_14118;
  assign v_14117 = mux_14117(v_14103);
  assign v_14118 = mux_14118(v_14119);
  assign v_14119 = ~v_14103;
  assign v_14120 = v_14121 & 1'h1;
  assign v_14121 = v_14122 & v_14123;
  assign v_14122 = ~act_14102;
  assign v_14123 = v_14124 | v_14132;
  assign v_14124 = v_14125 | v_14130;
  assign v_14125 = mux_14125(v_14126);
  assign v_14126 = v_14099 & v_14127;
  assign v_14127 = v_14128 & 1'h1;
  assign v_14128 = v_14129 | 1'h0;
  assign v_14129 = ~v_14092;
  assign v_14130 = mux_14130(v_14131);
  assign v_14131 = ~v_14126;
  assign v_14132 = ~v_14099;
  assign v_14133 = v_14134 | v_14135;
  assign v_14134 = mux_14134(v_14101);
  assign v_14135 = mux_14135(v_14120);
  assign v_14137 = v_14138 | v_14157;
  assign v_14138 = act_14139 & 1'h1;
  assign act_14139 = v_14140 | v_14146;
  assign v_14140 = v_14141 & v_14147;
  assign v_14141 = v_14142 & vout_canPeek_14152;
  assign v_14142 = ~vout_canPeek_14143;
  pebbles_core
    pebbles_core_14143
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14144),
       .in0_consume_en(vin0_consume_en_14143),
       .out_canPeek(vout_canPeek_14143),
       .out_peek(vout_peek_14143));
  assign v_14144 = v_14145 | v_14150;
  assign v_14145 = mux_14145(v_14146);
  assign v_14146 = vout_canPeek_14143 & v_14147;
  assign v_14147 = v_14148 & 1'h1;
  assign v_14148 = v_14149 | 1'h0;
  assign v_14149 = ~v_14136;
  assign v_14150 = mux_14150(v_14151);
  assign v_14151 = ~v_14146;
  pebbles_core
    pebbles_core_14152
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14153),
       .in0_consume_en(vin0_consume_en_14152),
       .out_canPeek(vout_canPeek_14152),
       .out_peek(vout_peek_14152));
  assign v_14153 = v_14154 | v_14155;
  assign v_14154 = mux_14154(v_14140);
  assign v_14155 = mux_14155(v_14156);
  assign v_14156 = ~v_14140;
  assign v_14157 = v_14158 & 1'h1;
  assign v_14158 = v_14159 & v_14160;
  assign v_14159 = ~act_14139;
  assign v_14160 = v_14161 | v_14165;
  assign v_14161 = v_14162 | v_14163;
  assign v_14162 = mux_14162(v_14096);
  assign v_14163 = mux_14163(v_14164);
  assign v_14164 = ~v_14096;
  assign v_14165 = ~v_14136;
  assign v_14166 = v_14167 | v_14168;
  assign v_14167 = mux_14167(v_14138);
  assign v_14168 = mux_14168(v_14157);
  assign v_14169 = v_14170 & 1'h1;
  assign v_14170 = v_14171 & v_14172;
  assign v_14171 = ~act_14095;
  assign v_14172 = v_14173 | v_14177;
  assign v_14173 = v_14174 | v_14175;
  assign v_14174 = mux_14174(v_13996);
  assign v_14175 = mux_14175(v_14176);
  assign v_14176 = ~v_13996;
  assign v_14177 = ~v_14092;
  assign v_14178 = v_14179 | v_14180;
  assign v_14179 = mux_14179(v_14094);
  assign v_14180 = mux_14180(v_14169);
  assign v_14181 = v_14182 & 1'h1;
  assign v_14182 = v_14183 & v_14184;
  assign v_14183 = ~act_13995;
  assign v_14184 = v_14185 | v_14189;
  assign v_14185 = v_14186 | v_14187;
  assign v_14186 = mux_14186(v_13784);
  assign v_14187 = mux_14187(v_14188);
  assign v_14188 = ~v_13784;
  assign v_14189 = ~v_13992;
  assign v_14190 = v_14191 | v_14192;
  assign v_14191 = mux_14191(v_13994);
  assign v_14192 = mux_14192(v_14181);
  assign v_14193 = v_14194 & 1'h1;
  assign v_14194 = v_14195 & v_14196;
  assign v_14195 = ~act_13783;
  assign v_14196 = v_14197 | v_14201;
  assign v_14197 = v_14198 | v_14199;
  assign v_14198 = mux_14198(v_13348);
  assign v_14199 = mux_14199(v_14200);
  assign v_14200 = ~v_13348;
  assign v_14201 = ~v_13780;
  assign v_14202 = v_14203 | v_14204;
  assign v_14203 = mux_14203(v_13782);
  assign v_14204 = mux_14204(v_14193);
  assign v_14205 = v_14206 & 1'h1;
  assign v_14206 = v_14207 & v_14208;
  assign v_14207 = ~act_13347;
  assign v_14208 = v_14209 | v_14217;
  assign v_14209 = v_14210 | v_14215;
  assign v_14210 = mux_14210(v_14211);
  assign v_14211 = v_13344 & v_14212;
  assign v_14212 = v_14213 & 1'h1;
  assign v_14213 = v_14214 | 1'h0;
  assign v_14214 = ~v_13337;
  assign v_14215 = mux_14215(v_14216);
  assign v_14216 = ~v_14211;
  assign v_14217 = ~v_13344;
  assign v_14218 = v_14219 | v_14220;
  assign v_14219 = mux_14219(v_13346);
  assign v_14220 = mux_14220(v_14205);
  assign v_14222 = v_14223 | v_15082;
  assign v_14223 = act_14224 & 1'h1;
  assign act_14224 = v_14225 | v_14647;
  assign v_14225 = v_14226 & v_14648;
  assign v_14226 = v_14227 & v_14657;
  assign v_14227 = ~v_14228;
  assign v_14229 = v_14230 | v_14641;
  assign v_14230 = act_14231 & 1'h1;
  assign act_14231 = v_14232 | v_14430;
  assign v_14232 = v_14233 & v_14431;
  assign v_14233 = v_14234 & v_14440;
  assign v_14234 = ~v_14235;
  assign v_14236 = v_14237 | v_14424;
  assign v_14237 = act_14238 & 1'h1;
  assign act_14238 = v_14239 | v_14325;
  assign v_14239 = v_14240 & v_14326;
  assign v_14240 = v_14241 & v_14335;
  assign v_14241 = ~v_14242;
  assign v_14243 = v_14244 | v_14319;
  assign v_14244 = act_14245 & 1'h1;
  assign act_14245 = v_14246 | v_14276;
  assign v_14246 = v_14247 & v_14277;
  assign v_14247 = v_14248 & v_14286;
  assign v_14248 = ~v_14249;
  assign v_14250 = v_14251 | v_14270;
  assign v_14251 = act_14252 & 1'h1;
  assign act_14252 = v_14253 | v_14259;
  assign v_14253 = v_14254 & v_14260;
  assign v_14254 = v_14255 & vout_canPeek_14265;
  assign v_14255 = ~vout_canPeek_14256;
  pebbles_core
    pebbles_core_14256
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14257),
       .in0_consume_en(vin0_consume_en_14256),
       .out_canPeek(vout_canPeek_14256),
       .out_peek(vout_peek_14256));
  assign v_14257 = v_14258 | v_14263;
  assign v_14258 = mux_14258(v_14259);
  assign v_14259 = vout_canPeek_14256 & v_14260;
  assign v_14260 = v_14261 & 1'h1;
  assign v_14261 = v_14262 | 1'h0;
  assign v_14262 = ~v_14249;
  assign v_14263 = mux_14263(v_14264);
  assign v_14264 = ~v_14259;
  pebbles_core
    pebbles_core_14265
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14266),
       .in0_consume_en(vin0_consume_en_14265),
       .out_canPeek(vout_canPeek_14265),
       .out_peek(vout_peek_14265));
  assign v_14266 = v_14267 | v_14268;
  assign v_14267 = mux_14267(v_14253);
  assign v_14268 = mux_14268(v_14269);
  assign v_14269 = ~v_14253;
  assign v_14270 = v_14271 & 1'h1;
  assign v_14271 = v_14272 & v_14273;
  assign v_14272 = ~act_14252;
  assign v_14273 = v_14274 | v_14282;
  assign v_14274 = v_14275 | v_14280;
  assign v_14275 = mux_14275(v_14276);
  assign v_14276 = v_14249 & v_14277;
  assign v_14277 = v_14278 & 1'h1;
  assign v_14278 = v_14279 | 1'h0;
  assign v_14279 = ~v_14242;
  assign v_14280 = mux_14280(v_14281);
  assign v_14281 = ~v_14276;
  assign v_14282 = ~v_14249;
  assign v_14283 = v_14284 | v_14285;
  assign v_14284 = mux_14284(v_14251);
  assign v_14285 = mux_14285(v_14270);
  assign v_14287 = v_14288 | v_14307;
  assign v_14288 = act_14289 & 1'h1;
  assign act_14289 = v_14290 | v_14296;
  assign v_14290 = v_14291 & v_14297;
  assign v_14291 = v_14292 & vout_canPeek_14302;
  assign v_14292 = ~vout_canPeek_14293;
  pebbles_core
    pebbles_core_14293
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14294),
       .in0_consume_en(vin0_consume_en_14293),
       .out_canPeek(vout_canPeek_14293),
       .out_peek(vout_peek_14293));
  assign v_14294 = v_14295 | v_14300;
  assign v_14295 = mux_14295(v_14296);
  assign v_14296 = vout_canPeek_14293 & v_14297;
  assign v_14297 = v_14298 & 1'h1;
  assign v_14298 = v_14299 | 1'h0;
  assign v_14299 = ~v_14286;
  assign v_14300 = mux_14300(v_14301);
  assign v_14301 = ~v_14296;
  pebbles_core
    pebbles_core_14302
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14303),
       .in0_consume_en(vin0_consume_en_14302),
       .out_canPeek(vout_canPeek_14302),
       .out_peek(vout_peek_14302));
  assign v_14303 = v_14304 | v_14305;
  assign v_14304 = mux_14304(v_14290);
  assign v_14305 = mux_14305(v_14306);
  assign v_14306 = ~v_14290;
  assign v_14307 = v_14308 & 1'h1;
  assign v_14308 = v_14309 & v_14310;
  assign v_14309 = ~act_14289;
  assign v_14310 = v_14311 | v_14315;
  assign v_14311 = v_14312 | v_14313;
  assign v_14312 = mux_14312(v_14246);
  assign v_14313 = mux_14313(v_14314);
  assign v_14314 = ~v_14246;
  assign v_14315 = ~v_14286;
  assign v_14316 = v_14317 | v_14318;
  assign v_14317 = mux_14317(v_14288);
  assign v_14318 = mux_14318(v_14307);
  assign v_14319 = v_14320 & 1'h1;
  assign v_14320 = v_14321 & v_14322;
  assign v_14321 = ~act_14245;
  assign v_14322 = v_14323 | v_14331;
  assign v_14323 = v_14324 | v_14329;
  assign v_14324 = mux_14324(v_14325);
  assign v_14325 = v_14242 & v_14326;
  assign v_14326 = v_14327 & 1'h1;
  assign v_14327 = v_14328 | 1'h0;
  assign v_14328 = ~v_14235;
  assign v_14329 = mux_14329(v_14330);
  assign v_14330 = ~v_14325;
  assign v_14331 = ~v_14242;
  assign v_14332 = v_14333 | v_14334;
  assign v_14333 = mux_14333(v_14244);
  assign v_14334 = mux_14334(v_14319);
  assign v_14336 = v_14337 | v_14412;
  assign v_14337 = act_14338 & 1'h1;
  assign act_14338 = v_14339 | v_14369;
  assign v_14339 = v_14340 & v_14370;
  assign v_14340 = v_14341 & v_14379;
  assign v_14341 = ~v_14342;
  assign v_14343 = v_14344 | v_14363;
  assign v_14344 = act_14345 & 1'h1;
  assign act_14345 = v_14346 | v_14352;
  assign v_14346 = v_14347 & v_14353;
  assign v_14347 = v_14348 & vout_canPeek_14358;
  assign v_14348 = ~vout_canPeek_14349;
  pebbles_core
    pebbles_core_14349
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14350),
       .in0_consume_en(vin0_consume_en_14349),
       .out_canPeek(vout_canPeek_14349),
       .out_peek(vout_peek_14349));
  assign v_14350 = v_14351 | v_14356;
  assign v_14351 = mux_14351(v_14352);
  assign v_14352 = vout_canPeek_14349 & v_14353;
  assign v_14353 = v_14354 & 1'h1;
  assign v_14354 = v_14355 | 1'h0;
  assign v_14355 = ~v_14342;
  assign v_14356 = mux_14356(v_14357);
  assign v_14357 = ~v_14352;
  pebbles_core
    pebbles_core_14358
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14359),
       .in0_consume_en(vin0_consume_en_14358),
       .out_canPeek(vout_canPeek_14358),
       .out_peek(vout_peek_14358));
  assign v_14359 = v_14360 | v_14361;
  assign v_14360 = mux_14360(v_14346);
  assign v_14361 = mux_14361(v_14362);
  assign v_14362 = ~v_14346;
  assign v_14363 = v_14364 & 1'h1;
  assign v_14364 = v_14365 & v_14366;
  assign v_14365 = ~act_14345;
  assign v_14366 = v_14367 | v_14375;
  assign v_14367 = v_14368 | v_14373;
  assign v_14368 = mux_14368(v_14369);
  assign v_14369 = v_14342 & v_14370;
  assign v_14370 = v_14371 & 1'h1;
  assign v_14371 = v_14372 | 1'h0;
  assign v_14372 = ~v_14335;
  assign v_14373 = mux_14373(v_14374);
  assign v_14374 = ~v_14369;
  assign v_14375 = ~v_14342;
  assign v_14376 = v_14377 | v_14378;
  assign v_14377 = mux_14377(v_14344);
  assign v_14378 = mux_14378(v_14363);
  assign v_14380 = v_14381 | v_14400;
  assign v_14381 = act_14382 & 1'h1;
  assign act_14382 = v_14383 | v_14389;
  assign v_14383 = v_14384 & v_14390;
  assign v_14384 = v_14385 & vout_canPeek_14395;
  assign v_14385 = ~vout_canPeek_14386;
  pebbles_core
    pebbles_core_14386
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14387),
       .in0_consume_en(vin0_consume_en_14386),
       .out_canPeek(vout_canPeek_14386),
       .out_peek(vout_peek_14386));
  assign v_14387 = v_14388 | v_14393;
  assign v_14388 = mux_14388(v_14389);
  assign v_14389 = vout_canPeek_14386 & v_14390;
  assign v_14390 = v_14391 & 1'h1;
  assign v_14391 = v_14392 | 1'h0;
  assign v_14392 = ~v_14379;
  assign v_14393 = mux_14393(v_14394);
  assign v_14394 = ~v_14389;
  pebbles_core
    pebbles_core_14395
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14396),
       .in0_consume_en(vin0_consume_en_14395),
       .out_canPeek(vout_canPeek_14395),
       .out_peek(vout_peek_14395));
  assign v_14396 = v_14397 | v_14398;
  assign v_14397 = mux_14397(v_14383);
  assign v_14398 = mux_14398(v_14399);
  assign v_14399 = ~v_14383;
  assign v_14400 = v_14401 & 1'h1;
  assign v_14401 = v_14402 & v_14403;
  assign v_14402 = ~act_14382;
  assign v_14403 = v_14404 | v_14408;
  assign v_14404 = v_14405 | v_14406;
  assign v_14405 = mux_14405(v_14339);
  assign v_14406 = mux_14406(v_14407);
  assign v_14407 = ~v_14339;
  assign v_14408 = ~v_14379;
  assign v_14409 = v_14410 | v_14411;
  assign v_14410 = mux_14410(v_14381);
  assign v_14411 = mux_14411(v_14400);
  assign v_14412 = v_14413 & 1'h1;
  assign v_14413 = v_14414 & v_14415;
  assign v_14414 = ~act_14338;
  assign v_14415 = v_14416 | v_14420;
  assign v_14416 = v_14417 | v_14418;
  assign v_14417 = mux_14417(v_14239);
  assign v_14418 = mux_14418(v_14419);
  assign v_14419 = ~v_14239;
  assign v_14420 = ~v_14335;
  assign v_14421 = v_14422 | v_14423;
  assign v_14422 = mux_14422(v_14337);
  assign v_14423 = mux_14423(v_14412);
  assign v_14424 = v_14425 & 1'h1;
  assign v_14425 = v_14426 & v_14427;
  assign v_14426 = ~act_14238;
  assign v_14427 = v_14428 | v_14436;
  assign v_14428 = v_14429 | v_14434;
  assign v_14429 = mux_14429(v_14430);
  assign v_14430 = v_14235 & v_14431;
  assign v_14431 = v_14432 & 1'h1;
  assign v_14432 = v_14433 | 1'h0;
  assign v_14433 = ~v_14228;
  assign v_14434 = mux_14434(v_14435);
  assign v_14435 = ~v_14430;
  assign v_14436 = ~v_14235;
  assign v_14437 = v_14438 | v_14439;
  assign v_14438 = mux_14438(v_14237);
  assign v_14439 = mux_14439(v_14424);
  assign v_14441 = v_14442 | v_14629;
  assign v_14442 = act_14443 & 1'h1;
  assign act_14443 = v_14444 | v_14530;
  assign v_14444 = v_14445 & v_14531;
  assign v_14445 = v_14446 & v_14540;
  assign v_14446 = ~v_14447;
  assign v_14448 = v_14449 | v_14524;
  assign v_14449 = act_14450 & 1'h1;
  assign act_14450 = v_14451 | v_14481;
  assign v_14451 = v_14452 & v_14482;
  assign v_14452 = v_14453 & v_14491;
  assign v_14453 = ~v_14454;
  assign v_14455 = v_14456 | v_14475;
  assign v_14456 = act_14457 & 1'h1;
  assign act_14457 = v_14458 | v_14464;
  assign v_14458 = v_14459 & v_14465;
  assign v_14459 = v_14460 & vout_canPeek_14470;
  assign v_14460 = ~vout_canPeek_14461;
  pebbles_core
    pebbles_core_14461
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14462),
       .in0_consume_en(vin0_consume_en_14461),
       .out_canPeek(vout_canPeek_14461),
       .out_peek(vout_peek_14461));
  assign v_14462 = v_14463 | v_14468;
  assign v_14463 = mux_14463(v_14464);
  assign v_14464 = vout_canPeek_14461 & v_14465;
  assign v_14465 = v_14466 & 1'h1;
  assign v_14466 = v_14467 | 1'h0;
  assign v_14467 = ~v_14454;
  assign v_14468 = mux_14468(v_14469);
  assign v_14469 = ~v_14464;
  pebbles_core
    pebbles_core_14470
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14471),
       .in0_consume_en(vin0_consume_en_14470),
       .out_canPeek(vout_canPeek_14470),
       .out_peek(vout_peek_14470));
  assign v_14471 = v_14472 | v_14473;
  assign v_14472 = mux_14472(v_14458);
  assign v_14473 = mux_14473(v_14474);
  assign v_14474 = ~v_14458;
  assign v_14475 = v_14476 & 1'h1;
  assign v_14476 = v_14477 & v_14478;
  assign v_14477 = ~act_14457;
  assign v_14478 = v_14479 | v_14487;
  assign v_14479 = v_14480 | v_14485;
  assign v_14480 = mux_14480(v_14481);
  assign v_14481 = v_14454 & v_14482;
  assign v_14482 = v_14483 & 1'h1;
  assign v_14483 = v_14484 | 1'h0;
  assign v_14484 = ~v_14447;
  assign v_14485 = mux_14485(v_14486);
  assign v_14486 = ~v_14481;
  assign v_14487 = ~v_14454;
  assign v_14488 = v_14489 | v_14490;
  assign v_14489 = mux_14489(v_14456);
  assign v_14490 = mux_14490(v_14475);
  assign v_14492 = v_14493 | v_14512;
  assign v_14493 = act_14494 & 1'h1;
  assign act_14494 = v_14495 | v_14501;
  assign v_14495 = v_14496 & v_14502;
  assign v_14496 = v_14497 & vout_canPeek_14507;
  assign v_14497 = ~vout_canPeek_14498;
  pebbles_core
    pebbles_core_14498
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14499),
       .in0_consume_en(vin0_consume_en_14498),
       .out_canPeek(vout_canPeek_14498),
       .out_peek(vout_peek_14498));
  assign v_14499 = v_14500 | v_14505;
  assign v_14500 = mux_14500(v_14501);
  assign v_14501 = vout_canPeek_14498 & v_14502;
  assign v_14502 = v_14503 & 1'h1;
  assign v_14503 = v_14504 | 1'h0;
  assign v_14504 = ~v_14491;
  assign v_14505 = mux_14505(v_14506);
  assign v_14506 = ~v_14501;
  pebbles_core
    pebbles_core_14507
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14508),
       .in0_consume_en(vin0_consume_en_14507),
       .out_canPeek(vout_canPeek_14507),
       .out_peek(vout_peek_14507));
  assign v_14508 = v_14509 | v_14510;
  assign v_14509 = mux_14509(v_14495);
  assign v_14510 = mux_14510(v_14511);
  assign v_14511 = ~v_14495;
  assign v_14512 = v_14513 & 1'h1;
  assign v_14513 = v_14514 & v_14515;
  assign v_14514 = ~act_14494;
  assign v_14515 = v_14516 | v_14520;
  assign v_14516 = v_14517 | v_14518;
  assign v_14517 = mux_14517(v_14451);
  assign v_14518 = mux_14518(v_14519);
  assign v_14519 = ~v_14451;
  assign v_14520 = ~v_14491;
  assign v_14521 = v_14522 | v_14523;
  assign v_14522 = mux_14522(v_14493);
  assign v_14523 = mux_14523(v_14512);
  assign v_14524 = v_14525 & 1'h1;
  assign v_14525 = v_14526 & v_14527;
  assign v_14526 = ~act_14450;
  assign v_14527 = v_14528 | v_14536;
  assign v_14528 = v_14529 | v_14534;
  assign v_14529 = mux_14529(v_14530);
  assign v_14530 = v_14447 & v_14531;
  assign v_14531 = v_14532 & 1'h1;
  assign v_14532 = v_14533 | 1'h0;
  assign v_14533 = ~v_14440;
  assign v_14534 = mux_14534(v_14535);
  assign v_14535 = ~v_14530;
  assign v_14536 = ~v_14447;
  assign v_14537 = v_14538 | v_14539;
  assign v_14538 = mux_14538(v_14449);
  assign v_14539 = mux_14539(v_14524);
  assign v_14541 = v_14542 | v_14617;
  assign v_14542 = act_14543 & 1'h1;
  assign act_14543 = v_14544 | v_14574;
  assign v_14544 = v_14545 & v_14575;
  assign v_14545 = v_14546 & v_14584;
  assign v_14546 = ~v_14547;
  assign v_14548 = v_14549 | v_14568;
  assign v_14549 = act_14550 & 1'h1;
  assign act_14550 = v_14551 | v_14557;
  assign v_14551 = v_14552 & v_14558;
  assign v_14552 = v_14553 & vout_canPeek_14563;
  assign v_14553 = ~vout_canPeek_14554;
  pebbles_core
    pebbles_core_14554
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14555),
       .in0_consume_en(vin0_consume_en_14554),
       .out_canPeek(vout_canPeek_14554),
       .out_peek(vout_peek_14554));
  assign v_14555 = v_14556 | v_14561;
  assign v_14556 = mux_14556(v_14557);
  assign v_14557 = vout_canPeek_14554 & v_14558;
  assign v_14558 = v_14559 & 1'h1;
  assign v_14559 = v_14560 | 1'h0;
  assign v_14560 = ~v_14547;
  assign v_14561 = mux_14561(v_14562);
  assign v_14562 = ~v_14557;
  pebbles_core
    pebbles_core_14563
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14564),
       .in0_consume_en(vin0_consume_en_14563),
       .out_canPeek(vout_canPeek_14563),
       .out_peek(vout_peek_14563));
  assign v_14564 = v_14565 | v_14566;
  assign v_14565 = mux_14565(v_14551);
  assign v_14566 = mux_14566(v_14567);
  assign v_14567 = ~v_14551;
  assign v_14568 = v_14569 & 1'h1;
  assign v_14569 = v_14570 & v_14571;
  assign v_14570 = ~act_14550;
  assign v_14571 = v_14572 | v_14580;
  assign v_14572 = v_14573 | v_14578;
  assign v_14573 = mux_14573(v_14574);
  assign v_14574 = v_14547 & v_14575;
  assign v_14575 = v_14576 & 1'h1;
  assign v_14576 = v_14577 | 1'h0;
  assign v_14577 = ~v_14540;
  assign v_14578 = mux_14578(v_14579);
  assign v_14579 = ~v_14574;
  assign v_14580 = ~v_14547;
  assign v_14581 = v_14582 | v_14583;
  assign v_14582 = mux_14582(v_14549);
  assign v_14583 = mux_14583(v_14568);
  assign v_14585 = v_14586 | v_14605;
  assign v_14586 = act_14587 & 1'h1;
  assign act_14587 = v_14588 | v_14594;
  assign v_14588 = v_14589 & v_14595;
  assign v_14589 = v_14590 & vout_canPeek_14600;
  assign v_14590 = ~vout_canPeek_14591;
  pebbles_core
    pebbles_core_14591
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14592),
       .in0_consume_en(vin0_consume_en_14591),
       .out_canPeek(vout_canPeek_14591),
       .out_peek(vout_peek_14591));
  assign v_14592 = v_14593 | v_14598;
  assign v_14593 = mux_14593(v_14594);
  assign v_14594 = vout_canPeek_14591 & v_14595;
  assign v_14595 = v_14596 & 1'h1;
  assign v_14596 = v_14597 | 1'h0;
  assign v_14597 = ~v_14584;
  assign v_14598 = mux_14598(v_14599);
  assign v_14599 = ~v_14594;
  pebbles_core
    pebbles_core_14600
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14601),
       .in0_consume_en(vin0_consume_en_14600),
       .out_canPeek(vout_canPeek_14600),
       .out_peek(vout_peek_14600));
  assign v_14601 = v_14602 | v_14603;
  assign v_14602 = mux_14602(v_14588);
  assign v_14603 = mux_14603(v_14604);
  assign v_14604 = ~v_14588;
  assign v_14605 = v_14606 & 1'h1;
  assign v_14606 = v_14607 & v_14608;
  assign v_14607 = ~act_14587;
  assign v_14608 = v_14609 | v_14613;
  assign v_14609 = v_14610 | v_14611;
  assign v_14610 = mux_14610(v_14544);
  assign v_14611 = mux_14611(v_14612);
  assign v_14612 = ~v_14544;
  assign v_14613 = ~v_14584;
  assign v_14614 = v_14615 | v_14616;
  assign v_14615 = mux_14615(v_14586);
  assign v_14616 = mux_14616(v_14605);
  assign v_14617 = v_14618 & 1'h1;
  assign v_14618 = v_14619 & v_14620;
  assign v_14619 = ~act_14543;
  assign v_14620 = v_14621 | v_14625;
  assign v_14621 = v_14622 | v_14623;
  assign v_14622 = mux_14622(v_14444);
  assign v_14623 = mux_14623(v_14624);
  assign v_14624 = ~v_14444;
  assign v_14625 = ~v_14540;
  assign v_14626 = v_14627 | v_14628;
  assign v_14627 = mux_14627(v_14542);
  assign v_14628 = mux_14628(v_14617);
  assign v_14629 = v_14630 & 1'h1;
  assign v_14630 = v_14631 & v_14632;
  assign v_14631 = ~act_14443;
  assign v_14632 = v_14633 | v_14637;
  assign v_14633 = v_14634 | v_14635;
  assign v_14634 = mux_14634(v_14232);
  assign v_14635 = mux_14635(v_14636);
  assign v_14636 = ~v_14232;
  assign v_14637 = ~v_14440;
  assign v_14638 = v_14639 | v_14640;
  assign v_14639 = mux_14639(v_14442);
  assign v_14640 = mux_14640(v_14629);
  assign v_14641 = v_14642 & 1'h1;
  assign v_14642 = v_14643 & v_14644;
  assign v_14643 = ~act_14231;
  assign v_14644 = v_14645 | v_14653;
  assign v_14645 = v_14646 | v_14651;
  assign v_14646 = mux_14646(v_14647);
  assign v_14647 = v_14228 & v_14648;
  assign v_14648 = v_14649 & 1'h1;
  assign v_14649 = v_14650 | 1'h0;
  assign v_14650 = ~v_14221;
  assign v_14651 = mux_14651(v_14652);
  assign v_14652 = ~v_14647;
  assign v_14653 = ~v_14228;
  assign v_14654 = v_14655 | v_14656;
  assign v_14655 = mux_14655(v_14230);
  assign v_14656 = mux_14656(v_14641);
  assign v_14658 = v_14659 | v_15070;
  assign v_14659 = act_14660 & 1'h1;
  assign act_14660 = v_14661 | v_14859;
  assign v_14661 = v_14662 & v_14860;
  assign v_14662 = v_14663 & v_14869;
  assign v_14663 = ~v_14664;
  assign v_14665 = v_14666 | v_14853;
  assign v_14666 = act_14667 & 1'h1;
  assign act_14667 = v_14668 | v_14754;
  assign v_14668 = v_14669 & v_14755;
  assign v_14669 = v_14670 & v_14764;
  assign v_14670 = ~v_14671;
  assign v_14672 = v_14673 | v_14748;
  assign v_14673 = act_14674 & 1'h1;
  assign act_14674 = v_14675 | v_14705;
  assign v_14675 = v_14676 & v_14706;
  assign v_14676 = v_14677 & v_14715;
  assign v_14677 = ~v_14678;
  assign v_14679 = v_14680 | v_14699;
  assign v_14680 = act_14681 & 1'h1;
  assign act_14681 = v_14682 | v_14688;
  assign v_14682 = v_14683 & v_14689;
  assign v_14683 = v_14684 & vout_canPeek_14694;
  assign v_14684 = ~vout_canPeek_14685;
  pebbles_core
    pebbles_core_14685
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14686),
       .in0_consume_en(vin0_consume_en_14685),
       .out_canPeek(vout_canPeek_14685),
       .out_peek(vout_peek_14685));
  assign v_14686 = v_14687 | v_14692;
  assign v_14687 = mux_14687(v_14688);
  assign v_14688 = vout_canPeek_14685 & v_14689;
  assign v_14689 = v_14690 & 1'h1;
  assign v_14690 = v_14691 | 1'h0;
  assign v_14691 = ~v_14678;
  assign v_14692 = mux_14692(v_14693);
  assign v_14693 = ~v_14688;
  pebbles_core
    pebbles_core_14694
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14695),
       .in0_consume_en(vin0_consume_en_14694),
       .out_canPeek(vout_canPeek_14694),
       .out_peek(vout_peek_14694));
  assign v_14695 = v_14696 | v_14697;
  assign v_14696 = mux_14696(v_14682);
  assign v_14697 = mux_14697(v_14698);
  assign v_14698 = ~v_14682;
  assign v_14699 = v_14700 & 1'h1;
  assign v_14700 = v_14701 & v_14702;
  assign v_14701 = ~act_14681;
  assign v_14702 = v_14703 | v_14711;
  assign v_14703 = v_14704 | v_14709;
  assign v_14704 = mux_14704(v_14705);
  assign v_14705 = v_14678 & v_14706;
  assign v_14706 = v_14707 & 1'h1;
  assign v_14707 = v_14708 | 1'h0;
  assign v_14708 = ~v_14671;
  assign v_14709 = mux_14709(v_14710);
  assign v_14710 = ~v_14705;
  assign v_14711 = ~v_14678;
  assign v_14712 = v_14713 | v_14714;
  assign v_14713 = mux_14713(v_14680);
  assign v_14714 = mux_14714(v_14699);
  assign v_14716 = v_14717 | v_14736;
  assign v_14717 = act_14718 & 1'h1;
  assign act_14718 = v_14719 | v_14725;
  assign v_14719 = v_14720 & v_14726;
  assign v_14720 = v_14721 & vout_canPeek_14731;
  assign v_14721 = ~vout_canPeek_14722;
  pebbles_core
    pebbles_core_14722
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14723),
       .in0_consume_en(vin0_consume_en_14722),
       .out_canPeek(vout_canPeek_14722),
       .out_peek(vout_peek_14722));
  assign v_14723 = v_14724 | v_14729;
  assign v_14724 = mux_14724(v_14725);
  assign v_14725 = vout_canPeek_14722 & v_14726;
  assign v_14726 = v_14727 & 1'h1;
  assign v_14727 = v_14728 | 1'h0;
  assign v_14728 = ~v_14715;
  assign v_14729 = mux_14729(v_14730);
  assign v_14730 = ~v_14725;
  pebbles_core
    pebbles_core_14731
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14732),
       .in0_consume_en(vin0_consume_en_14731),
       .out_canPeek(vout_canPeek_14731),
       .out_peek(vout_peek_14731));
  assign v_14732 = v_14733 | v_14734;
  assign v_14733 = mux_14733(v_14719);
  assign v_14734 = mux_14734(v_14735);
  assign v_14735 = ~v_14719;
  assign v_14736 = v_14737 & 1'h1;
  assign v_14737 = v_14738 & v_14739;
  assign v_14738 = ~act_14718;
  assign v_14739 = v_14740 | v_14744;
  assign v_14740 = v_14741 | v_14742;
  assign v_14741 = mux_14741(v_14675);
  assign v_14742 = mux_14742(v_14743);
  assign v_14743 = ~v_14675;
  assign v_14744 = ~v_14715;
  assign v_14745 = v_14746 | v_14747;
  assign v_14746 = mux_14746(v_14717);
  assign v_14747 = mux_14747(v_14736);
  assign v_14748 = v_14749 & 1'h1;
  assign v_14749 = v_14750 & v_14751;
  assign v_14750 = ~act_14674;
  assign v_14751 = v_14752 | v_14760;
  assign v_14752 = v_14753 | v_14758;
  assign v_14753 = mux_14753(v_14754);
  assign v_14754 = v_14671 & v_14755;
  assign v_14755 = v_14756 & 1'h1;
  assign v_14756 = v_14757 | 1'h0;
  assign v_14757 = ~v_14664;
  assign v_14758 = mux_14758(v_14759);
  assign v_14759 = ~v_14754;
  assign v_14760 = ~v_14671;
  assign v_14761 = v_14762 | v_14763;
  assign v_14762 = mux_14762(v_14673);
  assign v_14763 = mux_14763(v_14748);
  assign v_14765 = v_14766 | v_14841;
  assign v_14766 = act_14767 & 1'h1;
  assign act_14767 = v_14768 | v_14798;
  assign v_14768 = v_14769 & v_14799;
  assign v_14769 = v_14770 & v_14808;
  assign v_14770 = ~v_14771;
  assign v_14772 = v_14773 | v_14792;
  assign v_14773 = act_14774 & 1'h1;
  assign act_14774 = v_14775 | v_14781;
  assign v_14775 = v_14776 & v_14782;
  assign v_14776 = v_14777 & vout_canPeek_14787;
  assign v_14777 = ~vout_canPeek_14778;
  pebbles_core
    pebbles_core_14778
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14779),
       .in0_consume_en(vin0_consume_en_14778),
       .out_canPeek(vout_canPeek_14778),
       .out_peek(vout_peek_14778));
  assign v_14779 = v_14780 | v_14785;
  assign v_14780 = mux_14780(v_14781);
  assign v_14781 = vout_canPeek_14778 & v_14782;
  assign v_14782 = v_14783 & 1'h1;
  assign v_14783 = v_14784 | 1'h0;
  assign v_14784 = ~v_14771;
  assign v_14785 = mux_14785(v_14786);
  assign v_14786 = ~v_14781;
  pebbles_core
    pebbles_core_14787
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14788),
       .in0_consume_en(vin0_consume_en_14787),
       .out_canPeek(vout_canPeek_14787),
       .out_peek(vout_peek_14787));
  assign v_14788 = v_14789 | v_14790;
  assign v_14789 = mux_14789(v_14775);
  assign v_14790 = mux_14790(v_14791);
  assign v_14791 = ~v_14775;
  assign v_14792 = v_14793 & 1'h1;
  assign v_14793 = v_14794 & v_14795;
  assign v_14794 = ~act_14774;
  assign v_14795 = v_14796 | v_14804;
  assign v_14796 = v_14797 | v_14802;
  assign v_14797 = mux_14797(v_14798);
  assign v_14798 = v_14771 & v_14799;
  assign v_14799 = v_14800 & 1'h1;
  assign v_14800 = v_14801 | 1'h0;
  assign v_14801 = ~v_14764;
  assign v_14802 = mux_14802(v_14803);
  assign v_14803 = ~v_14798;
  assign v_14804 = ~v_14771;
  assign v_14805 = v_14806 | v_14807;
  assign v_14806 = mux_14806(v_14773);
  assign v_14807 = mux_14807(v_14792);
  assign v_14809 = v_14810 | v_14829;
  assign v_14810 = act_14811 & 1'h1;
  assign act_14811 = v_14812 | v_14818;
  assign v_14812 = v_14813 & v_14819;
  assign v_14813 = v_14814 & vout_canPeek_14824;
  assign v_14814 = ~vout_canPeek_14815;
  pebbles_core
    pebbles_core_14815
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14816),
       .in0_consume_en(vin0_consume_en_14815),
       .out_canPeek(vout_canPeek_14815),
       .out_peek(vout_peek_14815));
  assign v_14816 = v_14817 | v_14822;
  assign v_14817 = mux_14817(v_14818);
  assign v_14818 = vout_canPeek_14815 & v_14819;
  assign v_14819 = v_14820 & 1'h1;
  assign v_14820 = v_14821 | 1'h0;
  assign v_14821 = ~v_14808;
  assign v_14822 = mux_14822(v_14823);
  assign v_14823 = ~v_14818;
  pebbles_core
    pebbles_core_14824
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14825),
       .in0_consume_en(vin0_consume_en_14824),
       .out_canPeek(vout_canPeek_14824),
       .out_peek(vout_peek_14824));
  assign v_14825 = v_14826 | v_14827;
  assign v_14826 = mux_14826(v_14812);
  assign v_14827 = mux_14827(v_14828);
  assign v_14828 = ~v_14812;
  assign v_14829 = v_14830 & 1'h1;
  assign v_14830 = v_14831 & v_14832;
  assign v_14831 = ~act_14811;
  assign v_14832 = v_14833 | v_14837;
  assign v_14833 = v_14834 | v_14835;
  assign v_14834 = mux_14834(v_14768);
  assign v_14835 = mux_14835(v_14836);
  assign v_14836 = ~v_14768;
  assign v_14837 = ~v_14808;
  assign v_14838 = v_14839 | v_14840;
  assign v_14839 = mux_14839(v_14810);
  assign v_14840 = mux_14840(v_14829);
  assign v_14841 = v_14842 & 1'h1;
  assign v_14842 = v_14843 & v_14844;
  assign v_14843 = ~act_14767;
  assign v_14844 = v_14845 | v_14849;
  assign v_14845 = v_14846 | v_14847;
  assign v_14846 = mux_14846(v_14668);
  assign v_14847 = mux_14847(v_14848);
  assign v_14848 = ~v_14668;
  assign v_14849 = ~v_14764;
  assign v_14850 = v_14851 | v_14852;
  assign v_14851 = mux_14851(v_14766);
  assign v_14852 = mux_14852(v_14841);
  assign v_14853 = v_14854 & 1'h1;
  assign v_14854 = v_14855 & v_14856;
  assign v_14855 = ~act_14667;
  assign v_14856 = v_14857 | v_14865;
  assign v_14857 = v_14858 | v_14863;
  assign v_14858 = mux_14858(v_14859);
  assign v_14859 = v_14664 & v_14860;
  assign v_14860 = v_14861 & 1'h1;
  assign v_14861 = v_14862 | 1'h0;
  assign v_14862 = ~v_14657;
  assign v_14863 = mux_14863(v_14864);
  assign v_14864 = ~v_14859;
  assign v_14865 = ~v_14664;
  assign v_14866 = v_14867 | v_14868;
  assign v_14867 = mux_14867(v_14666);
  assign v_14868 = mux_14868(v_14853);
  assign v_14870 = v_14871 | v_15058;
  assign v_14871 = act_14872 & 1'h1;
  assign act_14872 = v_14873 | v_14959;
  assign v_14873 = v_14874 & v_14960;
  assign v_14874 = v_14875 & v_14969;
  assign v_14875 = ~v_14876;
  assign v_14877 = v_14878 | v_14953;
  assign v_14878 = act_14879 & 1'h1;
  assign act_14879 = v_14880 | v_14910;
  assign v_14880 = v_14881 & v_14911;
  assign v_14881 = v_14882 & v_14920;
  assign v_14882 = ~v_14883;
  assign v_14884 = v_14885 | v_14904;
  assign v_14885 = act_14886 & 1'h1;
  assign act_14886 = v_14887 | v_14893;
  assign v_14887 = v_14888 & v_14894;
  assign v_14888 = v_14889 & vout_canPeek_14899;
  assign v_14889 = ~vout_canPeek_14890;
  pebbles_core
    pebbles_core_14890
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14891),
       .in0_consume_en(vin0_consume_en_14890),
       .out_canPeek(vout_canPeek_14890),
       .out_peek(vout_peek_14890));
  assign v_14891 = v_14892 | v_14897;
  assign v_14892 = mux_14892(v_14893);
  assign v_14893 = vout_canPeek_14890 & v_14894;
  assign v_14894 = v_14895 & 1'h1;
  assign v_14895 = v_14896 | 1'h0;
  assign v_14896 = ~v_14883;
  assign v_14897 = mux_14897(v_14898);
  assign v_14898 = ~v_14893;
  pebbles_core
    pebbles_core_14899
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14900),
       .in0_consume_en(vin0_consume_en_14899),
       .out_canPeek(vout_canPeek_14899),
       .out_peek(vout_peek_14899));
  assign v_14900 = v_14901 | v_14902;
  assign v_14901 = mux_14901(v_14887);
  assign v_14902 = mux_14902(v_14903);
  assign v_14903 = ~v_14887;
  assign v_14904 = v_14905 & 1'h1;
  assign v_14905 = v_14906 & v_14907;
  assign v_14906 = ~act_14886;
  assign v_14907 = v_14908 | v_14916;
  assign v_14908 = v_14909 | v_14914;
  assign v_14909 = mux_14909(v_14910);
  assign v_14910 = v_14883 & v_14911;
  assign v_14911 = v_14912 & 1'h1;
  assign v_14912 = v_14913 | 1'h0;
  assign v_14913 = ~v_14876;
  assign v_14914 = mux_14914(v_14915);
  assign v_14915 = ~v_14910;
  assign v_14916 = ~v_14883;
  assign v_14917 = v_14918 | v_14919;
  assign v_14918 = mux_14918(v_14885);
  assign v_14919 = mux_14919(v_14904);
  assign v_14921 = v_14922 | v_14941;
  assign v_14922 = act_14923 & 1'h1;
  assign act_14923 = v_14924 | v_14930;
  assign v_14924 = v_14925 & v_14931;
  assign v_14925 = v_14926 & vout_canPeek_14936;
  assign v_14926 = ~vout_canPeek_14927;
  pebbles_core
    pebbles_core_14927
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14928),
       .in0_consume_en(vin0_consume_en_14927),
       .out_canPeek(vout_canPeek_14927),
       .out_peek(vout_peek_14927));
  assign v_14928 = v_14929 | v_14934;
  assign v_14929 = mux_14929(v_14930);
  assign v_14930 = vout_canPeek_14927 & v_14931;
  assign v_14931 = v_14932 & 1'h1;
  assign v_14932 = v_14933 | 1'h0;
  assign v_14933 = ~v_14920;
  assign v_14934 = mux_14934(v_14935);
  assign v_14935 = ~v_14930;
  pebbles_core
    pebbles_core_14936
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14937),
       .in0_consume_en(vin0_consume_en_14936),
       .out_canPeek(vout_canPeek_14936),
       .out_peek(vout_peek_14936));
  assign v_14937 = v_14938 | v_14939;
  assign v_14938 = mux_14938(v_14924);
  assign v_14939 = mux_14939(v_14940);
  assign v_14940 = ~v_14924;
  assign v_14941 = v_14942 & 1'h1;
  assign v_14942 = v_14943 & v_14944;
  assign v_14943 = ~act_14923;
  assign v_14944 = v_14945 | v_14949;
  assign v_14945 = v_14946 | v_14947;
  assign v_14946 = mux_14946(v_14880);
  assign v_14947 = mux_14947(v_14948);
  assign v_14948 = ~v_14880;
  assign v_14949 = ~v_14920;
  assign v_14950 = v_14951 | v_14952;
  assign v_14951 = mux_14951(v_14922);
  assign v_14952 = mux_14952(v_14941);
  assign v_14953 = v_14954 & 1'h1;
  assign v_14954 = v_14955 & v_14956;
  assign v_14955 = ~act_14879;
  assign v_14956 = v_14957 | v_14965;
  assign v_14957 = v_14958 | v_14963;
  assign v_14958 = mux_14958(v_14959);
  assign v_14959 = v_14876 & v_14960;
  assign v_14960 = v_14961 & 1'h1;
  assign v_14961 = v_14962 | 1'h0;
  assign v_14962 = ~v_14869;
  assign v_14963 = mux_14963(v_14964);
  assign v_14964 = ~v_14959;
  assign v_14965 = ~v_14876;
  assign v_14966 = v_14967 | v_14968;
  assign v_14967 = mux_14967(v_14878);
  assign v_14968 = mux_14968(v_14953);
  assign v_14970 = v_14971 | v_15046;
  assign v_14971 = act_14972 & 1'h1;
  assign act_14972 = v_14973 | v_15003;
  assign v_14973 = v_14974 & v_15004;
  assign v_14974 = v_14975 & v_15013;
  assign v_14975 = ~v_14976;
  assign v_14977 = v_14978 | v_14997;
  assign v_14978 = act_14979 & 1'h1;
  assign act_14979 = v_14980 | v_14986;
  assign v_14980 = v_14981 & v_14987;
  assign v_14981 = v_14982 & vout_canPeek_14992;
  assign v_14982 = ~vout_canPeek_14983;
  pebbles_core
    pebbles_core_14983
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14984),
       .in0_consume_en(vin0_consume_en_14983),
       .out_canPeek(vout_canPeek_14983),
       .out_peek(vout_peek_14983));
  assign v_14984 = v_14985 | v_14990;
  assign v_14985 = mux_14985(v_14986);
  assign v_14986 = vout_canPeek_14983 & v_14987;
  assign v_14987 = v_14988 & 1'h1;
  assign v_14988 = v_14989 | 1'h0;
  assign v_14989 = ~v_14976;
  assign v_14990 = mux_14990(v_14991);
  assign v_14991 = ~v_14986;
  pebbles_core
    pebbles_core_14992
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14993),
       .in0_consume_en(vin0_consume_en_14992),
       .out_canPeek(vout_canPeek_14992),
       .out_peek(vout_peek_14992));
  assign v_14993 = v_14994 | v_14995;
  assign v_14994 = mux_14994(v_14980);
  assign v_14995 = mux_14995(v_14996);
  assign v_14996 = ~v_14980;
  assign v_14997 = v_14998 & 1'h1;
  assign v_14998 = v_14999 & v_15000;
  assign v_14999 = ~act_14979;
  assign v_15000 = v_15001 | v_15009;
  assign v_15001 = v_15002 | v_15007;
  assign v_15002 = mux_15002(v_15003);
  assign v_15003 = v_14976 & v_15004;
  assign v_15004 = v_15005 & 1'h1;
  assign v_15005 = v_15006 | 1'h0;
  assign v_15006 = ~v_14969;
  assign v_15007 = mux_15007(v_15008);
  assign v_15008 = ~v_15003;
  assign v_15009 = ~v_14976;
  assign v_15010 = v_15011 | v_15012;
  assign v_15011 = mux_15011(v_14978);
  assign v_15012 = mux_15012(v_14997);
  assign v_15014 = v_15015 | v_15034;
  assign v_15015 = act_15016 & 1'h1;
  assign act_15016 = v_15017 | v_15023;
  assign v_15017 = v_15018 & v_15024;
  assign v_15018 = v_15019 & vout_canPeek_15029;
  assign v_15019 = ~vout_canPeek_15020;
  pebbles_core
    pebbles_core_15020
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15021),
       .in0_consume_en(vin0_consume_en_15020),
       .out_canPeek(vout_canPeek_15020),
       .out_peek(vout_peek_15020));
  assign v_15021 = v_15022 | v_15027;
  assign v_15022 = mux_15022(v_15023);
  assign v_15023 = vout_canPeek_15020 & v_15024;
  assign v_15024 = v_15025 & 1'h1;
  assign v_15025 = v_15026 | 1'h0;
  assign v_15026 = ~v_15013;
  assign v_15027 = mux_15027(v_15028);
  assign v_15028 = ~v_15023;
  pebbles_core
    pebbles_core_15029
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15030),
       .in0_consume_en(vin0_consume_en_15029),
       .out_canPeek(vout_canPeek_15029),
       .out_peek(vout_peek_15029));
  assign v_15030 = v_15031 | v_15032;
  assign v_15031 = mux_15031(v_15017);
  assign v_15032 = mux_15032(v_15033);
  assign v_15033 = ~v_15017;
  assign v_15034 = v_15035 & 1'h1;
  assign v_15035 = v_15036 & v_15037;
  assign v_15036 = ~act_15016;
  assign v_15037 = v_15038 | v_15042;
  assign v_15038 = v_15039 | v_15040;
  assign v_15039 = mux_15039(v_14973);
  assign v_15040 = mux_15040(v_15041);
  assign v_15041 = ~v_14973;
  assign v_15042 = ~v_15013;
  assign v_15043 = v_15044 | v_15045;
  assign v_15044 = mux_15044(v_15015);
  assign v_15045 = mux_15045(v_15034);
  assign v_15046 = v_15047 & 1'h1;
  assign v_15047 = v_15048 & v_15049;
  assign v_15048 = ~act_14972;
  assign v_15049 = v_15050 | v_15054;
  assign v_15050 = v_15051 | v_15052;
  assign v_15051 = mux_15051(v_14873);
  assign v_15052 = mux_15052(v_15053);
  assign v_15053 = ~v_14873;
  assign v_15054 = ~v_14969;
  assign v_15055 = v_15056 | v_15057;
  assign v_15056 = mux_15056(v_14971);
  assign v_15057 = mux_15057(v_15046);
  assign v_15058 = v_15059 & 1'h1;
  assign v_15059 = v_15060 & v_15061;
  assign v_15060 = ~act_14872;
  assign v_15061 = v_15062 | v_15066;
  assign v_15062 = v_15063 | v_15064;
  assign v_15063 = mux_15063(v_14661);
  assign v_15064 = mux_15064(v_15065);
  assign v_15065 = ~v_14661;
  assign v_15066 = ~v_14869;
  assign v_15067 = v_15068 | v_15069;
  assign v_15068 = mux_15068(v_14871);
  assign v_15069 = mux_15069(v_15058);
  assign v_15070 = v_15071 & 1'h1;
  assign v_15071 = v_15072 & v_15073;
  assign v_15072 = ~act_14660;
  assign v_15073 = v_15074 | v_15078;
  assign v_15074 = v_15075 | v_15076;
  assign v_15075 = mux_15075(v_14225);
  assign v_15076 = mux_15076(v_15077);
  assign v_15077 = ~v_14225;
  assign v_15078 = ~v_14657;
  assign v_15079 = v_15080 | v_15081;
  assign v_15080 = mux_15080(v_14659);
  assign v_15081 = mux_15081(v_15070);
  assign v_15082 = v_15083 & 1'h1;
  assign v_15083 = v_15084 & v_15085;
  assign v_15084 = ~act_14224;
  assign v_15085 = v_15086 | v_15090;
  assign v_15086 = v_15087 | v_15088;
  assign v_15087 = mux_15087(v_13341);
  assign v_15088 = mux_15088(v_15089);
  assign v_15089 = ~v_13341;
  assign v_15090 = ~v_14221;
  assign v_15091 = v_15092 | v_15093;
  assign v_15092 = mux_15092(v_14223);
  assign v_15093 = mux_15093(v_15082);
  assign v_15094 = v_15095 & 1'h1;
  assign v_15095 = v_15096 & v_15097;
  assign v_15096 = ~act_13340;
  assign v_15097 = v_15098 | v_15102;
  assign v_15098 = v_15099 | v_15100;
  assign v_15099 = mux_15099(v_11561);
  assign v_15100 = mux_15100(v_15101);
  assign v_15101 = ~v_11561;
  assign v_15102 = ~v_13337;
  assign v_15103 = v_15104 | v_15105;
  assign v_15104 = mux_15104(v_13339);
  assign v_15105 = mux_15105(v_15094);
  assign v_15106 = v_15107 & 1'h1;
  assign v_15107 = v_15108 & v_15109;
  assign v_15108 = ~act_11560;
  assign v_15109 = v_15110 | v_15114;
  assign v_15110 = v_15111 | v_15112;
  assign v_15111 = mux_15111(v_7989);
  assign v_15112 = mux_15112(v_15113);
  assign v_15113 = ~v_7989;
  assign v_15114 = ~v_11557;
  assign v_15115 = v_15116 | v_15117;
  assign v_15116 = mux_15116(v_11559);
  assign v_15117 = mux_15117(v_15106);
  assign v_15118 = v_15119 & 1'h1;
  assign v_15119 = v_15120 & v_15121;
  assign v_15120 = ~act_7988;
  assign v_15121 = v_15122 | v_15130;
  assign v_15122 = v_15123 | v_15128;
  assign v_15123 = mux_15123(v_15124);
  assign v_15124 = v_7985 & v_15125;
  assign v_15125 = v_15126 & 1'h1;
  assign v_15126 = v_15127 | 1'h0;
  assign v_15127 = ~v_7978;
  assign v_15128 = mux_15128(v_15129);
  assign v_15129 = ~v_15124;
  assign v_15130 = ~v_7985;
  assign v_15131 = v_15132 | v_15133;
  assign v_15132 = mux_15132(v_7987);
  assign v_15133 = mux_15133(v_15118);
  assign v_15135 = v_15136 | v_22267;
  assign v_15136 = act_15137 & 1'h1;
  assign act_15137 = v_15138 | v_18696;
  assign v_15138 = v_15139 & v_18697;
  assign v_15139 = v_15140 & v_18706;
  assign v_15140 = ~v_15141;
  assign v_15142 = v_15143 | v_18690;
  assign v_15143 = act_15144 & 1'h1;
  assign act_15144 = v_15145 | v_16911;
  assign v_15145 = v_15146 & v_16912;
  assign v_15146 = v_15147 & v_16921;
  assign v_15147 = ~v_15148;
  assign v_15149 = v_15150 | v_16905;
  assign v_15150 = act_15151 & 1'h1;
  assign act_15151 = v_15152 | v_16022;
  assign v_15152 = v_15153 & v_16023;
  assign v_15153 = v_15154 & v_16032;
  assign v_15154 = ~v_15155;
  assign v_15156 = v_15157 | v_16016;
  assign v_15157 = act_15158 & 1'h1;
  assign act_15158 = v_15159 | v_15581;
  assign v_15159 = v_15160 & v_15582;
  assign v_15160 = v_15161 & v_15591;
  assign v_15161 = ~v_15162;
  assign v_15163 = v_15164 | v_15575;
  assign v_15164 = act_15165 & 1'h1;
  assign act_15165 = v_15166 | v_15364;
  assign v_15166 = v_15167 & v_15365;
  assign v_15167 = v_15168 & v_15374;
  assign v_15168 = ~v_15169;
  assign v_15170 = v_15171 | v_15358;
  assign v_15171 = act_15172 & 1'h1;
  assign act_15172 = v_15173 | v_15259;
  assign v_15173 = v_15174 & v_15260;
  assign v_15174 = v_15175 & v_15269;
  assign v_15175 = ~v_15176;
  assign v_15177 = v_15178 | v_15253;
  assign v_15178 = act_15179 & 1'h1;
  assign act_15179 = v_15180 | v_15210;
  assign v_15180 = v_15181 & v_15211;
  assign v_15181 = v_15182 & v_15220;
  assign v_15182 = ~v_15183;
  assign v_15184 = v_15185 | v_15204;
  assign v_15185 = act_15186 & 1'h1;
  assign act_15186 = v_15187 | v_15193;
  assign v_15187 = v_15188 & v_15194;
  assign v_15188 = v_15189 & vout_canPeek_15199;
  assign v_15189 = ~vout_canPeek_15190;
  pebbles_core
    pebbles_core_15190
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15191),
       .in0_consume_en(vin0_consume_en_15190),
       .out_canPeek(vout_canPeek_15190),
       .out_peek(vout_peek_15190));
  assign v_15191 = v_15192 | v_15197;
  assign v_15192 = mux_15192(v_15193);
  assign v_15193 = vout_canPeek_15190 & v_15194;
  assign v_15194 = v_15195 & 1'h1;
  assign v_15195 = v_15196 | 1'h0;
  assign v_15196 = ~v_15183;
  assign v_15197 = mux_15197(v_15198);
  assign v_15198 = ~v_15193;
  pebbles_core
    pebbles_core_15199
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15200),
       .in0_consume_en(vin0_consume_en_15199),
       .out_canPeek(vout_canPeek_15199),
       .out_peek(vout_peek_15199));
  assign v_15200 = v_15201 | v_15202;
  assign v_15201 = mux_15201(v_15187);
  assign v_15202 = mux_15202(v_15203);
  assign v_15203 = ~v_15187;
  assign v_15204 = v_15205 & 1'h1;
  assign v_15205 = v_15206 & v_15207;
  assign v_15206 = ~act_15186;
  assign v_15207 = v_15208 | v_15216;
  assign v_15208 = v_15209 | v_15214;
  assign v_15209 = mux_15209(v_15210);
  assign v_15210 = v_15183 & v_15211;
  assign v_15211 = v_15212 & 1'h1;
  assign v_15212 = v_15213 | 1'h0;
  assign v_15213 = ~v_15176;
  assign v_15214 = mux_15214(v_15215);
  assign v_15215 = ~v_15210;
  assign v_15216 = ~v_15183;
  assign v_15217 = v_15218 | v_15219;
  assign v_15218 = mux_15218(v_15185);
  assign v_15219 = mux_15219(v_15204);
  assign v_15221 = v_15222 | v_15241;
  assign v_15222 = act_15223 & 1'h1;
  assign act_15223 = v_15224 | v_15230;
  assign v_15224 = v_15225 & v_15231;
  assign v_15225 = v_15226 & vout_canPeek_15236;
  assign v_15226 = ~vout_canPeek_15227;
  pebbles_core
    pebbles_core_15227
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15228),
       .in0_consume_en(vin0_consume_en_15227),
       .out_canPeek(vout_canPeek_15227),
       .out_peek(vout_peek_15227));
  assign v_15228 = v_15229 | v_15234;
  assign v_15229 = mux_15229(v_15230);
  assign v_15230 = vout_canPeek_15227 & v_15231;
  assign v_15231 = v_15232 & 1'h1;
  assign v_15232 = v_15233 | 1'h0;
  assign v_15233 = ~v_15220;
  assign v_15234 = mux_15234(v_15235);
  assign v_15235 = ~v_15230;
  pebbles_core
    pebbles_core_15236
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15237),
       .in0_consume_en(vin0_consume_en_15236),
       .out_canPeek(vout_canPeek_15236),
       .out_peek(vout_peek_15236));
  assign v_15237 = v_15238 | v_15239;
  assign v_15238 = mux_15238(v_15224);
  assign v_15239 = mux_15239(v_15240);
  assign v_15240 = ~v_15224;
  assign v_15241 = v_15242 & 1'h1;
  assign v_15242 = v_15243 & v_15244;
  assign v_15243 = ~act_15223;
  assign v_15244 = v_15245 | v_15249;
  assign v_15245 = v_15246 | v_15247;
  assign v_15246 = mux_15246(v_15180);
  assign v_15247 = mux_15247(v_15248);
  assign v_15248 = ~v_15180;
  assign v_15249 = ~v_15220;
  assign v_15250 = v_15251 | v_15252;
  assign v_15251 = mux_15251(v_15222);
  assign v_15252 = mux_15252(v_15241);
  assign v_15253 = v_15254 & 1'h1;
  assign v_15254 = v_15255 & v_15256;
  assign v_15255 = ~act_15179;
  assign v_15256 = v_15257 | v_15265;
  assign v_15257 = v_15258 | v_15263;
  assign v_15258 = mux_15258(v_15259);
  assign v_15259 = v_15176 & v_15260;
  assign v_15260 = v_15261 & 1'h1;
  assign v_15261 = v_15262 | 1'h0;
  assign v_15262 = ~v_15169;
  assign v_15263 = mux_15263(v_15264);
  assign v_15264 = ~v_15259;
  assign v_15265 = ~v_15176;
  assign v_15266 = v_15267 | v_15268;
  assign v_15267 = mux_15267(v_15178);
  assign v_15268 = mux_15268(v_15253);
  assign v_15270 = v_15271 | v_15346;
  assign v_15271 = act_15272 & 1'h1;
  assign act_15272 = v_15273 | v_15303;
  assign v_15273 = v_15274 & v_15304;
  assign v_15274 = v_15275 & v_15313;
  assign v_15275 = ~v_15276;
  assign v_15277 = v_15278 | v_15297;
  assign v_15278 = act_15279 & 1'h1;
  assign act_15279 = v_15280 | v_15286;
  assign v_15280 = v_15281 & v_15287;
  assign v_15281 = v_15282 & vout_canPeek_15292;
  assign v_15282 = ~vout_canPeek_15283;
  pebbles_core
    pebbles_core_15283
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15284),
       .in0_consume_en(vin0_consume_en_15283),
       .out_canPeek(vout_canPeek_15283),
       .out_peek(vout_peek_15283));
  assign v_15284 = v_15285 | v_15290;
  assign v_15285 = mux_15285(v_15286);
  assign v_15286 = vout_canPeek_15283 & v_15287;
  assign v_15287 = v_15288 & 1'h1;
  assign v_15288 = v_15289 | 1'h0;
  assign v_15289 = ~v_15276;
  assign v_15290 = mux_15290(v_15291);
  assign v_15291 = ~v_15286;
  pebbles_core
    pebbles_core_15292
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15293),
       .in0_consume_en(vin0_consume_en_15292),
       .out_canPeek(vout_canPeek_15292),
       .out_peek(vout_peek_15292));
  assign v_15293 = v_15294 | v_15295;
  assign v_15294 = mux_15294(v_15280);
  assign v_15295 = mux_15295(v_15296);
  assign v_15296 = ~v_15280;
  assign v_15297 = v_15298 & 1'h1;
  assign v_15298 = v_15299 & v_15300;
  assign v_15299 = ~act_15279;
  assign v_15300 = v_15301 | v_15309;
  assign v_15301 = v_15302 | v_15307;
  assign v_15302 = mux_15302(v_15303);
  assign v_15303 = v_15276 & v_15304;
  assign v_15304 = v_15305 & 1'h1;
  assign v_15305 = v_15306 | 1'h0;
  assign v_15306 = ~v_15269;
  assign v_15307 = mux_15307(v_15308);
  assign v_15308 = ~v_15303;
  assign v_15309 = ~v_15276;
  assign v_15310 = v_15311 | v_15312;
  assign v_15311 = mux_15311(v_15278);
  assign v_15312 = mux_15312(v_15297);
  assign v_15314 = v_15315 | v_15334;
  assign v_15315 = act_15316 & 1'h1;
  assign act_15316 = v_15317 | v_15323;
  assign v_15317 = v_15318 & v_15324;
  assign v_15318 = v_15319 & vout_canPeek_15329;
  assign v_15319 = ~vout_canPeek_15320;
  pebbles_core
    pebbles_core_15320
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15321),
       .in0_consume_en(vin0_consume_en_15320),
       .out_canPeek(vout_canPeek_15320),
       .out_peek(vout_peek_15320));
  assign v_15321 = v_15322 | v_15327;
  assign v_15322 = mux_15322(v_15323);
  assign v_15323 = vout_canPeek_15320 & v_15324;
  assign v_15324 = v_15325 & 1'h1;
  assign v_15325 = v_15326 | 1'h0;
  assign v_15326 = ~v_15313;
  assign v_15327 = mux_15327(v_15328);
  assign v_15328 = ~v_15323;
  pebbles_core
    pebbles_core_15329
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15330),
       .in0_consume_en(vin0_consume_en_15329),
       .out_canPeek(vout_canPeek_15329),
       .out_peek(vout_peek_15329));
  assign v_15330 = v_15331 | v_15332;
  assign v_15331 = mux_15331(v_15317);
  assign v_15332 = mux_15332(v_15333);
  assign v_15333 = ~v_15317;
  assign v_15334 = v_15335 & 1'h1;
  assign v_15335 = v_15336 & v_15337;
  assign v_15336 = ~act_15316;
  assign v_15337 = v_15338 | v_15342;
  assign v_15338 = v_15339 | v_15340;
  assign v_15339 = mux_15339(v_15273);
  assign v_15340 = mux_15340(v_15341);
  assign v_15341 = ~v_15273;
  assign v_15342 = ~v_15313;
  assign v_15343 = v_15344 | v_15345;
  assign v_15344 = mux_15344(v_15315);
  assign v_15345 = mux_15345(v_15334);
  assign v_15346 = v_15347 & 1'h1;
  assign v_15347 = v_15348 & v_15349;
  assign v_15348 = ~act_15272;
  assign v_15349 = v_15350 | v_15354;
  assign v_15350 = v_15351 | v_15352;
  assign v_15351 = mux_15351(v_15173);
  assign v_15352 = mux_15352(v_15353);
  assign v_15353 = ~v_15173;
  assign v_15354 = ~v_15269;
  assign v_15355 = v_15356 | v_15357;
  assign v_15356 = mux_15356(v_15271);
  assign v_15357 = mux_15357(v_15346);
  assign v_15358 = v_15359 & 1'h1;
  assign v_15359 = v_15360 & v_15361;
  assign v_15360 = ~act_15172;
  assign v_15361 = v_15362 | v_15370;
  assign v_15362 = v_15363 | v_15368;
  assign v_15363 = mux_15363(v_15364);
  assign v_15364 = v_15169 & v_15365;
  assign v_15365 = v_15366 & 1'h1;
  assign v_15366 = v_15367 | 1'h0;
  assign v_15367 = ~v_15162;
  assign v_15368 = mux_15368(v_15369);
  assign v_15369 = ~v_15364;
  assign v_15370 = ~v_15169;
  assign v_15371 = v_15372 | v_15373;
  assign v_15372 = mux_15372(v_15171);
  assign v_15373 = mux_15373(v_15358);
  assign v_15375 = v_15376 | v_15563;
  assign v_15376 = act_15377 & 1'h1;
  assign act_15377 = v_15378 | v_15464;
  assign v_15378 = v_15379 & v_15465;
  assign v_15379 = v_15380 & v_15474;
  assign v_15380 = ~v_15381;
  assign v_15382 = v_15383 | v_15458;
  assign v_15383 = act_15384 & 1'h1;
  assign act_15384 = v_15385 | v_15415;
  assign v_15385 = v_15386 & v_15416;
  assign v_15386 = v_15387 & v_15425;
  assign v_15387 = ~v_15388;
  assign v_15389 = v_15390 | v_15409;
  assign v_15390 = act_15391 & 1'h1;
  assign act_15391 = v_15392 | v_15398;
  assign v_15392 = v_15393 & v_15399;
  assign v_15393 = v_15394 & vout_canPeek_15404;
  assign v_15394 = ~vout_canPeek_15395;
  pebbles_core
    pebbles_core_15395
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15396),
       .in0_consume_en(vin0_consume_en_15395),
       .out_canPeek(vout_canPeek_15395),
       .out_peek(vout_peek_15395));
  assign v_15396 = v_15397 | v_15402;
  assign v_15397 = mux_15397(v_15398);
  assign v_15398 = vout_canPeek_15395 & v_15399;
  assign v_15399 = v_15400 & 1'h1;
  assign v_15400 = v_15401 | 1'h0;
  assign v_15401 = ~v_15388;
  assign v_15402 = mux_15402(v_15403);
  assign v_15403 = ~v_15398;
  pebbles_core
    pebbles_core_15404
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15405),
       .in0_consume_en(vin0_consume_en_15404),
       .out_canPeek(vout_canPeek_15404),
       .out_peek(vout_peek_15404));
  assign v_15405 = v_15406 | v_15407;
  assign v_15406 = mux_15406(v_15392);
  assign v_15407 = mux_15407(v_15408);
  assign v_15408 = ~v_15392;
  assign v_15409 = v_15410 & 1'h1;
  assign v_15410 = v_15411 & v_15412;
  assign v_15411 = ~act_15391;
  assign v_15412 = v_15413 | v_15421;
  assign v_15413 = v_15414 | v_15419;
  assign v_15414 = mux_15414(v_15415);
  assign v_15415 = v_15388 & v_15416;
  assign v_15416 = v_15417 & 1'h1;
  assign v_15417 = v_15418 | 1'h0;
  assign v_15418 = ~v_15381;
  assign v_15419 = mux_15419(v_15420);
  assign v_15420 = ~v_15415;
  assign v_15421 = ~v_15388;
  assign v_15422 = v_15423 | v_15424;
  assign v_15423 = mux_15423(v_15390);
  assign v_15424 = mux_15424(v_15409);
  assign v_15426 = v_15427 | v_15446;
  assign v_15427 = act_15428 & 1'h1;
  assign act_15428 = v_15429 | v_15435;
  assign v_15429 = v_15430 & v_15436;
  assign v_15430 = v_15431 & vout_canPeek_15441;
  assign v_15431 = ~vout_canPeek_15432;
  pebbles_core
    pebbles_core_15432
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15433),
       .in0_consume_en(vin0_consume_en_15432),
       .out_canPeek(vout_canPeek_15432),
       .out_peek(vout_peek_15432));
  assign v_15433 = v_15434 | v_15439;
  assign v_15434 = mux_15434(v_15435);
  assign v_15435 = vout_canPeek_15432 & v_15436;
  assign v_15436 = v_15437 & 1'h1;
  assign v_15437 = v_15438 | 1'h0;
  assign v_15438 = ~v_15425;
  assign v_15439 = mux_15439(v_15440);
  assign v_15440 = ~v_15435;
  pebbles_core
    pebbles_core_15441
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15442),
       .in0_consume_en(vin0_consume_en_15441),
       .out_canPeek(vout_canPeek_15441),
       .out_peek(vout_peek_15441));
  assign v_15442 = v_15443 | v_15444;
  assign v_15443 = mux_15443(v_15429);
  assign v_15444 = mux_15444(v_15445);
  assign v_15445 = ~v_15429;
  assign v_15446 = v_15447 & 1'h1;
  assign v_15447 = v_15448 & v_15449;
  assign v_15448 = ~act_15428;
  assign v_15449 = v_15450 | v_15454;
  assign v_15450 = v_15451 | v_15452;
  assign v_15451 = mux_15451(v_15385);
  assign v_15452 = mux_15452(v_15453);
  assign v_15453 = ~v_15385;
  assign v_15454 = ~v_15425;
  assign v_15455 = v_15456 | v_15457;
  assign v_15456 = mux_15456(v_15427);
  assign v_15457 = mux_15457(v_15446);
  assign v_15458 = v_15459 & 1'h1;
  assign v_15459 = v_15460 & v_15461;
  assign v_15460 = ~act_15384;
  assign v_15461 = v_15462 | v_15470;
  assign v_15462 = v_15463 | v_15468;
  assign v_15463 = mux_15463(v_15464);
  assign v_15464 = v_15381 & v_15465;
  assign v_15465 = v_15466 & 1'h1;
  assign v_15466 = v_15467 | 1'h0;
  assign v_15467 = ~v_15374;
  assign v_15468 = mux_15468(v_15469);
  assign v_15469 = ~v_15464;
  assign v_15470 = ~v_15381;
  assign v_15471 = v_15472 | v_15473;
  assign v_15472 = mux_15472(v_15383);
  assign v_15473 = mux_15473(v_15458);
  assign v_15475 = v_15476 | v_15551;
  assign v_15476 = act_15477 & 1'h1;
  assign act_15477 = v_15478 | v_15508;
  assign v_15478 = v_15479 & v_15509;
  assign v_15479 = v_15480 & v_15518;
  assign v_15480 = ~v_15481;
  assign v_15482 = v_15483 | v_15502;
  assign v_15483 = act_15484 & 1'h1;
  assign act_15484 = v_15485 | v_15491;
  assign v_15485 = v_15486 & v_15492;
  assign v_15486 = v_15487 & vout_canPeek_15497;
  assign v_15487 = ~vout_canPeek_15488;
  pebbles_core
    pebbles_core_15488
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15489),
       .in0_consume_en(vin0_consume_en_15488),
       .out_canPeek(vout_canPeek_15488),
       .out_peek(vout_peek_15488));
  assign v_15489 = v_15490 | v_15495;
  assign v_15490 = mux_15490(v_15491);
  assign v_15491 = vout_canPeek_15488 & v_15492;
  assign v_15492 = v_15493 & 1'h1;
  assign v_15493 = v_15494 | 1'h0;
  assign v_15494 = ~v_15481;
  assign v_15495 = mux_15495(v_15496);
  assign v_15496 = ~v_15491;
  pebbles_core
    pebbles_core_15497
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15498),
       .in0_consume_en(vin0_consume_en_15497),
       .out_canPeek(vout_canPeek_15497),
       .out_peek(vout_peek_15497));
  assign v_15498 = v_15499 | v_15500;
  assign v_15499 = mux_15499(v_15485);
  assign v_15500 = mux_15500(v_15501);
  assign v_15501 = ~v_15485;
  assign v_15502 = v_15503 & 1'h1;
  assign v_15503 = v_15504 & v_15505;
  assign v_15504 = ~act_15484;
  assign v_15505 = v_15506 | v_15514;
  assign v_15506 = v_15507 | v_15512;
  assign v_15507 = mux_15507(v_15508);
  assign v_15508 = v_15481 & v_15509;
  assign v_15509 = v_15510 & 1'h1;
  assign v_15510 = v_15511 | 1'h0;
  assign v_15511 = ~v_15474;
  assign v_15512 = mux_15512(v_15513);
  assign v_15513 = ~v_15508;
  assign v_15514 = ~v_15481;
  assign v_15515 = v_15516 | v_15517;
  assign v_15516 = mux_15516(v_15483);
  assign v_15517 = mux_15517(v_15502);
  assign v_15519 = v_15520 | v_15539;
  assign v_15520 = act_15521 & 1'h1;
  assign act_15521 = v_15522 | v_15528;
  assign v_15522 = v_15523 & v_15529;
  assign v_15523 = v_15524 & vout_canPeek_15534;
  assign v_15524 = ~vout_canPeek_15525;
  pebbles_core
    pebbles_core_15525
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15526),
       .in0_consume_en(vin0_consume_en_15525),
       .out_canPeek(vout_canPeek_15525),
       .out_peek(vout_peek_15525));
  assign v_15526 = v_15527 | v_15532;
  assign v_15527 = mux_15527(v_15528);
  assign v_15528 = vout_canPeek_15525 & v_15529;
  assign v_15529 = v_15530 & 1'h1;
  assign v_15530 = v_15531 | 1'h0;
  assign v_15531 = ~v_15518;
  assign v_15532 = mux_15532(v_15533);
  assign v_15533 = ~v_15528;
  pebbles_core
    pebbles_core_15534
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15535),
       .in0_consume_en(vin0_consume_en_15534),
       .out_canPeek(vout_canPeek_15534),
       .out_peek(vout_peek_15534));
  assign v_15535 = v_15536 | v_15537;
  assign v_15536 = mux_15536(v_15522);
  assign v_15537 = mux_15537(v_15538);
  assign v_15538 = ~v_15522;
  assign v_15539 = v_15540 & 1'h1;
  assign v_15540 = v_15541 & v_15542;
  assign v_15541 = ~act_15521;
  assign v_15542 = v_15543 | v_15547;
  assign v_15543 = v_15544 | v_15545;
  assign v_15544 = mux_15544(v_15478);
  assign v_15545 = mux_15545(v_15546);
  assign v_15546 = ~v_15478;
  assign v_15547 = ~v_15518;
  assign v_15548 = v_15549 | v_15550;
  assign v_15549 = mux_15549(v_15520);
  assign v_15550 = mux_15550(v_15539);
  assign v_15551 = v_15552 & 1'h1;
  assign v_15552 = v_15553 & v_15554;
  assign v_15553 = ~act_15477;
  assign v_15554 = v_15555 | v_15559;
  assign v_15555 = v_15556 | v_15557;
  assign v_15556 = mux_15556(v_15378);
  assign v_15557 = mux_15557(v_15558);
  assign v_15558 = ~v_15378;
  assign v_15559 = ~v_15474;
  assign v_15560 = v_15561 | v_15562;
  assign v_15561 = mux_15561(v_15476);
  assign v_15562 = mux_15562(v_15551);
  assign v_15563 = v_15564 & 1'h1;
  assign v_15564 = v_15565 & v_15566;
  assign v_15565 = ~act_15377;
  assign v_15566 = v_15567 | v_15571;
  assign v_15567 = v_15568 | v_15569;
  assign v_15568 = mux_15568(v_15166);
  assign v_15569 = mux_15569(v_15570);
  assign v_15570 = ~v_15166;
  assign v_15571 = ~v_15374;
  assign v_15572 = v_15573 | v_15574;
  assign v_15573 = mux_15573(v_15376);
  assign v_15574 = mux_15574(v_15563);
  assign v_15575 = v_15576 & 1'h1;
  assign v_15576 = v_15577 & v_15578;
  assign v_15577 = ~act_15165;
  assign v_15578 = v_15579 | v_15587;
  assign v_15579 = v_15580 | v_15585;
  assign v_15580 = mux_15580(v_15581);
  assign v_15581 = v_15162 & v_15582;
  assign v_15582 = v_15583 & 1'h1;
  assign v_15583 = v_15584 | 1'h0;
  assign v_15584 = ~v_15155;
  assign v_15585 = mux_15585(v_15586);
  assign v_15586 = ~v_15581;
  assign v_15587 = ~v_15162;
  assign v_15588 = v_15589 | v_15590;
  assign v_15589 = mux_15589(v_15164);
  assign v_15590 = mux_15590(v_15575);
  assign v_15592 = v_15593 | v_16004;
  assign v_15593 = act_15594 & 1'h1;
  assign act_15594 = v_15595 | v_15793;
  assign v_15595 = v_15596 & v_15794;
  assign v_15596 = v_15597 & v_15803;
  assign v_15597 = ~v_15598;
  assign v_15599 = v_15600 | v_15787;
  assign v_15600 = act_15601 & 1'h1;
  assign act_15601 = v_15602 | v_15688;
  assign v_15602 = v_15603 & v_15689;
  assign v_15603 = v_15604 & v_15698;
  assign v_15604 = ~v_15605;
  assign v_15606 = v_15607 | v_15682;
  assign v_15607 = act_15608 & 1'h1;
  assign act_15608 = v_15609 | v_15639;
  assign v_15609 = v_15610 & v_15640;
  assign v_15610 = v_15611 & v_15649;
  assign v_15611 = ~v_15612;
  assign v_15613 = v_15614 | v_15633;
  assign v_15614 = act_15615 & 1'h1;
  assign act_15615 = v_15616 | v_15622;
  assign v_15616 = v_15617 & v_15623;
  assign v_15617 = v_15618 & vout_canPeek_15628;
  assign v_15618 = ~vout_canPeek_15619;
  pebbles_core
    pebbles_core_15619
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15620),
       .in0_consume_en(vin0_consume_en_15619),
       .out_canPeek(vout_canPeek_15619),
       .out_peek(vout_peek_15619));
  assign v_15620 = v_15621 | v_15626;
  assign v_15621 = mux_15621(v_15622);
  assign v_15622 = vout_canPeek_15619 & v_15623;
  assign v_15623 = v_15624 & 1'h1;
  assign v_15624 = v_15625 | 1'h0;
  assign v_15625 = ~v_15612;
  assign v_15626 = mux_15626(v_15627);
  assign v_15627 = ~v_15622;
  pebbles_core
    pebbles_core_15628
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15629),
       .in0_consume_en(vin0_consume_en_15628),
       .out_canPeek(vout_canPeek_15628),
       .out_peek(vout_peek_15628));
  assign v_15629 = v_15630 | v_15631;
  assign v_15630 = mux_15630(v_15616);
  assign v_15631 = mux_15631(v_15632);
  assign v_15632 = ~v_15616;
  assign v_15633 = v_15634 & 1'h1;
  assign v_15634 = v_15635 & v_15636;
  assign v_15635 = ~act_15615;
  assign v_15636 = v_15637 | v_15645;
  assign v_15637 = v_15638 | v_15643;
  assign v_15638 = mux_15638(v_15639);
  assign v_15639 = v_15612 & v_15640;
  assign v_15640 = v_15641 & 1'h1;
  assign v_15641 = v_15642 | 1'h0;
  assign v_15642 = ~v_15605;
  assign v_15643 = mux_15643(v_15644);
  assign v_15644 = ~v_15639;
  assign v_15645 = ~v_15612;
  assign v_15646 = v_15647 | v_15648;
  assign v_15647 = mux_15647(v_15614);
  assign v_15648 = mux_15648(v_15633);
  assign v_15650 = v_15651 | v_15670;
  assign v_15651 = act_15652 & 1'h1;
  assign act_15652 = v_15653 | v_15659;
  assign v_15653 = v_15654 & v_15660;
  assign v_15654 = v_15655 & vout_canPeek_15665;
  assign v_15655 = ~vout_canPeek_15656;
  pebbles_core
    pebbles_core_15656
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15657),
       .in0_consume_en(vin0_consume_en_15656),
       .out_canPeek(vout_canPeek_15656),
       .out_peek(vout_peek_15656));
  assign v_15657 = v_15658 | v_15663;
  assign v_15658 = mux_15658(v_15659);
  assign v_15659 = vout_canPeek_15656 & v_15660;
  assign v_15660 = v_15661 & 1'h1;
  assign v_15661 = v_15662 | 1'h0;
  assign v_15662 = ~v_15649;
  assign v_15663 = mux_15663(v_15664);
  assign v_15664 = ~v_15659;
  pebbles_core
    pebbles_core_15665
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15666),
       .in0_consume_en(vin0_consume_en_15665),
       .out_canPeek(vout_canPeek_15665),
       .out_peek(vout_peek_15665));
  assign v_15666 = v_15667 | v_15668;
  assign v_15667 = mux_15667(v_15653);
  assign v_15668 = mux_15668(v_15669);
  assign v_15669 = ~v_15653;
  assign v_15670 = v_15671 & 1'h1;
  assign v_15671 = v_15672 & v_15673;
  assign v_15672 = ~act_15652;
  assign v_15673 = v_15674 | v_15678;
  assign v_15674 = v_15675 | v_15676;
  assign v_15675 = mux_15675(v_15609);
  assign v_15676 = mux_15676(v_15677);
  assign v_15677 = ~v_15609;
  assign v_15678 = ~v_15649;
  assign v_15679 = v_15680 | v_15681;
  assign v_15680 = mux_15680(v_15651);
  assign v_15681 = mux_15681(v_15670);
  assign v_15682 = v_15683 & 1'h1;
  assign v_15683 = v_15684 & v_15685;
  assign v_15684 = ~act_15608;
  assign v_15685 = v_15686 | v_15694;
  assign v_15686 = v_15687 | v_15692;
  assign v_15687 = mux_15687(v_15688);
  assign v_15688 = v_15605 & v_15689;
  assign v_15689 = v_15690 & 1'h1;
  assign v_15690 = v_15691 | 1'h0;
  assign v_15691 = ~v_15598;
  assign v_15692 = mux_15692(v_15693);
  assign v_15693 = ~v_15688;
  assign v_15694 = ~v_15605;
  assign v_15695 = v_15696 | v_15697;
  assign v_15696 = mux_15696(v_15607);
  assign v_15697 = mux_15697(v_15682);
  assign v_15699 = v_15700 | v_15775;
  assign v_15700 = act_15701 & 1'h1;
  assign act_15701 = v_15702 | v_15732;
  assign v_15702 = v_15703 & v_15733;
  assign v_15703 = v_15704 & v_15742;
  assign v_15704 = ~v_15705;
  assign v_15706 = v_15707 | v_15726;
  assign v_15707 = act_15708 & 1'h1;
  assign act_15708 = v_15709 | v_15715;
  assign v_15709 = v_15710 & v_15716;
  assign v_15710 = v_15711 & vout_canPeek_15721;
  assign v_15711 = ~vout_canPeek_15712;
  pebbles_core
    pebbles_core_15712
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15713),
       .in0_consume_en(vin0_consume_en_15712),
       .out_canPeek(vout_canPeek_15712),
       .out_peek(vout_peek_15712));
  assign v_15713 = v_15714 | v_15719;
  assign v_15714 = mux_15714(v_15715);
  assign v_15715 = vout_canPeek_15712 & v_15716;
  assign v_15716 = v_15717 & 1'h1;
  assign v_15717 = v_15718 | 1'h0;
  assign v_15718 = ~v_15705;
  assign v_15719 = mux_15719(v_15720);
  assign v_15720 = ~v_15715;
  pebbles_core
    pebbles_core_15721
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15722),
       .in0_consume_en(vin0_consume_en_15721),
       .out_canPeek(vout_canPeek_15721),
       .out_peek(vout_peek_15721));
  assign v_15722 = v_15723 | v_15724;
  assign v_15723 = mux_15723(v_15709);
  assign v_15724 = mux_15724(v_15725);
  assign v_15725 = ~v_15709;
  assign v_15726 = v_15727 & 1'h1;
  assign v_15727 = v_15728 & v_15729;
  assign v_15728 = ~act_15708;
  assign v_15729 = v_15730 | v_15738;
  assign v_15730 = v_15731 | v_15736;
  assign v_15731 = mux_15731(v_15732);
  assign v_15732 = v_15705 & v_15733;
  assign v_15733 = v_15734 & 1'h1;
  assign v_15734 = v_15735 | 1'h0;
  assign v_15735 = ~v_15698;
  assign v_15736 = mux_15736(v_15737);
  assign v_15737 = ~v_15732;
  assign v_15738 = ~v_15705;
  assign v_15739 = v_15740 | v_15741;
  assign v_15740 = mux_15740(v_15707);
  assign v_15741 = mux_15741(v_15726);
  assign v_15743 = v_15744 | v_15763;
  assign v_15744 = act_15745 & 1'h1;
  assign act_15745 = v_15746 | v_15752;
  assign v_15746 = v_15747 & v_15753;
  assign v_15747 = v_15748 & vout_canPeek_15758;
  assign v_15748 = ~vout_canPeek_15749;
  pebbles_core
    pebbles_core_15749
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15750),
       .in0_consume_en(vin0_consume_en_15749),
       .out_canPeek(vout_canPeek_15749),
       .out_peek(vout_peek_15749));
  assign v_15750 = v_15751 | v_15756;
  assign v_15751 = mux_15751(v_15752);
  assign v_15752 = vout_canPeek_15749 & v_15753;
  assign v_15753 = v_15754 & 1'h1;
  assign v_15754 = v_15755 | 1'h0;
  assign v_15755 = ~v_15742;
  assign v_15756 = mux_15756(v_15757);
  assign v_15757 = ~v_15752;
  pebbles_core
    pebbles_core_15758
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15759),
       .in0_consume_en(vin0_consume_en_15758),
       .out_canPeek(vout_canPeek_15758),
       .out_peek(vout_peek_15758));
  assign v_15759 = v_15760 | v_15761;
  assign v_15760 = mux_15760(v_15746);
  assign v_15761 = mux_15761(v_15762);
  assign v_15762 = ~v_15746;
  assign v_15763 = v_15764 & 1'h1;
  assign v_15764 = v_15765 & v_15766;
  assign v_15765 = ~act_15745;
  assign v_15766 = v_15767 | v_15771;
  assign v_15767 = v_15768 | v_15769;
  assign v_15768 = mux_15768(v_15702);
  assign v_15769 = mux_15769(v_15770);
  assign v_15770 = ~v_15702;
  assign v_15771 = ~v_15742;
  assign v_15772 = v_15773 | v_15774;
  assign v_15773 = mux_15773(v_15744);
  assign v_15774 = mux_15774(v_15763);
  assign v_15775 = v_15776 & 1'h1;
  assign v_15776 = v_15777 & v_15778;
  assign v_15777 = ~act_15701;
  assign v_15778 = v_15779 | v_15783;
  assign v_15779 = v_15780 | v_15781;
  assign v_15780 = mux_15780(v_15602);
  assign v_15781 = mux_15781(v_15782);
  assign v_15782 = ~v_15602;
  assign v_15783 = ~v_15698;
  assign v_15784 = v_15785 | v_15786;
  assign v_15785 = mux_15785(v_15700);
  assign v_15786 = mux_15786(v_15775);
  assign v_15787 = v_15788 & 1'h1;
  assign v_15788 = v_15789 & v_15790;
  assign v_15789 = ~act_15601;
  assign v_15790 = v_15791 | v_15799;
  assign v_15791 = v_15792 | v_15797;
  assign v_15792 = mux_15792(v_15793);
  assign v_15793 = v_15598 & v_15794;
  assign v_15794 = v_15795 & 1'h1;
  assign v_15795 = v_15796 | 1'h0;
  assign v_15796 = ~v_15591;
  assign v_15797 = mux_15797(v_15798);
  assign v_15798 = ~v_15793;
  assign v_15799 = ~v_15598;
  assign v_15800 = v_15801 | v_15802;
  assign v_15801 = mux_15801(v_15600);
  assign v_15802 = mux_15802(v_15787);
  assign v_15804 = v_15805 | v_15992;
  assign v_15805 = act_15806 & 1'h1;
  assign act_15806 = v_15807 | v_15893;
  assign v_15807 = v_15808 & v_15894;
  assign v_15808 = v_15809 & v_15903;
  assign v_15809 = ~v_15810;
  assign v_15811 = v_15812 | v_15887;
  assign v_15812 = act_15813 & 1'h1;
  assign act_15813 = v_15814 | v_15844;
  assign v_15814 = v_15815 & v_15845;
  assign v_15815 = v_15816 & v_15854;
  assign v_15816 = ~v_15817;
  assign v_15818 = v_15819 | v_15838;
  assign v_15819 = act_15820 & 1'h1;
  assign act_15820 = v_15821 | v_15827;
  assign v_15821 = v_15822 & v_15828;
  assign v_15822 = v_15823 & vout_canPeek_15833;
  assign v_15823 = ~vout_canPeek_15824;
  pebbles_core
    pebbles_core_15824
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15825),
       .in0_consume_en(vin0_consume_en_15824),
       .out_canPeek(vout_canPeek_15824),
       .out_peek(vout_peek_15824));
  assign v_15825 = v_15826 | v_15831;
  assign v_15826 = mux_15826(v_15827);
  assign v_15827 = vout_canPeek_15824 & v_15828;
  assign v_15828 = v_15829 & 1'h1;
  assign v_15829 = v_15830 | 1'h0;
  assign v_15830 = ~v_15817;
  assign v_15831 = mux_15831(v_15832);
  assign v_15832 = ~v_15827;
  pebbles_core
    pebbles_core_15833
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15834),
       .in0_consume_en(vin0_consume_en_15833),
       .out_canPeek(vout_canPeek_15833),
       .out_peek(vout_peek_15833));
  assign v_15834 = v_15835 | v_15836;
  assign v_15835 = mux_15835(v_15821);
  assign v_15836 = mux_15836(v_15837);
  assign v_15837 = ~v_15821;
  assign v_15838 = v_15839 & 1'h1;
  assign v_15839 = v_15840 & v_15841;
  assign v_15840 = ~act_15820;
  assign v_15841 = v_15842 | v_15850;
  assign v_15842 = v_15843 | v_15848;
  assign v_15843 = mux_15843(v_15844);
  assign v_15844 = v_15817 & v_15845;
  assign v_15845 = v_15846 & 1'h1;
  assign v_15846 = v_15847 | 1'h0;
  assign v_15847 = ~v_15810;
  assign v_15848 = mux_15848(v_15849);
  assign v_15849 = ~v_15844;
  assign v_15850 = ~v_15817;
  assign v_15851 = v_15852 | v_15853;
  assign v_15852 = mux_15852(v_15819);
  assign v_15853 = mux_15853(v_15838);
  assign v_15855 = v_15856 | v_15875;
  assign v_15856 = act_15857 & 1'h1;
  assign act_15857 = v_15858 | v_15864;
  assign v_15858 = v_15859 & v_15865;
  assign v_15859 = v_15860 & vout_canPeek_15870;
  assign v_15860 = ~vout_canPeek_15861;
  pebbles_core
    pebbles_core_15861
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15862),
       .in0_consume_en(vin0_consume_en_15861),
       .out_canPeek(vout_canPeek_15861),
       .out_peek(vout_peek_15861));
  assign v_15862 = v_15863 | v_15868;
  assign v_15863 = mux_15863(v_15864);
  assign v_15864 = vout_canPeek_15861 & v_15865;
  assign v_15865 = v_15866 & 1'h1;
  assign v_15866 = v_15867 | 1'h0;
  assign v_15867 = ~v_15854;
  assign v_15868 = mux_15868(v_15869);
  assign v_15869 = ~v_15864;
  pebbles_core
    pebbles_core_15870
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15871),
       .in0_consume_en(vin0_consume_en_15870),
       .out_canPeek(vout_canPeek_15870),
       .out_peek(vout_peek_15870));
  assign v_15871 = v_15872 | v_15873;
  assign v_15872 = mux_15872(v_15858);
  assign v_15873 = mux_15873(v_15874);
  assign v_15874 = ~v_15858;
  assign v_15875 = v_15876 & 1'h1;
  assign v_15876 = v_15877 & v_15878;
  assign v_15877 = ~act_15857;
  assign v_15878 = v_15879 | v_15883;
  assign v_15879 = v_15880 | v_15881;
  assign v_15880 = mux_15880(v_15814);
  assign v_15881 = mux_15881(v_15882);
  assign v_15882 = ~v_15814;
  assign v_15883 = ~v_15854;
  assign v_15884 = v_15885 | v_15886;
  assign v_15885 = mux_15885(v_15856);
  assign v_15886 = mux_15886(v_15875);
  assign v_15887 = v_15888 & 1'h1;
  assign v_15888 = v_15889 & v_15890;
  assign v_15889 = ~act_15813;
  assign v_15890 = v_15891 | v_15899;
  assign v_15891 = v_15892 | v_15897;
  assign v_15892 = mux_15892(v_15893);
  assign v_15893 = v_15810 & v_15894;
  assign v_15894 = v_15895 & 1'h1;
  assign v_15895 = v_15896 | 1'h0;
  assign v_15896 = ~v_15803;
  assign v_15897 = mux_15897(v_15898);
  assign v_15898 = ~v_15893;
  assign v_15899 = ~v_15810;
  assign v_15900 = v_15901 | v_15902;
  assign v_15901 = mux_15901(v_15812);
  assign v_15902 = mux_15902(v_15887);
  assign v_15904 = v_15905 | v_15980;
  assign v_15905 = act_15906 & 1'h1;
  assign act_15906 = v_15907 | v_15937;
  assign v_15907 = v_15908 & v_15938;
  assign v_15908 = v_15909 & v_15947;
  assign v_15909 = ~v_15910;
  assign v_15911 = v_15912 | v_15931;
  assign v_15912 = act_15913 & 1'h1;
  assign act_15913 = v_15914 | v_15920;
  assign v_15914 = v_15915 & v_15921;
  assign v_15915 = v_15916 & vout_canPeek_15926;
  assign v_15916 = ~vout_canPeek_15917;
  pebbles_core
    pebbles_core_15917
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15918),
       .in0_consume_en(vin0_consume_en_15917),
       .out_canPeek(vout_canPeek_15917),
       .out_peek(vout_peek_15917));
  assign v_15918 = v_15919 | v_15924;
  assign v_15919 = mux_15919(v_15920);
  assign v_15920 = vout_canPeek_15917 & v_15921;
  assign v_15921 = v_15922 & 1'h1;
  assign v_15922 = v_15923 | 1'h0;
  assign v_15923 = ~v_15910;
  assign v_15924 = mux_15924(v_15925);
  assign v_15925 = ~v_15920;
  pebbles_core
    pebbles_core_15926
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15927),
       .in0_consume_en(vin0_consume_en_15926),
       .out_canPeek(vout_canPeek_15926),
       .out_peek(vout_peek_15926));
  assign v_15927 = v_15928 | v_15929;
  assign v_15928 = mux_15928(v_15914);
  assign v_15929 = mux_15929(v_15930);
  assign v_15930 = ~v_15914;
  assign v_15931 = v_15932 & 1'h1;
  assign v_15932 = v_15933 & v_15934;
  assign v_15933 = ~act_15913;
  assign v_15934 = v_15935 | v_15943;
  assign v_15935 = v_15936 | v_15941;
  assign v_15936 = mux_15936(v_15937);
  assign v_15937 = v_15910 & v_15938;
  assign v_15938 = v_15939 & 1'h1;
  assign v_15939 = v_15940 | 1'h0;
  assign v_15940 = ~v_15903;
  assign v_15941 = mux_15941(v_15942);
  assign v_15942 = ~v_15937;
  assign v_15943 = ~v_15910;
  assign v_15944 = v_15945 | v_15946;
  assign v_15945 = mux_15945(v_15912);
  assign v_15946 = mux_15946(v_15931);
  assign v_15948 = v_15949 | v_15968;
  assign v_15949 = act_15950 & 1'h1;
  assign act_15950 = v_15951 | v_15957;
  assign v_15951 = v_15952 & v_15958;
  assign v_15952 = v_15953 & vout_canPeek_15963;
  assign v_15953 = ~vout_canPeek_15954;
  pebbles_core
    pebbles_core_15954
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15955),
       .in0_consume_en(vin0_consume_en_15954),
       .out_canPeek(vout_canPeek_15954),
       .out_peek(vout_peek_15954));
  assign v_15955 = v_15956 | v_15961;
  assign v_15956 = mux_15956(v_15957);
  assign v_15957 = vout_canPeek_15954 & v_15958;
  assign v_15958 = v_15959 & 1'h1;
  assign v_15959 = v_15960 | 1'h0;
  assign v_15960 = ~v_15947;
  assign v_15961 = mux_15961(v_15962);
  assign v_15962 = ~v_15957;
  pebbles_core
    pebbles_core_15963
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_15964),
       .in0_consume_en(vin0_consume_en_15963),
       .out_canPeek(vout_canPeek_15963),
       .out_peek(vout_peek_15963));
  assign v_15964 = v_15965 | v_15966;
  assign v_15965 = mux_15965(v_15951);
  assign v_15966 = mux_15966(v_15967);
  assign v_15967 = ~v_15951;
  assign v_15968 = v_15969 & 1'h1;
  assign v_15969 = v_15970 & v_15971;
  assign v_15970 = ~act_15950;
  assign v_15971 = v_15972 | v_15976;
  assign v_15972 = v_15973 | v_15974;
  assign v_15973 = mux_15973(v_15907);
  assign v_15974 = mux_15974(v_15975);
  assign v_15975 = ~v_15907;
  assign v_15976 = ~v_15947;
  assign v_15977 = v_15978 | v_15979;
  assign v_15978 = mux_15978(v_15949);
  assign v_15979 = mux_15979(v_15968);
  assign v_15980 = v_15981 & 1'h1;
  assign v_15981 = v_15982 & v_15983;
  assign v_15982 = ~act_15906;
  assign v_15983 = v_15984 | v_15988;
  assign v_15984 = v_15985 | v_15986;
  assign v_15985 = mux_15985(v_15807);
  assign v_15986 = mux_15986(v_15987);
  assign v_15987 = ~v_15807;
  assign v_15988 = ~v_15903;
  assign v_15989 = v_15990 | v_15991;
  assign v_15990 = mux_15990(v_15905);
  assign v_15991 = mux_15991(v_15980);
  assign v_15992 = v_15993 & 1'h1;
  assign v_15993 = v_15994 & v_15995;
  assign v_15994 = ~act_15806;
  assign v_15995 = v_15996 | v_16000;
  assign v_15996 = v_15997 | v_15998;
  assign v_15997 = mux_15997(v_15595);
  assign v_15998 = mux_15998(v_15999);
  assign v_15999 = ~v_15595;
  assign v_16000 = ~v_15803;
  assign v_16001 = v_16002 | v_16003;
  assign v_16002 = mux_16002(v_15805);
  assign v_16003 = mux_16003(v_15992);
  assign v_16004 = v_16005 & 1'h1;
  assign v_16005 = v_16006 & v_16007;
  assign v_16006 = ~act_15594;
  assign v_16007 = v_16008 | v_16012;
  assign v_16008 = v_16009 | v_16010;
  assign v_16009 = mux_16009(v_15159);
  assign v_16010 = mux_16010(v_16011);
  assign v_16011 = ~v_15159;
  assign v_16012 = ~v_15591;
  assign v_16013 = v_16014 | v_16015;
  assign v_16014 = mux_16014(v_15593);
  assign v_16015 = mux_16015(v_16004);
  assign v_16016 = v_16017 & 1'h1;
  assign v_16017 = v_16018 & v_16019;
  assign v_16018 = ~act_15158;
  assign v_16019 = v_16020 | v_16028;
  assign v_16020 = v_16021 | v_16026;
  assign v_16021 = mux_16021(v_16022);
  assign v_16022 = v_15155 & v_16023;
  assign v_16023 = v_16024 & 1'h1;
  assign v_16024 = v_16025 | 1'h0;
  assign v_16025 = ~v_15148;
  assign v_16026 = mux_16026(v_16027);
  assign v_16027 = ~v_16022;
  assign v_16028 = ~v_15155;
  assign v_16029 = v_16030 | v_16031;
  assign v_16030 = mux_16030(v_15157);
  assign v_16031 = mux_16031(v_16016);
  assign v_16033 = v_16034 | v_16893;
  assign v_16034 = act_16035 & 1'h1;
  assign act_16035 = v_16036 | v_16458;
  assign v_16036 = v_16037 & v_16459;
  assign v_16037 = v_16038 & v_16468;
  assign v_16038 = ~v_16039;
  assign v_16040 = v_16041 | v_16452;
  assign v_16041 = act_16042 & 1'h1;
  assign act_16042 = v_16043 | v_16241;
  assign v_16043 = v_16044 & v_16242;
  assign v_16044 = v_16045 & v_16251;
  assign v_16045 = ~v_16046;
  assign v_16047 = v_16048 | v_16235;
  assign v_16048 = act_16049 & 1'h1;
  assign act_16049 = v_16050 | v_16136;
  assign v_16050 = v_16051 & v_16137;
  assign v_16051 = v_16052 & v_16146;
  assign v_16052 = ~v_16053;
  assign v_16054 = v_16055 | v_16130;
  assign v_16055 = act_16056 & 1'h1;
  assign act_16056 = v_16057 | v_16087;
  assign v_16057 = v_16058 & v_16088;
  assign v_16058 = v_16059 & v_16097;
  assign v_16059 = ~v_16060;
  assign v_16061 = v_16062 | v_16081;
  assign v_16062 = act_16063 & 1'h1;
  assign act_16063 = v_16064 | v_16070;
  assign v_16064 = v_16065 & v_16071;
  assign v_16065 = v_16066 & vout_canPeek_16076;
  assign v_16066 = ~vout_canPeek_16067;
  pebbles_core
    pebbles_core_16067
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16068),
       .in0_consume_en(vin0_consume_en_16067),
       .out_canPeek(vout_canPeek_16067),
       .out_peek(vout_peek_16067));
  assign v_16068 = v_16069 | v_16074;
  assign v_16069 = mux_16069(v_16070);
  assign v_16070 = vout_canPeek_16067 & v_16071;
  assign v_16071 = v_16072 & 1'h1;
  assign v_16072 = v_16073 | 1'h0;
  assign v_16073 = ~v_16060;
  assign v_16074 = mux_16074(v_16075);
  assign v_16075 = ~v_16070;
  pebbles_core
    pebbles_core_16076
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16077),
       .in0_consume_en(vin0_consume_en_16076),
       .out_canPeek(vout_canPeek_16076),
       .out_peek(vout_peek_16076));
  assign v_16077 = v_16078 | v_16079;
  assign v_16078 = mux_16078(v_16064);
  assign v_16079 = mux_16079(v_16080);
  assign v_16080 = ~v_16064;
  assign v_16081 = v_16082 & 1'h1;
  assign v_16082 = v_16083 & v_16084;
  assign v_16083 = ~act_16063;
  assign v_16084 = v_16085 | v_16093;
  assign v_16085 = v_16086 | v_16091;
  assign v_16086 = mux_16086(v_16087);
  assign v_16087 = v_16060 & v_16088;
  assign v_16088 = v_16089 & 1'h1;
  assign v_16089 = v_16090 | 1'h0;
  assign v_16090 = ~v_16053;
  assign v_16091 = mux_16091(v_16092);
  assign v_16092 = ~v_16087;
  assign v_16093 = ~v_16060;
  assign v_16094 = v_16095 | v_16096;
  assign v_16095 = mux_16095(v_16062);
  assign v_16096 = mux_16096(v_16081);
  assign v_16098 = v_16099 | v_16118;
  assign v_16099 = act_16100 & 1'h1;
  assign act_16100 = v_16101 | v_16107;
  assign v_16101 = v_16102 & v_16108;
  assign v_16102 = v_16103 & vout_canPeek_16113;
  assign v_16103 = ~vout_canPeek_16104;
  pebbles_core
    pebbles_core_16104
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16105),
       .in0_consume_en(vin0_consume_en_16104),
       .out_canPeek(vout_canPeek_16104),
       .out_peek(vout_peek_16104));
  assign v_16105 = v_16106 | v_16111;
  assign v_16106 = mux_16106(v_16107);
  assign v_16107 = vout_canPeek_16104 & v_16108;
  assign v_16108 = v_16109 & 1'h1;
  assign v_16109 = v_16110 | 1'h0;
  assign v_16110 = ~v_16097;
  assign v_16111 = mux_16111(v_16112);
  assign v_16112 = ~v_16107;
  pebbles_core
    pebbles_core_16113
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16114),
       .in0_consume_en(vin0_consume_en_16113),
       .out_canPeek(vout_canPeek_16113),
       .out_peek(vout_peek_16113));
  assign v_16114 = v_16115 | v_16116;
  assign v_16115 = mux_16115(v_16101);
  assign v_16116 = mux_16116(v_16117);
  assign v_16117 = ~v_16101;
  assign v_16118 = v_16119 & 1'h1;
  assign v_16119 = v_16120 & v_16121;
  assign v_16120 = ~act_16100;
  assign v_16121 = v_16122 | v_16126;
  assign v_16122 = v_16123 | v_16124;
  assign v_16123 = mux_16123(v_16057);
  assign v_16124 = mux_16124(v_16125);
  assign v_16125 = ~v_16057;
  assign v_16126 = ~v_16097;
  assign v_16127 = v_16128 | v_16129;
  assign v_16128 = mux_16128(v_16099);
  assign v_16129 = mux_16129(v_16118);
  assign v_16130 = v_16131 & 1'h1;
  assign v_16131 = v_16132 & v_16133;
  assign v_16132 = ~act_16056;
  assign v_16133 = v_16134 | v_16142;
  assign v_16134 = v_16135 | v_16140;
  assign v_16135 = mux_16135(v_16136);
  assign v_16136 = v_16053 & v_16137;
  assign v_16137 = v_16138 & 1'h1;
  assign v_16138 = v_16139 | 1'h0;
  assign v_16139 = ~v_16046;
  assign v_16140 = mux_16140(v_16141);
  assign v_16141 = ~v_16136;
  assign v_16142 = ~v_16053;
  assign v_16143 = v_16144 | v_16145;
  assign v_16144 = mux_16144(v_16055);
  assign v_16145 = mux_16145(v_16130);
  assign v_16147 = v_16148 | v_16223;
  assign v_16148 = act_16149 & 1'h1;
  assign act_16149 = v_16150 | v_16180;
  assign v_16150 = v_16151 & v_16181;
  assign v_16151 = v_16152 & v_16190;
  assign v_16152 = ~v_16153;
  assign v_16154 = v_16155 | v_16174;
  assign v_16155 = act_16156 & 1'h1;
  assign act_16156 = v_16157 | v_16163;
  assign v_16157 = v_16158 & v_16164;
  assign v_16158 = v_16159 & vout_canPeek_16169;
  assign v_16159 = ~vout_canPeek_16160;
  pebbles_core
    pebbles_core_16160
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16161),
       .in0_consume_en(vin0_consume_en_16160),
       .out_canPeek(vout_canPeek_16160),
       .out_peek(vout_peek_16160));
  assign v_16161 = v_16162 | v_16167;
  assign v_16162 = mux_16162(v_16163);
  assign v_16163 = vout_canPeek_16160 & v_16164;
  assign v_16164 = v_16165 & 1'h1;
  assign v_16165 = v_16166 | 1'h0;
  assign v_16166 = ~v_16153;
  assign v_16167 = mux_16167(v_16168);
  assign v_16168 = ~v_16163;
  pebbles_core
    pebbles_core_16169
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16170),
       .in0_consume_en(vin0_consume_en_16169),
       .out_canPeek(vout_canPeek_16169),
       .out_peek(vout_peek_16169));
  assign v_16170 = v_16171 | v_16172;
  assign v_16171 = mux_16171(v_16157);
  assign v_16172 = mux_16172(v_16173);
  assign v_16173 = ~v_16157;
  assign v_16174 = v_16175 & 1'h1;
  assign v_16175 = v_16176 & v_16177;
  assign v_16176 = ~act_16156;
  assign v_16177 = v_16178 | v_16186;
  assign v_16178 = v_16179 | v_16184;
  assign v_16179 = mux_16179(v_16180);
  assign v_16180 = v_16153 & v_16181;
  assign v_16181 = v_16182 & 1'h1;
  assign v_16182 = v_16183 | 1'h0;
  assign v_16183 = ~v_16146;
  assign v_16184 = mux_16184(v_16185);
  assign v_16185 = ~v_16180;
  assign v_16186 = ~v_16153;
  assign v_16187 = v_16188 | v_16189;
  assign v_16188 = mux_16188(v_16155);
  assign v_16189 = mux_16189(v_16174);
  assign v_16191 = v_16192 | v_16211;
  assign v_16192 = act_16193 & 1'h1;
  assign act_16193 = v_16194 | v_16200;
  assign v_16194 = v_16195 & v_16201;
  assign v_16195 = v_16196 & vout_canPeek_16206;
  assign v_16196 = ~vout_canPeek_16197;
  pebbles_core
    pebbles_core_16197
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16198),
       .in0_consume_en(vin0_consume_en_16197),
       .out_canPeek(vout_canPeek_16197),
       .out_peek(vout_peek_16197));
  assign v_16198 = v_16199 | v_16204;
  assign v_16199 = mux_16199(v_16200);
  assign v_16200 = vout_canPeek_16197 & v_16201;
  assign v_16201 = v_16202 & 1'h1;
  assign v_16202 = v_16203 | 1'h0;
  assign v_16203 = ~v_16190;
  assign v_16204 = mux_16204(v_16205);
  assign v_16205 = ~v_16200;
  pebbles_core
    pebbles_core_16206
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16207),
       .in0_consume_en(vin0_consume_en_16206),
       .out_canPeek(vout_canPeek_16206),
       .out_peek(vout_peek_16206));
  assign v_16207 = v_16208 | v_16209;
  assign v_16208 = mux_16208(v_16194);
  assign v_16209 = mux_16209(v_16210);
  assign v_16210 = ~v_16194;
  assign v_16211 = v_16212 & 1'h1;
  assign v_16212 = v_16213 & v_16214;
  assign v_16213 = ~act_16193;
  assign v_16214 = v_16215 | v_16219;
  assign v_16215 = v_16216 | v_16217;
  assign v_16216 = mux_16216(v_16150);
  assign v_16217 = mux_16217(v_16218);
  assign v_16218 = ~v_16150;
  assign v_16219 = ~v_16190;
  assign v_16220 = v_16221 | v_16222;
  assign v_16221 = mux_16221(v_16192);
  assign v_16222 = mux_16222(v_16211);
  assign v_16223 = v_16224 & 1'h1;
  assign v_16224 = v_16225 & v_16226;
  assign v_16225 = ~act_16149;
  assign v_16226 = v_16227 | v_16231;
  assign v_16227 = v_16228 | v_16229;
  assign v_16228 = mux_16228(v_16050);
  assign v_16229 = mux_16229(v_16230);
  assign v_16230 = ~v_16050;
  assign v_16231 = ~v_16146;
  assign v_16232 = v_16233 | v_16234;
  assign v_16233 = mux_16233(v_16148);
  assign v_16234 = mux_16234(v_16223);
  assign v_16235 = v_16236 & 1'h1;
  assign v_16236 = v_16237 & v_16238;
  assign v_16237 = ~act_16049;
  assign v_16238 = v_16239 | v_16247;
  assign v_16239 = v_16240 | v_16245;
  assign v_16240 = mux_16240(v_16241);
  assign v_16241 = v_16046 & v_16242;
  assign v_16242 = v_16243 & 1'h1;
  assign v_16243 = v_16244 | 1'h0;
  assign v_16244 = ~v_16039;
  assign v_16245 = mux_16245(v_16246);
  assign v_16246 = ~v_16241;
  assign v_16247 = ~v_16046;
  assign v_16248 = v_16249 | v_16250;
  assign v_16249 = mux_16249(v_16048);
  assign v_16250 = mux_16250(v_16235);
  assign v_16252 = v_16253 | v_16440;
  assign v_16253 = act_16254 & 1'h1;
  assign act_16254 = v_16255 | v_16341;
  assign v_16255 = v_16256 & v_16342;
  assign v_16256 = v_16257 & v_16351;
  assign v_16257 = ~v_16258;
  assign v_16259 = v_16260 | v_16335;
  assign v_16260 = act_16261 & 1'h1;
  assign act_16261 = v_16262 | v_16292;
  assign v_16262 = v_16263 & v_16293;
  assign v_16263 = v_16264 & v_16302;
  assign v_16264 = ~v_16265;
  assign v_16266 = v_16267 | v_16286;
  assign v_16267 = act_16268 & 1'h1;
  assign act_16268 = v_16269 | v_16275;
  assign v_16269 = v_16270 & v_16276;
  assign v_16270 = v_16271 & vout_canPeek_16281;
  assign v_16271 = ~vout_canPeek_16272;
  pebbles_core
    pebbles_core_16272
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16273),
       .in0_consume_en(vin0_consume_en_16272),
       .out_canPeek(vout_canPeek_16272),
       .out_peek(vout_peek_16272));
  assign v_16273 = v_16274 | v_16279;
  assign v_16274 = mux_16274(v_16275);
  assign v_16275 = vout_canPeek_16272 & v_16276;
  assign v_16276 = v_16277 & 1'h1;
  assign v_16277 = v_16278 | 1'h0;
  assign v_16278 = ~v_16265;
  assign v_16279 = mux_16279(v_16280);
  assign v_16280 = ~v_16275;
  pebbles_core
    pebbles_core_16281
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16282),
       .in0_consume_en(vin0_consume_en_16281),
       .out_canPeek(vout_canPeek_16281),
       .out_peek(vout_peek_16281));
  assign v_16282 = v_16283 | v_16284;
  assign v_16283 = mux_16283(v_16269);
  assign v_16284 = mux_16284(v_16285);
  assign v_16285 = ~v_16269;
  assign v_16286 = v_16287 & 1'h1;
  assign v_16287 = v_16288 & v_16289;
  assign v_16288 = ~act_16268;
  assign v_16289 = v_16290 | v_16298;
  assign v_16290 = v_16291 | v_16296;
  assign v_16291 = mux_16291(v_16292);
  assign v_16292 = v_16265 & v_16293;
  assign v_16293 = v_16294 & 1'h1;
  assign v_16294 = v_16295 | 1'h0;
  assign v_16295 = ~v_16258;
  assign v_16296 = mux_16296(v_16297);
  assign v_16297 = ~v_16292;
  assign v_16298 = ~v_16265;
  assign v_16299 = v_16300 | v_16301;
  assign v_16300 = mux_16300(v_16267);
  assign v_16301 = mux_16301(v_16286);
  assign v_16303 = v_16304 | v_16323;
  assign v_16304 = act_16305 & 1'h1;
  assign act_16305 = v_16306 | v_16312;
  assign v_16306 = v_16307 & v_16313;
  assign v_16307 = v_16308 & vout_canPeek_16318;
  assign v_16308 = ~vout_canPeek_16309;
  pebbles_core
    pebbles_core_16309
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16310),
       .in0_consume_en(vin0_consume_en_16309),
       .out_canPeek(vout_canPeek_16309),
       .out_peek(vout_peek_16309));
  assign v_16310 = v_16311 | v_16316;
  assign v_16311 = mux_16311(v_16312);
  assign v_16312 = vout_canPeek_16309 & v_16313;
  assign v_16313 = v_16314 & 1'h1;
  assign v_16314 = v_16315 | 1'h0;
  assign v_16315 = ~v_16302;
  assign v_16316 = mux_16316(v_16317);
  assign v_16317 = ~v_16312;
  pebbles_core
    pebbles_core_16318
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16319),
       .in0_consume_en(vin0_consume_en_16318),
       .out_canPeek(vout_canPeek_16318),
       .out_peek(vout_peek_16318));
  assign v_16319 = v_16320 | v_16321;
  assign v_16320 = mux_16320(v_16306);
  assign v_16321 = mux_16321(v_16322);
  assign v_16322 = ~v_16306;
  assign v_16323 = v_16324 & 1'h1;
  assign v_16324 = v_16325 & v_16326;
  assign v_16325 = ~act_16305;
  assign v_16326 = v_16327 | v_16331;
  assign v_16327 = v_16328 | v_16329;
  assign v_16328 = mux_16328(v_16262);
  assign v_16329 = mux_16329(v_16330);
  assign v_16330 = ~v_16262;
  assign v_16331 = ~v_16302;
  assign v_16332 = v_16333 | v_16334;
  assign v_16333 = mux_16333(v_16304);
  assign v_16334 = mux_16334(v_16323);
  assign v_16335 = v_16336 & 1'h1;
  assign v_16336 = v_16337 & v_16338;
  assign v_16337 = ~act_16261;
  assign v_16338 = v_16339 | v_16347;
  assign v_16339 = v_16340 | v_16345;
  assign v_16340 = mux_16340(v_16341);
  assign v_16341 = v_16258 & v_16342;
  assign v_16342 = v_16343 & 1'h1;
  assign v_16343 = v_16344 | 1'h0;
  assign v_16344 = ~v_16251;
  assign v_16345 = mux_16345(v_16346);
  assign v_16346 = ~v_16341;
  assign v_16347 = ~v_16258;
  assign v_16348 = v_16349 | v_16350;
  assign v_16349 = mux_16349(v_16260);
  assign v_16350 = mux_16350(v_16335);
  assign v_16352 = v_16353 | v_16428;
  assign v_16353 = act_16354 & 1'h1;
  assign act_16354 = v_16355 | v_16385;
  assign v_16355 = v_16356 & v_16386;
  assign v_16356 = v_16357 & v_16395;
  assign v_16357 = ~v_16358;
  assign v_16359 = v_16360 | v_16379;
  assign v_16360 = act_16361 & 1'h1;
  assign act_16361 = v_16362 | v_16368;
  assign v_16362 = v_16363 & v_16369;
  assign v_16363 = v_16364 & vout_canPeek_16374;
  assign v_16364 = ~vout_canPeek_16365;
  pebbles_core
    pebbles_core_16365
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16366),
       .in0_consume_en(vin0_consume_en_16365),
       .out_canPeek(vout_canPeek_16365),
       .out_peek(vout_peek_16365));
  assign v_16366 = v_16367 | v_16372;
  assign v_16367 = mux_16367(v_16368);
  assign v_16368 = vout_canPeek_16365 & v_16369;
  assign v_16369 = v_16370 & 1'h1;
  assign v_16370 = v_16371 | 1'h0;
  assign v_16371 = ~v_16358;
  assign v_16372 = mux_16372(v_16373);
  assign v_16373 = ~v_16368;
  pebbles_core
    pebbles_core_16374
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16375),
       .in0_consume_en(vin0_consume_en_16374),
       .out_canPeek(vout_canPeek_16374),
       .out_peek(vout_peek_16374));
  assign v_16375 = v_16376 | v_16377;
  assign v_16376 = mux_16376(v_16362);
  assign v_16377 = mux_16377(v_16378);
  assign v_16378 = ~v_16362;
  assign v_16379 = v_16380 & 1'h1;
  assign v_16380 = v_16381 & v_16382;
  assign v_16381 = ~act_16361;
  assign v_16382 = v_16383 | v_16391;
  assign v_16383 = v_16384 | v_16389;
  assign v_16384 = mux_16384(v_16385);
  assign v_16385 = v_16358 & v_16386;
  assign v_16386 = v_16387 & 1'h1;
  assign v_16387 = v_16388 | 1'h0;
  assign v_16388 = ~v_16351;
  assign v_16389 = mux_16389(v_16390);
  assign v_16390 = ~v_16385;
  assign v_16391 = ~v_16358;
  assign v_16392 = v_16393 | v_16394;
  assign v_16393 = mux_16393(v_16360);
  assign v_16394 = mux_16394(v_16379);
  assign v_16396 = v_16397 | v_16416;
  assign v_16397 = act_16398 & 1'h1;
  assign act_16398 = v_16399 | v_16405;
  assign v_16399 = v_16400 & v_16406;
  assign v_16400 = v_16401 & vout_canPeek_16411;
  assign v_16401 = ~vout_canPeek_16402;
  pebbles_core
    pebbles_core_16402
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16403),
       .in0_consume_en(vin0_consume_en_16402),
       .out_canPeek(vout_canPeek_16402),
       .out_peek(vout_peek_16402));
  assign v_16403 = v_16404 | v_16409;
  assign v_16404 = mux_16404(v_16405);
  assign v_16405 = vout_canPeek_16402 & v_16406;
  assign v_16406 = v_16407 & 1'h1;
  assign v_16407 = v_16408 | 1'h0;
  assign v_16408 = ~v_16395;
  assign v_16409 = mux_16409(v_16410);
  assign v_16410 = ~v_16405;
  pebbles_core
    pebbles_core_16411
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16412),
       .in0_consume_en(vin0_consume_en_16411),
       .out_canPeek(vout_canPeek_16411),
       .out_peek(vout_peek_16411));
  assign v_16412 = v_16413 | v_16414;
  assign v_16413 = mux_16413(v_16399);
  assign v_16414 = mux_16414(v_16415);
  assign v_16415 = ~v_16399;
  assign v_16416 = v_16417 & 1'h1;
  assign v_16417 = v_16418 & v_16419;
  assign v_16418 = ~act_16398;
  assign v_16419 = v_16420 | v_16424;
  assign v_16420 = v_16421 | v_16422;
  assign v_16421 = mux_16421(v_16355);
  assign v_16422 = mux_16422(v_16423);
  assign v_16423 = ~v_16355;
  assign v_16424 = ~v_16395;
  assign v_16425 = v_16426 | v_16427;
  assign v_16426 = mux_16426(v_16397);
  assign v_16427 = mux_16427(v_16416);
  assign v_16428 = v_16429 & 1'h1;
  assign v_16429 = v_16430 & v_16431;
  assign v_16430 = ~act_16354;
  assign v_16431 = v_16432 | v_16436;
  assign v_16432 = v_16433 | v_16434;
  assign v_16433 = mux_16433(v_16255);
  assign v_16434 = mux_16434(v_16435);
  assign v_16435 = ~v_16255;
  assign v_16436 = ~v_16351;
  assign v_16437 = v_16438 | v_16439;
  assign v_16438 = mux_16438(v_16353);
  assign v_16439 = mux_16439(v_16428);
  assign v_16440 = v_16441 & 1'h1;
  assign v_16441 = v_16442 & v_16443;
  assign v_16442 = ~act_16254;
  assign v_16443 = v_16444 | v_16448;
  assign v_16444 = v_16445 | v_16446;
  assign v_16445 = mux_16445(v_16043);
  assign v_16446 = mux_16446(v_16447);
  assign v_16447 = ~v_16043;
  assign v_16448 = ~v_16251;
  assign v_16449 = v_16450 | v_16451;
  assign v_16450 = mux_16450(v_16253);
  assign v_16451 = mux_16451(v_16440);
  assign v_16452 = v_16453 & 1'h1;
  assign v_16453 = v_16454 & v_16455;
  assign v_16454 = ~act_16042;
  assign v_16455 = v_16456 | v_16464;
  assign v_16456 = v_16457 | v_16462;
  assign v_16457 = mux_16457(v_16458);
  assign v_16458 = v_16039 & v_16459;
  assign v_16459 = v_16460 & 1'h1;
  assign v_16460 = v_16461 | 1'h0;
  assign v_16461 = ~v_16032;
  assign v_16462 = mux_16462(v_16463);
  assign v_16463 = ~v_16458;
  assign v_16464 = ~v_16039;
  assign v_16465 = v_16466 | v_16467;
  assign v_16466 = mux_16466(v_16041);
  assign v_16467 = mux_16467(v_16452);
  assign v_16469 = v_16470 | v_16881;
  assign v_16470 = act_16471 & 1'h1;
  assign act_16471 = v_16472 | v_16670;
  assign v_16472 = v_16473 & v_16671;
  assign v_16473 = v_16474 & v_16680;
  assign v_16474 = ~v_16475;
  assign v_16476 = v_16477 | v_16664;
  assign v_16477 = act_16478 & 1'h1;
  assign act_16478 = v_16479 | v_16565;
  assign v_16479 = v_16480 & v_16566;
  assign v_16480 = v_16481 & v_16575;
  assign v_16481 = ~v_16482;
  assign v_16483 = v_16484 | v_16559;
  assign v_16484 = act_16485 & 1'h1;
  assign act_16485 = v_16486 | v_16516;
  assign v_16486 = v_16487 & v_16517;
  assign v_16487 = v_16488 & v_16526;
  assign v_16488 = ~v_16489;
  assign v_16490 = v_16491 | v_16510;
  assign v_16491 = act_16492 & 1'h1;
  assign act_16492 = v_16493 | v_16499;
  assign v_16493 = v_16494 & v_16500;
  assign v_16494 = v_16495 & vout_canPeek_16505;
  assign v_16495 = ~vout_canPeek_16496;
  pebbles_core
    pebbles_core_16496
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16497),
       .in0_consume_en(vin0_consume_en_16496),
       .out_canPeek(vout_canPeek_16496),
       .out_peek(vout_peek_16496));
  assign v_16497 = v_16498 | v_16503;
  assign v_16498 = mux_16498(v_16499);
  assign v_16499 = vout_canPeek_16496 & v_16500;
  assign v_16500 = v_16501 & 1'h1;
  assign v_16501 = v_16502 | 1'h0;
  assign v_16502 = ~v_16489;
  assign v_16503 = mux_16503(v_16504);
  assign v_16504 = ~v_16499;
  pebbles_core
    pebbles_core_16505
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16506),
       .in0_consume_en(vin0_consume_en_16505),
       .out_canPeek(vout_canPeek_16505),
       .out_peek(vout_peek_16505));
  assign v_16506 = v_16507 | v_16508;
  assign v_16507 = mux_16507(v_16493);
  assign v_16508 = mux_16508(v_16509);
  assign v_16509 = ~v_16493;
  assign v_16510 = v_16511 & 1'h1;
  assign v_16511 = v_16512 & v_16513;
  assign v_16512 = ~act_16492;
  assign v_16513 = v_16514 | v_16522;
  assign v_16514 = v_16515 | v_16520;
  assign v_16515 = mux_16515(v_16516);
  assign v_16516 = v_16489 & v_16517;
  assign v_16517 = v_16518 & 1'h1;
  assign v_16518 = v_16519 | 1'h0;
  assign v_16519 = ~v_16482;
  assign v_16520 = mux_16520(v_16521);
  assign v_16521 = ~v_16516;
  assign v_16522 = ~v_16489;
  assign v_16523 = v_16524 | v_16525;
  assign v_16524 = mux_16524(v_16491);
  assign v_16525 = mux_16525(v_16510);
  assign v_16527 = v_16528 | v_16547;
  assign v_16528 = act_16529 & 1'h1;
  assign act_16529 = v_16530 | v_16536;
  assign v_16530 = v_16531 & v_16537;
  assign v_16531 = v_16532 & vout_canPeek_16542;
  assign v_16532 = ~vout_canPeek_16533;
  pebbles_core
    pebbles_core_16533
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16534),
       .in0_consume_en(vin0_consume_en_16533),
       .out_canPeek(vout_canPeek_16533),
       .out_peek(vout_peek_16533));
  assign v_16534 = v_16535 | v_16540;
  assign v_16535 = mux_16535(v_16536);
  assign v_16536 = vout_canPeek_16533 & v_16537;
  assign v_16537 = v_16538 & 1'h1;
  assign v_16538 = v_16539 | 1'h0;
  assign v_16539 = ~v_16526;
  assign v_16540 = mux_16540(v_16541);
  assign v_16541 = ~v_16536;
  pebbles_core
    pebbles_core_16542
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16543),
       .in0_consume_en(vin0_consume_en_16542),
       .out_canPeek(vout_canPeek_16542),
       .out_peek(vout_peek_16542));
  assign v_16543 = v_16544 | v_16545;
  assign v_16544 = mux_16544(v_16530);
  assign v_16545 = mux_16545(v_16546);
  assign v_16546 = ~v_16530;
  assign v_16547 = v_16548 & 1'h1;
  assign v_16548 = v_16549 & v_16550;
  assign v_16549 = ~act_16529;
  assign v_16550 = v_16551 | v_16555;
  assign v_16551 = v_16552 | v_16553;
  assign v_16552 = mux_16552(v_16486);
  assign v_16553 = mux_16553(v_16554);
  assign v_16554 = ~v_16486;
  assign v_16555 = ~v_16526;
  assign v_16556 = v_16557 | v_16558;
  assign v_16557 = mux_16557(v_16528);
  assign v_16558 = mux_16558(v_16547);
  assign v_16559 = v_16560 & 1'h1;
  assign v_16560 = v_16561 & v_16562;
  assign v_16561 = ~act_16485;
  assign v_16562 = v_16563 | v_16571;
  assign v_16563 = v_16564 | v_16569;
  assign v_16564 = mux_16564(v_16565);
  assign v_16565 = v_16482 & v_16566;
  assign v_16566 = v_16567 & 1'h1;
  assign v_16567 = v_16568 | 1'h0;
  assign v_16568 = ~v_16475;
  assign v_16569 = mux_16569(v_16570);
  assign v_16570 = ~v_16565;
  assign v_16571 = ~v_16482;
  assign v_16572 = v_16573 | v_16574;
  assign v_16573 = mux_16573(v_16484);
  assign v_16574 = mux_16574(v_16559);
  assign v_16576 = v_16577 | v_16652;
  assign v_16577 = act_16578 & 1'h1;
  assign act_16578 = v_16579 | v_16609;
  assign v_16579 = v_16580 & v_16610;
  assign v_16580 = v_16581 & v_16619;
  assign v_16581 = ~v_16582;
  assign v_16583 = v_16584 | v_16603;
  assign v_16584 = act_16585 & 1'h1;
  assign act_16585 = v_16586 | v_16592;
  assign v_16586 = v_16587 & v_16593;
  assign v_16587 = v_16588 & vout_canPeek_16598;
  assign v_16588 = ~vout_canPeek_16589;
  pebbles_core
    pebbles_core_16589
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16590),
       .in0_consume_en(vin0_consume_en_16589),
       .out_canPeek(vout_canPeek_16589),
       .out_peek(vout_peek_16589));
  assign v_16590 = v_16591 | v_16596;
  assign v_16591 = mux_16591(v_16592);
  assign v_16592 = vout_canPeek_16589 & v_16593;
  assign v_16593 = v_16594 & 1'h1;
  assign v_16594 = v_16595 | 1'h0;
  assign v_16595 = ~v_16582;
  assign v_16596 = mux_16596(v_16597);
  assign v_16597 = ~v_16592;
  pebbles_core
    pebbles_core_16598
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16599),
       .in0_consume_en(vin0_consume_en_16598),
       .out_canPeek(vout_canPeek_16598),
       .out_peek(vout_peek_16598));
  assign v_16599 = v_16600 | v_16601;
  assign v_16600 = mux_16600(v_16586);
  assign v_16601 = mux_16601(v_16602);
  assign v_16602 = ~v_16586;
  assign v_16603 = v_16604 & 1'h1;
  assign v_16604 = v_16605 & v_16606;
  assign v_16605 = ~act_16585;
  assign v_16606 = v_16607 | v_16615;
  assign v_16607 = v_16608 | v_16613;
  assign v_16608 = mux_16608(v_16609);
  assign v_16609 = v_16582 & v_16610;
  assign v_16610 = v_16611 & 1'h1;
  assign v_16611 = v_16612 | 1'h0;
  assign v_16612 = ~v_16575;
  assign v_16613 = mux_16613(v_16614);
  assign v_16614 = ~v_16609;
  assign v_16615 = ~v_16582;
  assign v_16616 = v_16617 | v_16618;
  assign v_16617 = mux_16617(v_16584);
  assign v_16618 = mux_16618(v_16603);
  assign v_16620 = v_16621 | v_16640;
  assign v_16621 = act_16622 & 1'h1;
  assign act_16622 = v_16623 | v_16629;
  assign v_16623 = v_16624 & v_16630;
  assign v_16624 = v_16625 & vout_canPeek_16635;
  assign v_16625 = ~vout_canPeek_16626;
  pebbles_core
    pebbles_core_16626
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16627),
       .in0_consume_en(vin0_consume_en_16626),
       .out_canPeek(vout_canPeek_16626),
       .out_peek(vout_peek_16626));
  assign v_16627 = v_16628 | v_16633;
  assign v_16628 = mux_16628(v_16629);
  assign v_16629 = vout_canPeek_16626 & v_16630;
  assign v_16630 = v_16631 & 1'h1;
  assign v_16631 = v_16632 | 1'h0;
  assign v_16632 = ~v_16619;
  assign v_16633 = mux_16633(v_16634);
  assign v_16634 = ~v_16629;
  pebbles_core
    pebbles_core_16635
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16636),
       .in0_consume_en(vin0_consume_en_16635),
       .out_canPeek(vout_canPeek_16635),
       .out_peek(vout_peek_16635));
  assign v_16636 = v_16637 | v_16638;
  assign v_16637 = mux_16637(v_16623);
  assign v_16638 = mux_16638(v_16639);
  assign v_16639 = ~v_16623;
  assign v_16640 = v_16641 & 1'h1;
  assign v_16641 = v_16642 & v_16643;
  assign v_16642 = ~act_16622;
  assign v_16643 = v_16644 | v_16648;
  assign v_16644 = v_16645 | v_16646;
  assign v_16645 = mux_16645(v_16579);
  assign v_16646 = mux_16646(v_16647);
  assign v_16647 = ~v_16579;
  assign v_16648 = ~v_16619;
  assign v_16649 = v_16650 | v_16651;
  assign v_16650 = mux_16650(v_16621);
  assign v_16651 = mux_16651(v_16640);
  assign v_16652 = v_16653 & 1'h1;
  assign v_16653 = v_16654 & v_16655;
  assign v_16654 = ~act_16578;
  assign v_16655 = v_16656 | v_16660;
  assign v_16656 = v_16657 | v_16658;
  assign v_16657 = mux_16657(v_16479);
  assign v_16658 = mux_16658(v_16659);
  assign v_16659 = ~v_16479;
  assign v_16660 = ~v_16575;
  assign v_16661 = v_16662 | v_16663;
  assign v_16662 = mux_16662(v_16577);
  assign v_16663 = mux_16663(v_16652);
  assign v_16664 = v_16665 & 1'h1;
  assign v_16665 = v_16666 & v_16667;
  assign v_16666 = ~act_16478;
  assign v_16667 = v_16668 | v_16676;
  assign v_16668 = v_16669 | v_16674;
  assign v_16669 = mux_16669(v_16670);
  assign v_16670 = v_16475 & v_16671;
  assign v_16671 = v_16672 & 1'h1;
  assign v_16672 = v_16673 | 1'h0;
  assign v_16673 = ~v_16468;
  assign v_16674 = mux_16674(v_16675);
  assign v_16675 = ~v_16670;
  assign v_16676 = ~v_16475;
  assign v_16677 = v_16678 | v_16679;
  assign v_16678 = mux_16678(v_16477);
  assign v_16679 = mux_16679(v_16664);
  assign v_16681 = v_16682 | v_16869;
  assign v_16682 = act_16683 & 1'h1;
  assign act_16683 = v_16684 | v_16770;
  assign v_16684 = v_16685 & v_16771;
  assign v_16685 = v_16686 & v_16780;
  assign v_16686 = ~v_16687;
  assign v_16688 = v_16689 | v_16764;
  assign v_16689 = act_16690 & 1'h1;
  assign act_16690 = v_16691 | v_16721;
  assign v_16691 = v_16692 & v_16722;
  assign v_16692 = v_16693 & v_16731;
  assign v_16693 = ~v_16694;
  assign v_16695 = v_16696 | v_16715;
  assign v_16696 = act_16697 & 1'h1;
  assign act_16697 = v_16698 | v_16704;
  assign v_16698 = v_16699 & v_16705;
  assign v_16699 = v_16700 & vout_canPeek_16710;
  assign v_16700 = ~vout_canPeek_16701;
  pebbles_core
    pebbles_core_16701
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16702),
       .in0_consume_en(vin0_consume_en_16701),
       .out_canPeek(vout_canPeek_16701),
       .out_peek(vout_peek_16701));
  assign v_16702 = v_16703 | v_16708;
  assign v_16703 = mux_16703(v_16704);
  assign v_16704 = vout_canPeek_16701 & v_16705;
  assign v_16705 = v_16706 & 1'h1;
  assign v_16706 = v_16707 | 1'h0;
  assign v_16707 = ~v_16694;
  assign v_16708 = mux_16708(v_16709);
  assign v_16709 = ~v_16704;
  pebbles_core
    pebbles_core_16710
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16711),
       .in0_consume_en(vin0_consume_en_16710),
       .out_canPeek(vout_canPeek_16710),
       .out_peek(vout_peek_16710));
  assign v_16711 = v_16712 | v_16713;
  assign v_16712 = mux_16712(v_16698);
  assign v_16713 = mux_16713(v_16714);
  assign v_16714 = ~v_16698;
  assign v_16715 = v_16716 & 1'h1;
  assign v_16716 = v_16717 & v_16718;
  assign v_16717 = ~act_16697;
  assign v_16718 = v_16719 | v_16727;
  assign v_16719 = v_16720 | v_16725;
  assign v_16720 = mux_16720(v_16721);
  assign v_16721 = v_16694 & v_16722;
  assign v_16722 = v_16723 & 1'h1;
  assign v_16723 = v_16724 | 1'h0;
  assign v_16724 = ~v_16687;
  assign v_16725 = mux_16725(v_16726);
  assign v_16726 = ~v_16721;
  assign v_16727 = ~v_16694;
  assign v_16728 = v_16729 | v_16730;
  assign v_16729 = mux_16729(v_16696);
  assign v_16730 = mux_16730(v_16715);
  assign v_16732 = v_16733 | v_16752;
  assign v_16733 = act_16734 & 1'h1;
  assign act_16734 = v_16735 | v_16741;
  assign v_16735 = v_16736 & v_16742;
  assign v_16736 = v_16737 & vout_canPeek_16747;
  assign v_16737 = ~vout_canPeek_16738;
  pebbles_core
    pebbles_core_16738
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16739),
       .in0_consume_en(vin0_consume_en_16738),
       .out_canPeek(vout_canPeek_16738),
       .out_peek(vout_peek_16738));
  assign v_16739 = v_16740 | v_16745;
  assign v_16740 = mux_16740(v_16741);
  assign v_16741 = vout_canPeek_16738 & v_16742;
  assign v_16742 = v_16743 & 1'h1;
  assign v_16743 = v_16744 | 1'h0;
  assign v_16744 = ~v_16731;
  assign v_16745 = mux_16745(v_16746);
  assign v_16746 = ~v_16741;
  pebbles_core
    pebbles_core_16747
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16748),
       .in0_consume_en(vin0_consume_en_16747),
       .out_canPeek(vout_canPeek_16747),
       .out_peek(vout_peek_16747));
  assign v_16748 = v_16749 | v_16750;
  assign v_16749 = mux_16749(v_16735);
  assign v_16750 = mux_16750(v_16751);
  assign v_16751 = ~v_16735;
  assign v_16752 = v_16753 & 1'h1;
  assign v_16753 = v_16754 & v_16755;
  assign v_16754 = ~act_16734;
  assign v_16755 = v_16756 | v_16760;
  assign v_16756 = v_16757 | v_16758;
  assign v_16757 = mux_16757(v_16691);
  assign v_16758 = mux_16758(v_16759);
  assign v_16759 = ~v_16691;
  assign v_16760 = ~v_16731;
  assign v_16761 = v_16762 | v_16763;
  assign v_16762 = mux_16762(v_16733);
  assign v_16763 = mux_16763(v_16752);
  assign v_16764 = v_16765 & 1'h1;
  assign v_16765 = v_16766 & v_16767;
  assign v_16766 = ~act_16690;
  assign v_16767 = v_16768 | v_16776;
  assign v_16768 = v_16769 | v_16774;
  assign v_16769 = mux_16769(v_16770);
  assign v_16770 = v_16687 & v_16771;
  assign v_16771 = v_16772 & 1'h1;
  assign v_16772 = v_16773 | 1'h0;
  assign v_16773 = ~v_16680;
  assign v_16774 = mux_16774(v_16775);
  assign v_16775 = ~v_16770;
  assign v_16776 = ~v_16687;
  assign v_16777 = v_16778 | v_16779;
  assign v_16778 = mux_16778(v_16689);
  assign v_16779 = mux_16779(v_16764);
  assign v_16781 = v_16782 | v_16857;
  assign v_16782 = act_16783 & 1'h1;
  assign act_16783 = v_16784 | v_16814;
  assign v_16784 = v_16785 & v_16815;
  assign v_16785 = v_16786 & v_16824;
  assign v_16786 = ~v_16787;
  assign v_16788 = v_16789 | v_16808;
  assign v_16789 = act_16790 & 1'h1;
  assign act_16790 = v_16791 | v_16797;
  assign v_16791 = v_16792 & v_16798;
  assign v_16792 = v_16793 & vout_canPeek_16803;
  assign v_16793 = ~vout_canPeek_16794;
  pebbles_core
    pebbles_core_16794
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16795),
       .in0_consume_en(vin0_consume_en_16794),
       .out_canPeek(vout_canPeek_16794),
       .out_peek(vout_peek_16794));
  assign v_16795 = v_16796 | v_16801;
  assign v_16796 = mux_16796(v_16797);
  assign v_16797 = vout_canPeek_16794 & v_16798;
  assign v_16798 = v_16799 & 1'h1;
  assign v_16799 = v_16800 | 1'h0;
  assign v_16800 = ~v_16787;
  assign v_16801 = mux_16801(v_16802);
  assign v_16802 = ~v_16797;
  pebbles_core
    pebbles_core_16803
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16804),
       .in0_consume_en(vin0_consume_en_16803),
       .out_canPeek(vout_canPeek_16803),
       .out_peek(vout_peek_16803));
  assign v_16804 = v_16805 | v_16806;
  assign v_16805 = mux_16805(v_16791);
  assign v_16806 = mux_16806(v_16807);
  assign v_16807 = ~v_16791;
  assign v_16808 = v_16809 & 1'h1;
  assign v_16809 = v_16810 & v_16811;
  assign v_16810 = ~act_16790;
  assign v_16811 = v_16812 | v_16820;
  assign v_16812 = v_16813 | v_16818;
  assign v_16813 = mux_16813(v_16814);
  assign v_16814 = v_16787 & v_16815;
  assign v_16815 = v_16816 & 1'h1;
  assign v_16816 = v_16817 | 1'h0;
  assign v_16817 = ~v_16780;
  assign v_16818 = mux_16818(v_16819);
  assign v_16819 = ~v_16814;
  assign v_16820 = ~v_16787;
  assign v_16821 = v_16822 | v_16823;
  assign v_16822 = mux_16822(v_16789);
  assign v_16823 = mux_16823(v_16808);
  assign v_16825 = v_16826 | v_16845;
  assign v_16826 = act_16827 & 1'h1;
  assign act_16827 = v_16828 | v_16834;
  assign v_16828 = v_16829 & v_16835;
  assign v_16829 = v_16830 & vout_canPeek_16840;
  assign v_16830 = ~vout_canPeek_16831;
  pebbles_core
    pebbles_core_16831
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16832),
       .in0_consume_en(vin0_consume_en_16831),
       .out_canPeek(vout_canPeek_16831),
       .out_peek(vout_peek_16831));
  assign v_16832 = v_16833 | v_16838;
  assign v_16833 = mux_16833(v_16834);
  assign v_16834 = vout_canPeek_16831 & v_16835;
  assign v_16835 = v_16836 & 1'h1;
  assign v_16836 = v_16837 | 1'h0;
  assign v_16837 = ~v_16824;
  assign v_16838 = mux_16838(v_16839);
  assign v_16839 = ~v_16834;
  pebbles_core
    pebbles_core_16840
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16841),
       .in0_consume_en(vin0_consume_en_16840),
       .out_canPeek(vout_canPeek_16840),
       .out_peek(vout_peek_16840));
  assign v_16841 = v_16842 | v_16843;
  assign v_16842 = mux_16842(v_16828);
  assign v_16843 = mux_16843(v_16844);
  assign v_16844 = ~v_16828;
  assign v_16845 = v_16846 & 1'h1;
  assign v_16846 = v_16847 & v_16848;
  assign v_16847 = ~act_16827;
  assign v_16848 = v_16849 | v_16853;
  assign v_16849 = v_16850 | v_16851;
  assign v_16850 = mux_16850(v_16784);
  assign v_16851 = mux_16851(v_16852);
  assign v_16852 = ~v_16784;
  assign v_16853 = ~v_16824;
  assign v_16854 = v_16855 | v_16856;
  assign v_16855 = mux_16855(v_16826);
  assign v_16856 = mux_16856(v_16845);
  assign v_16857 = v_16858 & 1'h1;
  assign v_16858 = v_16859 & v_16860;
  assign v_16859 = ~act_16783;
  assign v_16860 = v_16861 | v_16865;
  assign v_16861 = v_16862 | v_16863;
  assign v_16862 = mux_16862(v_16684);
  assign v_16863 = mux_16863(v_16864);
  assign v_16864 = ~v_16684;
  assign v_16865 = ~v_16780;
  assign v_16866 = v_16867 | v_16868;
  assign v_16867 = mux_16867(v_16782);
  assign v_16868 = mux_16868(v_16857);
  assign v_16869 = v_16870 & 1'h1;
  assign v_16870 = v_16871 & v_16872;
  assign v_16871 = ~act_16683;
  assign v_16872 = v_16873 | v_16877;
  assign v_16873 = v_16874 | v_16875;
  assign v_16874 = mux_16874(v_16472);
  assign v_16875 = mux_16875(v_16876);
  assign v_16876 = ~v_16472;
  assign v_16877 = ~v_16680;
  assign v_16878 = v_16879 | v_16880;
  assign v_16879 = mux_16879(v_16682);
  assign v_16880 = mux_16880(v_16869);
  assign v_16881 = v_16882 & 1'h1;
  assign v_16882 = v_16883 & v_16884;
  assign v_16883 = ~act_16471;
  assign v_16884 = v_16885 | v_16889;
  assign v_16885 = v_16886 | v_16887;
  assign v_16886 = mux_16886(v_16036);
  assign v_16887 = mux_16887(v_16888);
  assign v_16888 = ~v_16036;
  assign v_16889 = ~v_16468;
  assign v_16890 = v_16891 | v_16892;
  assign v_16891 = mux_16891(v_16470);
  assign v_16892 = mux_16892(v_16881);
  assign v_16893 = v_16894 & 1'h1;
  assign v_16894 = v_16895 & v_16896;
  assign v_16895 = ~act_16035;
  assign v_16896 = v_16897 | v_16901;
  assign v_16897 = v_16898 | v_16899;
  assign v_16898 = mux_16898(v_15152);
  assign v_16899 = mux_16899(v_16900);
  assign v_16900 = ~v_15152;
  assign v_16901 = ~v_16032;
  assign v_16902 = v_16903 | v_16904;
  assign v_16903 = mux_16903(v_16034);
  assign v_16904 = mux_16904(v_16893);
  assign v_16905 = v_16906 & 1'h1;
  assign v_16906 = v_16907 & v_16908;
  assign v_16907 = ~act_15151;
  assign v_16908 = v_16909 | v_16917;
  assign v_16909 = v_16910 | v_16915;
  assign v_16910 = mux_16910(v_16911);
  assign v_16911 = v_15148 & v_16912;
  assign v_16912 = v_16913 & 1'h1;
  assign v_16913 = v_16914 | 1'h0;
  assign v_16914 = ~v_15141;
  assign v_16915 = mux_16915(v_16916);
  assign v_16916 = ~v_16911;
  assign v_16917 = ~v_15148;
  assign v_16918 = v_16919 | v_16920;
  assign v_16919 = mux_16919(v_15150);
  assign v_16920 = mux_16920(v_16905);
  assign v_16922 = v_16923 | v_18678;
  assign v_16923 = act_16924 & 1'h1;
  assign act_16924 = v_16925 | v_17795;
  assign v_16925 = v_16926 & v_17796;
  assign v_16926 = v_16927 & v_17805;
  assign v_16927 = ~v_16928;
  assign v_16929 = v_16930 | v_17789;
  assign v_16930 = act_16931 & 1'h1;
  assign act_16931 = v_16932 | v_17354;
  assign v_16932 = v_16933 & v_17355;
  assign v_16933 = v_16934 & v_17364;
  assign v_16934 = ~v_16935;
  assign v_16936 = v_16937 | v_17348;
  assign v_16937 = act_16938 & 1'h1;
  assign act_16938 = v_16939 | v_17137;
  assign v_16939 = v_16940 & v_17138;
  assign v_16940 = v_16941 & v_17147;
  assign v_16941 = ~v_16942;
  assign v_16943 = v_16944 | v_17131;
  assign v_16944 = act_16945 & 1'h1;
  assign act_16945 = v_16946 | v_17032;
  assign v_16946 = v_16947 & v_17033;
  assign v_16947 = v_16948 & v_17042;
  assign v_16948 = ~v_16949;
  assign v_16950 = v_16951 | v_17026;
  assign v_16951 = act_16952 & 1'h1;
  assign act_16952 = v_16953 | v_16983;
  assign v_16953 = v_16954 & v_16984;
  assign v_16954 = v_16955 & v_16993;
  assign v_16955 = ~v_16956;
  assign v_16957 = v_16958 | v_16977;
  assign v_16958 = act_16959 & 1'h1;
  assign act_16959 = v_16960 | v_16966;
  assign v_16960 = v_16961 & v_16967;
  assign v_16961 = v_16962 & vout_canPeek_16972;
  assign v_16962 = ~vout_canPeek_16963;
  pebbles_core
    pebbles_core_16963
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16964),
       .in0_consume_en(vin0_consume_en_16963),
       .out_canPeek(vout_canPeek_16963),
       .out_peek(vout_peek_16963));
  assign v_16964 = v_16965 | v_16970;
  assign v_16965 = mux_16965(v_16966);
  assign v_16966 = vout_canPeek_16963 & v_16967;
  assign v_16967 = v_16968 & 1'h1;
  assign v_16968 = v_16969 | 1'h0;
  assign v_16969 = ~v_16956;
  assign v_16970 = mux_16970(v_16971);
  assign v_16971 = ~v_16966;
  pebbles_core
    pebbles_core_16972
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_16973),
       .in0_consume_en(vin0_consume_en_16972),
       .out_canPeek(vout_canPeek_16972),
       .out_peek(vout_peek_16972));
  assign v_16973 = v_16974 | v_16975;
  assign v_16974 = mux_16974(v_16960);
  assign v_16975 = mux_16975(v_16976);
  assign v_16976 = ~v_16960;
  assign v_16977 = v_16978 & 1'h1;
  assign v_16978 = v_16979 & v_16980;
  assign v_16979 = ~act_16959;
  assign v_16980 = v_16981 | v_16989;
  assign v_16981 = v_16982 | v_16987;
  assign v_16982 = mux_16982(v_16983);
  assign v_16983 = v_16956 & v_16984;
  assign v_16984 = v_16985 & 1'h1;
  assign v_16985 = v_16986 | 1'h0;
  assign v_16986 = ~v_16949;
  assign v_16987 = mux_16987(v_16988);
  assign v_16988 = ~v_16983;
  assign v_16989 = ~v_16956;
  assign v_16990 = v_16991 | v_16992;
  assign v_16991 = mux_16991(v_16958);
  assign v_16992 = mux_16992(v_16977);
  assign v_16994 = v_16995 | v_17014;
  assign v_16995 = act_16996 & 1'h1;
  assign act_16996 = v_16997 | v_17003;
  assign v_16997 = v_16998 & v_17004;
  assign v_16998 = v_16999 & vout_canPeek_17009;
  assign v_16999 = ~vout_canPeek_17000;
  pebbles_core
    pebbles_core_17000
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17001),
       .in0_consume_en(vin0_consume_en_17000),
       .out_canPeek(vout_canPeek_17000),
       .out_peek(vout_peek_17000));
  assign v_17001 = v_17002 | v_17007;
  assign v_17002 = mux_17002(v_17003);
  assign v_17003 = vout_canPeek_17000 & v_17004;
  assign v_17004 = v_17005 & 1'h1;
  assign v_17005 = v_17006 | 1'h0;
  assign v_17006 = ~v_16993;
  assign v_17007 = mux_17007(v_17008);
  assign v_17008 = ~v_17003;
  pebbles_core
    pebbles_core_17009
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17010),
       .in0_consume_en(vin0_consume_en_17009),
       .out_canPeek(vout_canPeek_17009),
       .out_peek(vout_peek_17009));
  assign v_17010 = v_17011 | v_17012;
  assign v_17011 = mux_17011(v_16997);
  assign v_17012 = mux_17012(v_17013);
  assign v_17013 = ~v_16997;
  assign v_17014 = v_17015 & 1'h1;
  assign v_17015 = v_17016 & v_17017;
  assign v_17016 = ~act_16996;
  assign v_17017 = v_17018 | v_17022;
  assign v_17018 = v_17019 | v_17020;
  assign v_17019 = mux_17019(v_16953);
  assign v_17020 = mux_17020(v_17021);
  assign v_17021 = ~v_16953;
  assign v_17022 = ~v_16993;
  assign v_17023 = v_17024 | v_17025;
  assign v_17024 = mux_17024(v_16995);
  assign v_17025 = mux_17025(v_17014);
  assign v_17026 = v_17027 & 1'h1;
  assign v_17027 = v_17028 & v_17029;
  assign v_17028 = ~act_16952;
  assign v_17029 = v_17030 | v_17038;
  assign v_17030 = v_17031 | v_17036;
  assign v_17031 = mux_17031(v_17032);
  assign v_17032 = v_16949 & v_17033;
  assign v_17033 = v_17034 & 1'h1;
  assign v_17034 = v_17035 | 1'h0;
  assign v_17035 = ~v_16942;
  assign v_17036 = mux_17036(v_17037);
  assign v_17037 = ~v_17032;
  assign v_17038 = ~v_16949;
  assign v_17039 = v_17040 | v_17041;
  assign v_17040 = mux_17040(v_16951);
  assign v_17041 = mux_17041(v_17026);
  assign v_17043 = v_17044 | v_17119;
  assign v_17044 = act_17045 & 1'h1;
  assign act_17045 = v_17046 | v_17076;
  assign v_17046 = v_17047 & v_17077;
  assign v_17047 = v_17048 & v_17086;
  assign v_17048 = ~v_17049;
  assign v_17050 = v_17051 | v_17070;
  assign v_17051 = act_17052 & 1'h1;
  assign act_17052 = v_17053 | v_17059;
  assign v_17053 = v_17054 & v_17060;
  assign v_17054 = v_17055 & vout_canPeek_17065;
  assign v_17055 = ~vout_canPeek_17056;
  pebbles_core
    pebbles_core_17056
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17057),
       .in0_consume_en(vin0_consume_en_17056),
       .out_canPeek(vout_canPeek_17056),
       .out_peek(vout_peek_17056));
  assign v_17057 = v_17058 | v_17063;
  assign v_17058 = mux_17058(v_17059);
  assign v_17059 = vout_canPeek_17056 & v_17060;
  assign v_17060 = v_17061 & 1'h1;
  assign v_17061 = v_17062 | 1'h0;
  assign v_17062 = ~v_17049;
  assign v_17063 = mux_17063(v_17064);
  assign v_17064 = ~v_17059;
  pebbles_core
    pebbles_core_17065
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17066),
       .in0_consume_en(vin0_consume_en_17065),
       .out_canPeek(vout_canPeek_17065),
       .out_peek(vout_peek_17065));
  assign v_17066 = v_17067 | v_17068;
  assign v_17067 = mux_17067(v_17053);
  assign v_17068 = mux_17068(v_17069);
  assign v_17069 = ~v_17053;
  assign v_17070 = v_17071 & 1'h1;
  assign v_17071 = v_17072 & v_17073;
  assign v_17072 = ~act_17052;
  assign v_17073 = v_17074 | v_17082;
  assign v_17074 = v_17075 | v_17080;
  assign v_17075 = mux_17075(v_17076);
  assign v_17076 = v_17049 & v_17077;
  assign v_17077 = v_17078 & 1'h1;
  assign v_17078 = v_17079 | 1'h0;
  assign v_17079 = ~v_17042;
  assign v_17080 = mux_17080(v_17081);
  assign v_17081 = ~v_17076;
  assign v_17082 = ~v_17049;
  assign v_17083 = v_17084 | v_17085;
  assign v_17084 = mux_17084(v_17051);
  assign v_17085 = mux_17085(v_17070);
  assign v_17087 = v_17088 | v_17107;
  assign v_17088 = act_17089 & 1'h1;
  assign act_17089 = v_17090 | v_17096;
  assign v_17090 = v_17091 & v_17097;
  assign v_17091 = v_17092 & vout_canPeek_17102;
  assign v_17092 = ~vout_canPeek_17093;
  pebbles_core
    pebbles_core_17093
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17094),
       .in0_consume_en(vin0_consume_en_17093),
       .out_canPeek(vout_canPeek_17093),
       .out_peek(vout_peek_17093));
  assign v_17094 = v_17095 | v_17100;
  assign v_17095 = mux_17095(v_17096);
  assign v_17096 = vout_canPeek_17093 & v_17097;
  assign v_17097 = v_17098 & 1'h1;
  assign v_17098 = v_17099 | 1'h0;
  assign v_17099 = ~v_17086;
  assign v_17100 = mux_17100(v_17101);
  assign v_17101 = ~v_17096;
  pebbles_core
    pebbles_core_17102
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17103),
       .in0_consume_en(vin0_consume_en_17102),
       .out_canPeek(vout_canPeek_17102),
       .out_peek(vout_peek_17102));
  assign v_17103 = v_17104 | v_17105;
  assign v_17104 = mux_17104(v_17090);
  assign v_17105 = mux_17105(v_17106);
  assign v_17106 = ~v_17090;
  assign v_17107 = v_17108 & 1'h1;
  assign v_17108 = v_17109 & v_17110;
  assign v_17109 = ~act_17089;
  assign v_17110 = v_17111 | v_17115;
  assign v_17111 = v_17112 | v_17113;
  assign v_17112 = mux_17112(v_17046);
  assign v_17113 = mux_17113(v_17114);
  assign v_17114 = ~v_17046;
  assign v_17115 = ~v_17086;
  assign v_17116 = v_17117 | v_17118;
  assign v_17117 = mux_17117(v_17088);
  assign v_17118 = mux_17118(v_17107);
  assign v_17119 = v_17120 & 1'h1;
  assign v_17120 = v_17121 & v_17122;
  assign v_17121 = ~act_17045;
  assign v_17122 = v_17123 | v_17127;
  assign v_17123 = v_17124 | v_17125;
  assign v_17124 = mux_17124(v_16946);
  assign v_17125 = mux_17125(v_17126);
  assign v_17126 = ~v_16946;
  assign v_17127 = ~v_17042;
  assign v_17128 = v_17129 | v_17130;
  assign v_17129 = mux_17129(v_17044);
  assign v_17130 = mux_17130(v_17119);
  assign v_17131 = v_17132 & 1'h1;
  assign v_17132 = v_17133 & v_17134;
  assign v_17133 = ~act_16945;
  assign v_17134 = v_17135 | v_17143;
  assign v_17135 = v_17136 | v_17141;
  assign v_17136 = mux_17136(v_17137);
  assign v_17137 = v_16942 & v_17138;
  assign v_17138 = v_17139 & 1'h1;
  assign v_17139 = v_17140 | 1'h0;
  assign v_17140 = ~v_16935;
  assign v_17141 = mux_17141(v_17142);
  assign v_17142 = ~v_17137;
  assign v_17143 = ~v_16942;
  assign v_17144 = v_17145 | v_17146;
  assign v_17145 = mux_17145(v_16944);
  assign v_17146 = mux_17146(v_17131);
  assign v_17148 = v_17149 | v_17336;
  assign v_17149 = act_17150 & 1'h1;
  assign act_17150 = v_17151 | v_17237;
  assign v_17151 = v_17152 & v_17238;
  assign v_17152 = v_17153 & v_17247;
  assign v_17153 = ~v_17154;
  assign v_17155 = v_17156 | v_17231;
  assign v_17156 = act_17157 & 1'h1;
  assign act_17157 = v_17158 | v_17188;
  assign v_17158 = v_17159 & v_17189;
  assign v_17159 = v_17160 & v_17198;
  assign v_17160 = ~v_17161;
  assign v_17162 = v_17163 | v_17182;
  assign v_17163 = act_17164 & 1'h1;
  assign act_17164 = v_17165 | v_17171;
  assign v_17165 = v_17166 & v_17172;
  assign v_17166 = v_17167 & vout_canPeek_17177;
  assign v_17167 = ~vout_canPeek_17168;
  pebbles_core
    pebbles_core_17168
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17169),
       .in0_consume_en(vin0_consume_en_17168),
       .out_canPeek(vout_canPeek_17168),
       .out_peek(vout_peek_17168));
  assign v_17169 = v_17170 | v_17175;
  assign v_17170 = mux_17170(v_17171);
  assign v_17171 = vout_canPeek_17168 & v_17172;
  assign v_17172 = v_17173 & 1'h1;
  assign v_17173 = v_17174 | 1'h0;
  assign v_17174 = ~v_17161;
  assign v_17175 = mux_17175(v_17176);
  assign v_17176 = ~v_17171;
  pebbles_core
    pebbles_core_17177
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17178),
       .in0_consume_en(vin0_consume_en_17177),
       .out_canPeek(vout_canPeek_17177),
       .out_peek(vout_peek_17177));
  assign v_17178 = v_17179 | v_17180;
  assign v_17179 = mux_17179(v_17165);
  assign v_17180 = mux_17180(v_17181);
  assign v_17181 = ~v_17165;
  assign v_17182 = v_17183 & 1'h1;
  assign v_17183 = v_17184 & v_17185;
  assign v_17184 = ~act_17164;
  assign v_17185 = v_17186 | v_17194;
  assign v_17186 = v_17187 | v_17192;
  assign v_17187 = mux_17187(v_17188);
  assign v_17188 = v_17161 & v_17189;
  assign v_17189 = v_17190 & 1'h1;
  assign v_17190 = v_17191 | 1'h0;
  assign v_17191 = ~v_17154;
  assign v_17192 = mux_17192(v_17193);
  assign v_17193 = ~v_17188;
  assign v_17194 = ~v_17161;
  assign v_17195 = v_17196 | v_17197;
  assign v_17196 = mux_17196(v_17163);
  assign v_17197 = mux_17197(v_17182);
  assign v_17199 = v_17200 | v_17219;
  assign v_17200 = act_17201 & 1'h1;
  assign act_17201 = v_17202 | v_17208;
  assign v_17202 = v_17203 & v_17209;
  assign v_17203 = v_17204 & vout_canPeek_17214;
  assign v_17204 = ~vout_canPeek_17205;
  pebbles_core
    pebbles_core_17205
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17206),
       .in0_consume_en(vin0_consume_en_17205),
       .out_canPeek(vout_canPeek_17205),
       .out_peek(vout_peek_17205));
  assign v_17206 = v_17207 | v_17212;
  assign v_17207 = mux_17207(v_17208);
  assign v_17208 = vout_canPeek_17205 & v_17209;
  assign v_17209 = v_17210 & 1'h1;
  assign v_17210 = v_17211 | 1'h0;
  assign v_17211 = ~v_17198;
  assign v_17212 = mux_17212(v_17213);
  assign v_17213 = ~v_17208;
  pebbles_core
    pebbles_core_17214
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17215),
       .in0_consume_en(vin0_consume_en_17214),
       .out_canPeek(vout_canPeek_17214),
       .out_peek(vout_peek_17214));
  assign v_17215 = v_17216 | v_17217;
  assign v_17216 = mux_17216(v_17202);
  assign v_17217 = mux_17217(v_17218);
  assign v_17218 = ~v_17202;
  assign v_17219 = v_17220 & 1'h1;
  assign v_17220 = v_17221 & v_17222;
  assign v_17221 = ~act_17201;
  assign v_17222 = v_17223 | v_17227;
  assign v_17223 = v_17224 | v_17225;
  assign v_17224 = mux_17224(v_17158);
  assign v_17225 = mux_17225(v_17226);
  assign v_17226 = ~v_17158;
  assign v_17227 = ~v_17198;
  assign v_17228 = v_17229 | v_17230;
  assign v_17229 = mux_17229(v_17200);
  assign v_17230 = mux_17230(v_17219);
  assign v_17231 = v_17232 & 1'h1;
  assign v_17232 = v_17233 & v_17234;
  assign v_17233 = ~act_17157;
  assign v_17234 = v_17235 | v_17243;
  assign v_17235 = v_17236 | v_17241;
  assign v_17236 = mux_17236(v_17237);
  assign v_17237 = v_17154 & v_17238;
  assign v_17238 = v_17239 & 1'h1;
  assign v_17239 = v_17240 | 1'h0;
  assign v_17240 = ~v_17147;
  assign v_17241 = mux_17241(v_17242);
  assign v_17242 = ~v_17237;
  assign v_17243 = ~v_17154;
  assign v_17244 = v_17245 | v_17246;
  assign v_17245 = mux_17245(v_17156);
  assign v_17246 = mux_17246(v_17231);
  assign v_17248 = v_17249 | v_17324;
  assign v_17249 = act_17250 & 1'h1;
  assign act_17250 = v_17251 | v_17281;
  assign v_17251 = v_17252 & v_17282;
  assign v_17252 = v_17253 & v_17291;
  assign v_17253 = ~v_17254;
  assign v_17255 = v_17256 | v_17275;
  assign v_17256 = act_17257 & 1'h1;
  assign act_17257 = v_17258 | v_17264;
  assign v_17258 = v_17259 & v_17265;
  assign v_17259 = v_17260 & vout_canPeek_17270;
  assign v_17260 = ~vout_canPeek_17261;
  pebbles_core
    pebbles_core_17261
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17262),
       .in0_consume_en(vin0_consume_en_17261),
       .out_canPeek(vout_canPeek_17261),
       .out_peek(vout_peek_17261));
  assign v_17262 = v_17263 | v_17268;
  assign v_17263 = mux_17263(v_17264);
  assign v_17264 = vout_canPeek_17261 & v_17265;
  assign v_17265 = v_17266 & 1'h1;
  assign v_17266 = v_17267 | 1'h0;
  assign v_17267 = ~v_17254;
  assign v_17268 = mux_17268(v_17269);
  assign v_17269 = ~v_17264;
  pebbles_core
    pebbles_core_17270
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17271),
       .in0_consume_en(vin0_consume_en_17270),
       .out_canPeek(vout_canPeek_17270),
       .out_peek(vout_peek_17270));
  assign v_17271 = v_17272 | v_17273;
  assign v_17272 = mux_17272(v_17258);
  assign v_17273 = mux_17273(v_17274);
  assign v_17274 = ~v_17258;
  assign v_17275 = v_17276 & 1'h1;
  assign v_17276 = v_17277 & v_17278;
  assign v_17277 = ~act_17257;
  assign v_17278 = v_17279 | v_17287;
  assign v_17279 = v_17280 | v_17285;
  assign v_17280 = mux_17280(v_17281);
  assign v_17281 = v_17254 & v_17282;
  assign v_17282 = v_17283 & 1'h1;
  assign v_17283 = v_17284 | 1'h0;
  assign v_17284 = ~v_17247;
  assign v_17285 = mux_17285(v_17286);
  assign v_17286 = ~v_17281;
  assign v_17287 = ~v_17254;
  assign v_17288 = v_17289 | v_17290;
  assign v_17289 = mux_17289(v_17256);
  assign v_17290 = mux_17290(v_17275);
  assign v_17292 = v_17293 | v_17312;
  assign v_17293 = act_17294 & 1'h1;
  assign act_17294 = v_17295 | v_17301;
  assign v_17295 = v_17296 & v_17302;
  assign v_17296 = v_17297 & vout_canPeek_17307;
  assign v_17297 = ~vout_canPeek_17298;
  pebbles_core
    pebbles_core_17298
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17299),
       .in0_consume_en(vin0_consume_en_17298),
       .out_canPeek(vout_canPeek_17298),
       .out_peek(vout_peek_17298));
  assign v_17299 = v_17300 | v_17305;
  assign v_17300 = mux_17300(v_17301);
  assign v_17301 = vout_canPeek_17298 & v_17302;
  assign v_17302 = v_17303 & 1'h1;
  assign v_17303 = v_17304 | 1'h0;
  assign v_17304 = ~v_17291;
  assign v_17305 = mux_17305(v_17306);
  assign v_17306 = ~v_17301;
  pebbles_core
    pebbles_core_17307
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17308),
       .in0_consume_en(vin0_consume_en_17307),
       .out_canPeek(vout_canPeek_17307),
       .out_peek(vout_peek_17307));
  assign v_17308 = v_17309 | v_17310;
  assign v_17309 = mux_17309(v_17295);
  assign v_17310 = mux_17310(v_17311);
  assign v_17311 = ~v_17295;
  assign v_17312 = v_17313 & 1'h1;
  assign v_17313 = v_17314 & v_17315;
  assign v_17314 = ~act_17294;
  assign v_17315 = v_17316 | v_17320;
  assign v_17316 = v_17317 | v_17318;
  assign v_17317 = mux_17317(v_17251);
  assign v_17318 = mux_17318(v_17319);
  assign v_17319 = ~v_17251;
  assign v_17320 = ~v_17291;
  assign v_17321 = v_17322 | v_17323;
  assign v_17322 = mux_17322(v_17293);
  assign v_17323 = mux_17323(v_17312);
  assign v_17324 = v_17325 & 1'h1;
  assign v_17325 = v_17326 & v_17327;
  assign v_17326 = ~act_17250;
  assign v_17327 = v_17328 | v_17332;
  assign v_17328 = v_17329 | v_17330;
  assign v_17329 = mux_17329(v_17151);
  assign v_17330 = mux_17330(v_17331);
  assign v_17331 = ~v_17151;
  assign v_17332 = ~v_17247;
  assign v_17333 = v_17334 | v_17335;
  assign v_17334 = mux_17334(v_17249);
  assign v_17335 = mux_17335(v_17324);
  assign v_17336 = v_17337 & 1'h1;
  assign v_17337 = v_17338 & v_17339;
  assign v_17338 = ~act_17150;
  assign v_17339 = v_17340 | v_17344;
  assign v_17340 = v_17341 | v_17342;
  assign v_17341 = mux_17341(v_16939);
  assign v_17342 = mux_17342(v_17343);
  assign v_17343 = ~v_16939;
  assign v_17344 = ~v_17147;
  assign v_17345 = v_17346 | v_17347;
  assign v_17346 = mux_17346(v_17149);
  assign v_17347 = mux_17347(v_17336);
  assign v_17348 = v_17349 & 1'h1;
  assign v_17349 = v_17350 & v_17351;
  assign v_17350 = ~act_16938;
  assign v_17351 = v_17352 | v_17360;
  assign v_17352 = v_17353 | v_17358;
  assign v_17353 = mux_17353(v_17354);
  assign v_17354 = v_16935 & v_17355;
  assign v_17355 = v_17356 & 1'h1;
  assign v_17356 = v_17357 | 1'h0;
  assign v_17357 = ~v_16928;
  assign v_17358 = mux_17358(v_17359);
  assign v_17359 = ~v_17354;
  assign v_17360 = ~v_16935;
  assign v_17361 = v_17362 | v_17363;
  assign v_17362 = mux_17362(v_16937);
  assign v_17363 = mux_17363(v_17348);
  assign v_17365 = v_17366 | v_17777;
  assign v_17366 = act_17367 & 1'h1;
  assign act_17367 = v_17368 | v_17566;
  assign v_17368 = v_17369 & v_17567;
  assign v_17369 = v_17370 & v_17576;
  assign v_17370 = ~v_17371;
  assign v_17372 = v_17373 | v_17560;
  assign v_17373 = act_17374 & 1'h1;
  assign act_17374 = v_17375 | v_17461;
  assign v_17375 = v_17376 & v_17462;
  assign v_17376 = v_17377 & v_17471;
  assign v_17377 = ~v_17378;
  assign v_17379 = v_17380 | v_17455;
  assign v_17380 = act_17381 & 1'h1;
  assign act_17381 = v_17382 | v_17412;
  assign v_17382 = v_17383 & v_17413;
  assign v_17383 = v_17384 & v_17422;
  assign v_17384 = ~v_17385;
  assign v_17386 = v_17387 | v_17406;
  assign v_17387 = act_17388 & 1'h1;
  assign act_17388 = v_17389 | v_17395;
  assign v_17389 = v_17390 & v_17396;
  assign v_17390 = v_17391 & vout_canPeek_17401;
  assign v_17391 = ~vout_canPeek_17392;
  pebbles_core
    pebbles_core_17392
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17393),
       .in0_consume_en(vin0_consume_en_17392),
       .out_canPeek(vout_canPeek_17392),
       .out_peek(vout_peek_17392));
  assign v_17393 = v_17394 | v_17399;
  assign v_17394 = mux_17394(v_17395);
  assign v_17395 = vout_canPeek_17392 & v_17396;
  assign v_17396 = v_17397 & 1'h1;
  assign v_17397 = v_17398 | 1'h0;
  assign v_17398 = ~v_17385;
  assign v_17399 = mux_17399(v_17400);
  assign v_17400 = ~v_17395;
  pebbles_core
    pebbles_core_17401
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17402),
       .in0_consume_en(vin0_consume_en_17401),
       .out_canPeek(vout_canPeek_17401),
       .out_peek(vout_peek_17401));
  assign v_17402 = v_17403 | v_17404;
  assign v_17403 = mux_17403(v_17389);
  assign v_17404 = mux_17404(v_17405);
  assign v_17405 = ~v_17389;
  assign v_17406 = v_17407 & 1'h1;
  assign v_17407 = v_17408 & v_17409;
  assign v_17408 = ~act_17388;
  assign v_17409 = v_17410 | v_17418;
  assign v_17410 = v_17411 | v_17416;
  assign v_17411 = mux_17411(v_17412);
  assign v_17412 = v_17385 & v_17413;
  assign v_17413 = v_17414 & 1'h1;
  assign v_17414 = v_17415 | 1'h0;
  assign v_17415 = ~v_17378;
  assign v_17416 = mux_17416(v_17417);
  assign v_17417 = ~v_17412;
  assign v_17418 = ~v_17385;
  assign v_17419 = v_17420 | v_17421;
  assign v_17420 = mux_17420(v_17387);
  assign v_17421 = mux_17421(v_17406);
  assign v_17423 = v_17424 | v_17443;
  assign v_17424 = act_17425 & 1'h1;
  assign act_17425 = v_17426 | v_17432;
  assign v_17426 = v_17427 & v_17433;
  assign v_17427 = v_17428 & vout_canPeek_17438;
  assign v_17428 = ~vout_canPeek_17429;
  pebbles_core
    pebbles_core_17429
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17430),
       .in0_consume_en(vin0_consume_en_17429),
       .out_canPeek(vout_canPeek_17429),
       .out_peek(vout_peek_17429));
  assign v_17430 = v_17431 | v_17436;
  assign v_17431 = mux_17431(v_17432);
  assign v_17432 = vout_canPeek_17429 & v_17433;
  assign v_17433 = v_17434 & 1'h1;
  assign v_17434 = v_17435 | 1'h0;
  assign v_17435 = ~v_17422;
  assign v_17436 = mux_17436(v_17437);
  assign v_17437 = ~v_17432;
  pebbles_core
    pebbles_core_17438
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17439),
       .in0_consume_en(vin0_consume_en_17438),
       .out_canPeek(vout_canPeek_17438),
       .out_peek(vout_peek_17438));
  assign v_17439 = v_17440 | v_17441;
  assign v_17440 = mux_17440(v_17426);
  assign v_17441 = mux_17441(v_17442);
  assign v_17442 = ~v_17426;
  assign v_17443 = v_17444 & 1'h1;
  assign v_17444 = v_17445 & v_17446;
  assign v_17445 = ~act_17425;
  assign v_17446 = v_17447 | v_17451;
  assign v_17447 = v_17448 | v_17449;
  assign v_17448 = mux_17448(v_17382);
  assign v_17449 = mux_17449(v_17450);
  assign v_17450 = ~v_17382;
  assign v_17451 = ~v_17422;
  assign v_17452 = v_17453 | v_17454;
  assign v_17453 = mux_17453(v_17424);
  assign v_17454 = mux_17454(v_17443);
  assign v_17455 = v_17456 & 1'h1;
  assign v_17456 = v_17457 & v_17458;
  assign v_17457 = ~act_17381;
  assign v_17458 = v_17459 | v_17467;
  assign v_17459 = v_17460 | v_17465;
  assign v_17460 = mux_17460(v_17461);
  assign v_17461 = v_17378 & v_17462;
  assign v_17462 = v_17463 & 1'h1;
  assign v_17463 = v_17464 | 1'h0;
  assign v_17464 = ~v_17371;
  assign v_17465 = mux_17465(v_17466);
  assign v_17466 = ~v_17461;
  assign v_17467 = ~v_17378;
  assign v_17468 = v_17469 | v_17470;
  assign v_17469 = mux_17469(v_17380);
  assign v_17470 = mux_17470(v_17455);
  assign v_17472 = v_17473 | v_17548;
  assign v_17473 = act_17474 & 1'h1;
  assign act_17474 = v_17475 | v_17505;
  assign v_17475 = v_17476 & v_17506;
  assign v_17476 = v_17477 & v_17515;
  assign v_17477 = ~v_17478;
  assign v_17479 = v_17480 | v_17499;
  assign v_17480 = act_17481 & 1'h1;
  assign act_17481 = v_17482 | v_17488;
  assign v_17482 = v_17483 & v_17489;
  assign v_17483 = v_17484 & vout_canPeek_17494;
  assign v_17484 = ~vout_canPeek_17485;
  pebbles_core
    pebbles_core_17485
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17486),
       .in0_consume_en(vin0_consume_en_17485),
       .out_canPeek(vout_canPeek_17485),
       .out_peek(vout_peek_17485));
  assign v_17486 = v_17487 | v_17492;
  assign v_17487 = mux_17487(v_17488);
  assign v_17488 = vout_canPeek_17485 & v_17489;
  assign v_17489 = v_17490 & 1'h1;
  assign v_17490 = v_17491 | 1'h0;
  assign v_17491 = ~v_17478;
  assign v_17492 = mux_17492(v_17493);
  assign v_17493 = ~v_17488;
  pebbles_core
    pebbles_core_17494
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17495),
       .in0_consume_en(vin0_consume_en_17494),
       .out_canPeek(vout_canPeek_17494),
       .out_peek(vout_peek_17494));
  assign v_17495 = v_17496 | v_17497;
  assign v_17496 = mux_17496(v_17482);
  assign v_17497 = mux_17497(v_17498);
  assign v_17498 = ~v_17482;
  assign v_17499 = v_17500 & 1'h1;
  assign v_17500 = v_17501 & v_17502;
  assign v_17501 = ~act_17481;
  assign v_17502 = v_17503 | v_17511;
  assign v_17503 = v_17504 | v_17509;
  assign v_17504 = mux_17504(v_17505);
  assign v_17505 = v_17478 & v_17506;
  assign v_17506 = v_17507 & 1'h1;
  assign v_17507 = v_17508 | 1'h0;
  assign v_17508 = ~v_17471;
  assign v_17509 = mux_17509(v_17510);
  assign v_17510 = ~v_17505;
  assign v_17511 = ~v_17478;
  assign v_17512 = v_17513 | v_17514;
  assign v_17513 = mux_17513(v_17480);
  assign v_17514 = mux_17514(v_17499);
  assign v_17516 = v_17517 | v_17536;
  assign v_17517 = act_17518 & 1'h1;
  assign act_17518 = v_17519 | v_17525;
  assign v_17519 = v_17520 & v_17526;
  assign v_17520 = v_17521 & vout_canPeek_17531;
  assign v_17521 = ~vout_canPeek_17522;
  pebbles_core
    pebbles_core_17522
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17523),
       .in0_consume_en(vin0_consume_en_17522),
       .out_canPeek(vout_canPeek_17522),
       .out_peek(vout_peek_17522));
  assign v_17523 = v_17524 | v_17529;
  assign v_17524 = mux_17524(v_17525);
  assign v_17525 = vout_canPeek_17522 & v_17526;
  assign v_17526 = v_17527 & 1'h1;
  assign v_17527 = v_17528 | 1'h0;
  assign v_17528 = ~v_17515;
  assign v_17529 = mux_17529(v_17530);
  assign v_17530 = ~v_17525;
  pebbles_core
    pebbles_core_17531
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17532),
       .in0_consume_en(vin0_consume_en_17531),
       .out_canPeek(vout_canPeek_17531),
       .out_peek(vout_peek_17531));
  assign v_17532 = v_17533 | v_17534;
  assign v_17533 = mux_17533(v_17519);
  assign v_17534 = mux_17534(v_17535);
  assign v_17535 = ~v_17519;
  assign v_17536 = v_17537 & 1'h1;
  assign v_17537 = v_17538 & v_17539;
  assign v_17538 = ~act_17518;
  assign v_17539 = v_17540 | v_17544;
  assign v_17540 = v_17541 | v_17542;
  assign v_17541 = mux_17541(v_17475);
  assign v_17542 = mux_17542(v_17543);
  assign v_17543 = ~v_17475;
  assign v_17544 = ~v_17515;
  assign v_17545 = v_17546 | v_17547;
  assign v_17546 = mux_17546(v_17517);
  assign v_17547 = mux_17547(v_17536);
  assign v_17548 = v_17549 & 1'h1;
  assign v_17549 = v_17550 & v_17551;
  assign v_17550 = ~act_17474;
  assign v_17551 = v_17552 | v_17556;
  assign v_17552 = v_17553 | v_17554;
  assign v_17553 = mux_17553(v_17375);
  assign v_17554 = mux_17554(v_17555);
  assign v_17555 = ~v_17375;
  assign v_17556 = ~v_17471;
  assign v_17557 = v_17558 | v_17559;
  assign v_17558 = mux_17558(v_17473);
  assign v_17559 = mux_17559(v_17548);
  assign v_17560 = v_17561 & 1'h1;
  assign v_17561 = v_17562 & v_17563;
  assign v_17562 = ~act_17374;
  assign v_17563 = v_17564 | v_17572;
  assign v_17564 = v_17565 | v_17570;
  assign v_17565 = mux_17565(v_17566);
  assign v_17566 = v_17371 & v_17567;
  assign v_17567 = v_17568 & 1'h1;
  assign v_17568 = v_17569 | 1'h0;
  assign v_17569 = ~v_17364;
  assign v_17570 = mux_17570(v_17571);
  assign v_17571 = ~v_17566;
  assign v_17572 = ~v_17371;
  assign v_17573 = v_17574 | v_17575;
  assign v_17574 = mux_17574(v_17373);
  assign v_17575 = mux_17575(v_17560);
  assign v_17577 = v_17578 | v_17765;
  assign v_17578 = act_17579 & 1'h1;
  assign act_17579 = v_17580 | v_17666;
  assign v_17580 = v_17581 & v_17667;
  assign v_17581 = v_17582 & v_17676;
  assign v_17582 = ~v_17583;
  assign v_17584 = v_17585 | v_17660;
  assign v_17585 = act_17586 & 1'h1;
  assign act_17586 = v_17587 | v_17617;
  assign v_17587 = v_17588 & v_17618;
  assign v_17588 = v_17589 & v_17627;
  assign v_17589 = ~v_17590;
  assign v_17591 = v_17592 | v_17611;
  assign v_17592 = act_17593 & 1'h1;
  assign act_17593 = v_17594 | v_17600;
  assign v_17594 = v_17595 & v_17601;
  assign v_17595 = v_17596 & vout_canPeek_17606;
  assign v_17596 = ~vout_canPeek_17597;
  pebbles_core
    pebbles_core_17597
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17598),
       .in0_consume_en(vin0_consume_en_17597),
       .out_canPeek(vout_canPeek_17597),
       .out_peek(vout_peek_17597));
  assign v_17598 = v_17599 | v_17604;
  assign v_17599 = mux_17599(v_17600);
  assign v_17600 = vout_canPeek_17597 & v_17601;
  assign v_17601 = v_17602 & 1'h1;
  assign v_17602 = v_17603 | 1'h0;
  assign v_17603 = ~v_17590;
  assign v_17604 = mux_17604(v_17605);
  assign v_17605 = ~v_17600;
  pebbles_core
    pebbles_core_17606
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17607),
       .in0_consume_en(vin0_consume_en_17606),
       .out_canPeek(vout_canPeek_17606),
       .out_peek(vout_peek_17606));
  assign v_17607 = v_17608 | v_17609;
  assign v_17608 = mux_17608(v_17594);
  assign v_17609 = mux_17609(v_17610);
  assign v_17610 = ~v_17594;
  assign v_17611 = v_17612 & 1'h1;
  assign v_17612 = v_17613 & v_17614;
  assign v_17613 = ~act_17593;
  assign v_17614 = v_17615 | v_17623;
  assign v_17615 = v_17616 | v_17621;
  assign v_17616 = mux_17616(v_17617);
  assign v_17617 = v_17590 & v_17618;
  assign v_17618 = v_17619 & 1'h1;
  assign v_17619 = v_17620 | 1'h0;
  assign v_17620 = ~v_17583;
  assign v_17621 = mux_17621(v_17622);
  assign v_17622 = ~v_17617;
  assign v_17623 = ~v_17590;
  assign v_17624 = v_17625 | v_17626;
  assign v_17625 = mux_17625(v_17592);
  assign v_17626 = mux_17626(v_17611);
  assign v_17628 = v_17629 | v_17648;
  assign v_17629 = act_17630 & 1'h1;
  assign act_17630 = v_17631 | v_17637;
  assign v_17631 = v_17632 & v_17638;
  assign v_17632 = v_17633 & vout_canPeek_17643;
  assign v_17633 = ~vout_canPeek_17634;
  pebbles_core
    pebbles_core_17634
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17635),
       .in0_consume_en(vin0_consume_en_17634),
       .out_canPeek(vout_canPeek_17634),
       .out_peek(vout_peek_17634));
  assign v_17635 = v_17636 | v_17641;
  assign v_17636 = mux_17636(v_17637);
  assign v_17637 = vout_canPeek_17634 & v_17638;
  assign v_17638 = v_17639 & 1'h1;
  assign v_17639 = v_17640 | 1'h0;
  assign v_17640 = ~v_17627;
  assign v_17641 = mux_17641(v_17642);
  assign v_17642 = ~v_17637;
  pebbles_core
    pebbles_core_17643
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17644),
       .in0_consume_en(vin0_consume_en_17643),
       .out_canPeek(vout_canPeek_17643),
       .out_peek(vout_peek_17643));
  assign v_17644 = v_17645 | v_17646;
  assign v_17645 = mux_17645(v_17631);
  assign v_17646 = mux_17646(v_17647);
  assign v_17647 = ~v_17631;
  assign v_17648 = v_17649 & 1'h1;
  assign v_17649 = v_17650 & v_17651;
  assign v_17650 = ~act_17630;
  assign v_17651 = v_17652 | v_17656;
  assign v_17652 = v_17653 | v_17654;
  assign v_17653 = mux_17653(v_17587);
  assign v_17654 = mux_17654(v_17655);
  assign v_17655 = ~v_17587;
  assign v_17656 = ~v_17627;
  assign v_17657 = v_17658 | v_17659;
  assign v_17658 = mux_17658(v_17629);
  assign v_17659 = mux_17659(v_17648);
  assign v_17660 = v_17661 & 1'h1;
  assign v_17661 = v_17662 & v_17663;
  assign v_17662 = ~act_17586;
  assign v_17663 = v_17664 | v_17672;
  assign v_17664 = v_17665 | v_17670;
  assign v_17665 = mux_17665(v_17666);
  assign v_17666 = v_17583 & v_17667;
  assign v_17667 = v_17668 & 1'h1;
  assign v_17668 = v_17669 | 1'h0;
  assign v_17669 = ~v_17576;
  assign v_17670 = mux_17670(v_17671);
  assign v_17671 = ~v_17666;
  assign v_17672 = ~v_17583;
  assign v_17673 = v_17674 | v_17675;
  assign v_17674 = mux_17674(v_17585);
  assign v_17675 = mux_17675(v_17660);
  assign v_17677 = v_17678 | v_17753;
  assign v_17678 = act_17679 & 1'h1;
  assign act_17679 = v_17680 | v_17710;
  assign v_17680 = v_17681 & v_17711;
  assign v_17681 = v_17682 & v_17720;
  assign v_17682 = ~v_17683;
  assign v_17684 = v_17685 | v_17704;
  assign v_17685 = act_17686 & 1'h1;
  assign act_17686 = v_17687 | v_17693;
  assign v_17687 = v_17688 & v_17694;
  assign v_17688 = v_17689 & vout_canPeek_17699;
  assign v_17689 = ~vout_canPeek_17690;
  pebbles_core
    pebbles_core_17690
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17691),
       .in0_consume_en(vin0_consume_en_17690),
       .out_canPeek(vout_canPeek_17690),
       .out_peek(vout_peek_17690));
  assign v_17691 = v_17692 | v_17697;
  assign v_17692 = mux_17692(v_17693);
  assign v_17693 = vout_canPeek_17690 & v_17694;
  assign v_17694 = v_17695 & 1'h1;
  assign v_17695 = v_17696 | 1'h0;
  assign v_17696 = ~v_17683;
  assign v_17697 = mux_17697(v_17698);
  assign v_17698 = ~v_17693;
  pebbles_core
    pebbles_core_17699
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17700),
       .in0_consume_en(vin0_consume_en_17699),
       .out_canPeek(vout_canPeek_17699),
       .out_peek(vout_peek_17699));
  assign v_17700 = v_17701 | v_17702;
  assign v_17701 = mux_17701(v_17687);
  assign v_17702 = mux_17702(v_17703);
  assign v_17703 = ~v_17687;
  assign v_17704 = v_17705 & 1'h1;
  assign v_17705 = v_17706 & v_17707;
  assign v_17706 = ~act_17686;
  assign v_17707 = v_17708 | v_17716;
  assign v_17708 = v_17709 | v_17714;
  assign v_17709 = mux_17709(v_17710);
  assign v_17710 = v_17683 & v_17711;
  assign v_17711 = v_17712 & 1'h1;
  assign v_17712 = v_17713 | 1'h0;
  assign v_17713 = ~v_17676;
  assign v_17714 = mux_17714(v_17715);
  assign v_17715 = ~v_17710;
  assign v_17716 = ~v_17683;
  assign v_17717 = v_17718 | v_17719;
  assign v_17718 = mux_17718(v_17685);
  assign v_17719 = mux_17719(v_17704);
  assign v_17721 = v_17722 | v_17741;
  assign v_17722 = act_17723 & 1'h1;
  assign act_17723 = v_17724 | v_17730;
  assign v_17724 = v_17725 & v_17731;
  assign v_17725 = v_17726 & vout_canPeek_17736;
  assign v_17726 = ~vout_canPeek_17727;
  pebbles_core
    pebbles_core_17727
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17728),
       .in0_consume_en(vin0_consume_en_17727),
       .out_canPeek(vout_canPeek_17727),
       .out_peek(vout_peek_17727));
  assign v_17728 = v_17729 | v_17734;
  assign v_17729 = mux_17729(v_17730);
  assign v_17730 = vout_canPeek_17727 & v_17731;
  assign v_17731 = v_17732 & 1'h1;
  assign v_17732 = v_17733 | 1'h0;
  assign v_17733 = ~v_17720;
  assign v_17734 = mux_17734(v_17735);
  assign v_17735 = ~v_17730;
  pebbles_core
    pebbles_core_17736
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17737),
       .in0_consume_en(vin0_consume_en_17736),
       .out_canPeek(vout_canPeek_17736),
       .out_peek(vout_peek_17736));
  assign v_17737 = v_17738 | v_17739;
  assign v_17738 = mux_17738(v_17724);
  assign v_17739 = mux_17739(v_17740);
  assign v_17740 = ~v_17724;
  assign v_17741 = v_17742 & 1'h1;
  assign v_17742 = v_17743 & v_17744;
  assign v_17743 = ~act_17723;
  assign v_17744 = v_17745 | v_17749;
  assign v_17745 = v_17746 | v_17747;
  assign v_17746 = mux_17746(v_17680);
  assign v_17747 = mux_17747(v_17748);
  assign v_17748 = ~v_17680;
  assign v_17749 = ~v_17720;
  assign v_17750 = v_17751 | v_17752;
  assign v_17751 = mux_17751(v_17722);
  assign v_17752 = mux_17752(v_17741);
  assign v_17753 = v_17754 & 1'h1;
  assign v_17754 = v_17755 & v_17756;
  assign v_17755 = ~act_17679;
  assign v_17756 = v_17757 | v_17761;
  assign v_17757 = v_17758 | v_17759;
  assign v_17758 = mux_17758(v_17580);
  assign v_17759 = mux_17759(v_17760);
  assign v_17760 = ~v_17580;
  assign v_17761 = ~v_17676;
  assign v_17762 = v_17763 | v_17764;
  assign v_17763 = mux_17763(v_17678);
  assign v_17764 = mux_17764(v_17753);
  assign v_17765 = v_17766 & 1'h1;
  assign v_17766 = v_17767 & v_17768;
  assign v_17767 = ~act_17579;
  assign v_17768 = v_17769 | v_17773;
  assign v_17769 = v_17770 | v_17771;
  assign v_17770 = mux_17770(v_17368);
  assign v_17771 = mux_17771(v_17772);
  assign v_17772 = ~v_17368;
  assign v_17773 = ~v_17576;
  assign v_17774 = v_17775 | v_17776;
  assign v_17775 = mux_17775(v_17578);
  assign v_17776 = mux_17776(v_17765);
  assign v_17777 = v_17778 & 1'h1;
  assign v_17778 = v_17779 & v_17780;
  assign v_17779 = ~act_17367;
  assign v_17780 = v_17781 | v_17785;
  assign v_17781 = v_17782 | v_17783;
  assign v_17782 = mux_17782(v_16932);
  assign v_17783 = mux_17783(v_17784);
  assign v_17784 = ~v_16932;
  assign v_17785 = ~v_17364;
  assign v_17786 = v_17787 | v_17788;
  assign v_17787 = mux_17787(v_17366);
  assign v_17788 = mux_17788(v_17777);
  assign v_17789 = v_17790 & 1'h1;
  assign v_17790 = v_17791 & v_17792;
  assign v_17791 = ~act_16931;
  assign v_17792 = v_17793 | v_17801;
  assign v_17793 = v_17794 | v_17799;
  assign v_17794 = mux_17794(v_17795);
  assign v_17795 = v_16928 & v_17796;
  assign v_17796 = v_17797 & 1'h1;
  assign v_17797 = v_17798 | 1'h0;
  assign v_17798 = ~v_16921;
  assign v_17799 = mux_17799(v_17800);
  assign v_17800 = ~v_17795;
  assign v_17801 = ~v_16928;
  assign v_17802 = v_17803 | v_17804;
  assign v_17803 = mux_17803(v_16930);
  assign v_17804 = mux_17804(v_17789);
  assign v_17806 = v_17807 | v_18666;
  assign v_17807 = act_17808 & 1'h1;
  assign act_17808 = v_17809 | v_18231;
  assign v_17809 = v_17810 & v_18232;
  assign v_17810 = v_17811 & v_18241;
  assign v_17811 = ~v_17812;
  assign v_17813 = v_17814 | v_18225;
  assign v_17814 = act_17815 & 1'h1;
  assign act_17815 = v_17816 | v_18014;
  assign v_17816 = v_17817 & v_18015;
  assign v_17817 = v_17818 & v_18024;
  assign v_17818 = ~v_17819;
  assign v_17820 = v_17821 | v_18008;
  assign v_17821 = act_17822 & 1'h1;
  assign act_17822 = v_17823 | v_17909;
  assign v_17823 = v_17824 & v_17910;
  assign v_17824 = v_17825 & v_17919;
  assign v_17825 = ~v_17826;
  assign v_17827 = v_17828 | v_17903;
  assign v_17828 = act_17829 & 1'h1;
  assign act_17829 = v_17830 | v_17860;
  assign v_17830 = v_17831 & v_17861;
  assign v_17831 = v_17832 & v_17870;
  assign v_17832 = ~v_17833;
  assign v_17834 = v_17835 | v_17854;
  assign v_17835 = act_17836 & 1'h1;
  assign act_17836 = v_17837 | v_17843;
  assign v_17837 = v_17838 & v_17844;
  assign v_17838 = v_17839 & vout_canPeek_17849;
  assign v_17839 = ~vout_canPeek_17840;
  pebbles_core
    pebbles_core_17840
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17841),
       .in0_consume_en(vin0_consume_en_17840),
       .out_canPeek(vout_canPeek_17840),
       .out_peek(vout_peek_17840));
  assign v_17841 = v_17842 | v_17847;
  assign v_17842 = mux_17842(v_17843);
  assign v_17843 = vout_canPeek_17840 & v_17844;
  assign v_17844 = v_17845 & 1'h1;
  assign v_17845 = v_17846 | 1'h0;
  assign v_17846 = ~v_17833;
  assign v_17847 = mux_17847(v_17848);
  assign v_17848 = ~v_17843;
  pebbles_core
    pebbles_core_17849
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17850),
       .in0_consume_en(vin0_consume_en_17849),
       .out_canPeek(vout_canPeek_17849),
       .out_peek(vout_peek_17849));
  assign v_17850 = v_17851 | v_17852;
  assign v_17851 = mux_17851(v_17837);
  assign v_17852 = mux_17852(v_17853);
  assign v_17853 = ~v_17837;
  assign v_17854 = v_17855 & 1'h1;
  assign v_17855 = v_17856 & v_17857;
  assign v_17856 = ~act_17836;
  assign v_17857 = v_17858 | v_17866;
  assign v_17858 = v_17859 | v_17864;
  assign v_17859 = mux_17859(v_17860);
  assign v_17860 = v_17833 & v_17861;
  assign v_17861 = v_17862 & 1'h1;
  assign v_17862 = v_17863 | 1'h0;
  assign v_17863 = ~v_17826;
  assign v_17864 = mux_17864(v_17865);
  assign v_17865 = ~v_17860;
  assign v_17866 = ~v_17833;
  assign v_17867 = v_17868 | v_17869;
  assign v_17868 = mux_17868(v_17835);
  assign v_17869 = mux_17869(v_17854);
  assign v_17871 = v_17872 | v_17891;
  assign v_17872 = act_17873 & 1'h1;
  assign act_17873 = v_17874 | v_17880;
  assign v_17874 = v_17875 & v_17881;
  assign v_17875 = v_17876 & vout_canPeek_17886;
  assign v_17876 = ~vout_canPeek_17877;
  pebbles_core
    pebbles_core_17877
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17878),
       .in0_consume_en(vin0_consume_en_17877),
       .out_canPeek(vout_canPeek_17877),
       .out_peek(vout_peek_17877));
  assign v_17878 = v_17879 | v_17884;
  assign v_17879 = mux_17879(v_17880);
  assign v_17880 = vout_canPeek_17877 & v_17881;
  assign v_17881 = v_17882 & 1'h1;
  assign v_17882 = v_17883 | 1'h0;
  assign v_17883 = ~v_17870;
  assign v_17884 = mux_17884(v_17885);
  assign v_17885 = ~v_17880;
  pebbles_core
    pebbles_core_17886
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17887),
       .in0_consume_en(vin0_consume_en_17886),
       .out_canPeek(vout_canPeek_17886),
       .out_peek(vout_peek_17886));
  assign v_17887 = v_17888 | v_17889;
  assign v_17888 = mux_17888(v_17874);
  assign v_17889 = mux_17889(v_17890);
  assign v_17890 = ~v_17874;
  assign v_17891 = v_17892 & 1'h1;
  assign v_17892 = v_17893 & v_17894;
  assign v_17893 = ~act_17873;
  assign v_17894 = v_17895 | v_17899;
  assign v_17895 = v_17896 | v_17897;
  assign v_17896 = mux_17896(v_17830);
  assign v_17897 = mux_17897(v_17898);
  assign v_17898 = ~v_17830;
  assign v_17899 = ~v_17870;
  assign v_17900 = v_17901 | v_17902;
  assign v_17901 = mux_17901(v_17872);
  assign v_17902 = mux_17902(v_17891);
  assign v_17903 = v_17904 & 1'h1;
  assign v_17904 = v_17905 & v_17906;
  assign v_17905 = ~act_17829;
  assign v_17906 = v_17907 | v_17915;
  assign v_17907 = v_17908 | v_17913;
  assign v_17908 = mux_17908(v_17909);
  assign v_17909 = v_17826 & v_17910;
  assign v_17910 = v_17911 & 1'h1;
  assign v_17911 = v_17912 | 1'h0;
  assign v_17912 = ~v_17819;
  assign v_17913 = mux_17913(v_17914);
  assign v_17914 = ~v_17909;
  assign v_17915 = ~v_17826;
  assign v_17916 = v_17917 | v_17918;
  assign v_17917 = mux_17917(v_17828);
  assign v_17918 = mux_17918(v_17903);
  assign v_17920 = v_17921 | v_17996;
  assign v_17921 = act_17922 & 1'h1;
  assign act_17922 = v_17923 | v_17953;
  assign v_17923 = v_17924 & v_17954;
  assign v_17924 = v_17925 & v_17963;
  assign v_17925 = ~v_17926;
  assign v_17927 = v_17928 | v_17947;
  assign v_17928 = act_17929 & 1'h1;
  assign act_17929 = v_17930 | v_17936;
  assign v_17930 = v_17931 & v_17937;
  assign v_17931 = v_17932 & vout_canPeek_17942;
  assign v_17932 = ~vout_canPeek_17933;
  pebbles_core
    pebbles_core_17933
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17934),
       .in0_consume_en(vin0_consume_en_17933),
       .out_canPeek(vout_canPeek_17933),
       .out_peek(vout_peek_17933));
  assign v_17934 = v_17935 | v_17940;
  assign v_17935 = mux_17935(v_17936);
  assign v_17936 = vout_canPeek_17933 & v_17937;
  assign v_17937 = v_17938 & 1'h1;
  assign v_17938 = v_17939 | 1'h0;
  assign v_17939 = ~v_17926;
  assign v_17940 = mux_17940(v_17941);
  assign v_17941 = ~v_17936;
  pebbles_core
    pebbles_core_17942
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17943),
       .in0_consume_en(vin0_consume_en_17942),
       .out_canPeek(vout_canPeek_17942),
       .out_peek(vout_peek_17942));
  assign v_17943 = v_17944 | v_17945;
  assign v_17944 = mux_17944(v_17930);
  assign v_17945 = mux_17945(v_17946);
  assign v_17946 = ~v_17930;
  assign v_17947 = v_17948 & 1'h1;
  assign v_17948 = v_17949 & v_17950;
  assign v_17949 = ~act_17929;
  assign v_17950 = v_17951 | v_17959;
  assign v_17951 = v_17952 | v_17957;
  assign v_17952 = mux_17952(v_17953);
  assign v_17953 = v_17926 & v_17954;
  assign v_17954 = v_17955 & 1'h1;
  assign v_17955 = v_17956 | 1'h0;
  assign v_17956 = ~v_17919;
  assign v_17957 = mux_17957(v_17958);
  assign v_17958 = ~v_17953;
  assign v_17959 = ~v_17926;
  assign v_17960 = v_17961 | v_17962;
  assign v_17961 = mux_17961(v_17928);
  assign v_17962 = mux_17962(v_17947);
  assign v_17964 = v_17965 | v_17984;
  assign v_17965 = act_17966 & 1'h1;
  assign act_17966 = v_17967 | v_17973;
  assign v_17967 = v_17968 & v_17974;
  assign v_17968 = v_17969 & vout_canPeek_17979;
  assign v_17969 = ~vout_canPeek_17970;
  pebbles_core
    pebbles_core_17970
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17971),
       .in0_consume_en(vin0_consume_en_17970),
       .out_canPeek(vout_canPeek_17970),
       .out_peek(vout_peek_17970));
  assign v_17971 = v_17972 | v_17977;
  assign v_17972 = mux_17972(v_17973);
  assign v_17973 = vout_canPeek_17970 & v_17974;
  assign v_17974 = v_17975 & 1'h1;
  assign v_17975 = v_17976 | 1'h0;
  assign v_17976 = ~v_17963;
  assign v_17977 = mux_17977(v_17978);
  assign v_17978 = ~v_17973;
  pebbles_core
    pebbles_core_17979
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_17980),
       .in0_consume_en(vin0_consume_en_17979),
       .out_canPeek(vout_canPeek_17979),
       .out_peek(vout_peek_17979));
  assign v_17980 = v_17981 | v_17982;
  assign v_17981 = mux_17981(v_17967);
  assign v_17982 = mux_17982(v_17983);
  assign v_17983 = ~v_17967;
  assign v_17984 = v_17985 & 1'h1;
  assign v_17985 = v_17986 & v_17987;
  assign v_17986 = ~act_17966;
  assign v_17987 = v_17988 | v_17992;
  assign v_17988 = v_17989 | v_17990;
  assign v_17989 = mux_17989(v_17923);
  assign v_17990 = mux_17990(v_17991);
  assign v_17991 = ~v_17923;
  assign v_17992 = ~v_17963;
  assign v_17993 = v_17994 | v_17995;
  assign v_17994 = mux_17994(v_17965);
  assign v_17995 = mux_17995(v_17984);
  assign v_17996 = v_17997 & 1'h1;
  assign v_17997 = v_17998 & v_17999;
  assign v_17998 = ~act_17922;
  assign v_17999 = v_18000 | v_18004;
  assign v_18000 = v_18001 | v_18002;
  assign v_18001 = mux_18001(v_17823);
  assign v_18002 = mux_18002(v_18003);
  assign v_18003 = ~v_17823;
  assign v_18004 = ~v_17919;
  assign v_18005 = v_18006 | v_18007;
  assign v_18006 = mux_18006(v_17921);
  assign v_18007 = mux_18007(v_17996);
  assign v_18008 = v_18009 & 1'h1;
  assign v_18009 = v_18010 & v_18011;
  assign v_18010 = ~act_17822;
  assign v_18011 = v_18012 | v_18020;
  assign v_18012 = v_18013 | v_18018;
  assign v_18013 = mux_18013(v_18014);
  assign v_18014 = v_17819 & v_18015;
  assign v_18015 = v_18016 & 1'h1;
  assign v_18016 = v_18017 | 1'h0;
  assign v_18017 = ~v_17812;
  assign v_18018 = mux_18018(v_18019);
  assign v_18019 = ~v_18014;
  assign v_18020 = ~v_17819;
  assign v_18021 = v_18022 | v_18023;
  assign v_18022 = mux_18022(v_17821);
  assign v_18023 = mux_18023(v_18008);
  assign v_18025 = v_18026 | v_18213;
  assign v_18026 = act_18027 & 1'h1;
  assign act_18027 = v_18028 | v_18114;
  assign v_18028 = v_18029 & v_18115;
  assign v_18029 = v_18030 & v_18124;
  assign v_18030 = ~v_18031;
  assign v_18032 = v_18033 | v_18108;
  assign v_18033 = act_18034 & 1'h1;
  assign act_18034 = v_18035 | v_18065;
  assign v_18035 = v_18036 & v_18066;
  assign v_18036 = v_18037 & v_18075;
  assign v_18037 = ~v_18038;
  assign v_18039 = v_18040 | v_18059;
  assign v_18040 = act_18041 & 1'h1;
  assign act_18041 = v_18042 | v_18048;
  assign v_18042 = v_18043 & v_18049;
  assign v_18043 = v_18044 & vout_canPeek_18054;
  assign v_18044 = ~vout_canPeek_18045;
  pebbles_core
    pebbles_core_18045
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18046),
       .in0_consume_en(vin0_consume_en_18045),
       .out_canPeek(vout_canPeek_18045),
       .out_peek(vout_peek_18045));
  assign v_18046 = v_18047 | v_18052;
  assign v_18047 = mux_18047(v_18048);
  assign v_18048 = vout_canPeek_18045 & v_18049;
  assign v_18049 = v_18050 & 1'h1;
  assign v_18050 = v_18051 | 1'h0;
  assign v_18051 = ~v_18038;
  assign v_18052 = mux_18052(v_18053);
  assign v_18053 = ~v_18048;
  pebbles_core
    pebbles_core_18054
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18055),
       .in0_consume_en(vin0_consume_en_18054),
       .out_canPeek(vout_canPeek_18054),
       .out_peek(vout_peek_18054));
  assign v_18055 = v_18056 | v_18057;
  assign v_18056 = mux_18056(v_18042);
  assign v_18057 = mux_18057(v_18058);
  assign v_18058 = ~v_18042;
  assign v_18059 = v_18060 & 1'h1;
  assign v_18060 = v_18061 & v_18062;
  assign v_18061 = ~act_18041;
  assign v_18062 = v_18063 | v_18071;
  assign v_18063 = v_18064 | v_18069;
  assign v_18064 = mux_18064(v_18065);
  assign v_18065 = v_18038 & v_18066;
  assign v_18066 = v_18067 & 1'h1;
  assign v_18067 = v_18068 | 1'h0;
  assign v_18068 = ~v_18031;
  assign v_18069 = mux_18069(v_18070);
  assign v_18070 = ~v_18065;
  assign v_18071 = ~v_18038;
  assign v_18072 = v_18073 | v_18074;
  assign v_18073 = mux_18073(v_18040);
  assign v_18074 = mux_18074(v_18059);
  assign v_18076 = v_18077 | v_18096;
  assign v_18077 = act_18078 & 1'h1;
  assign act_18078 = v_18079 | v_18085;
  assign v_18079 = v_18080 & v_18086;
  assign v_18080 = v_18081 & vout_canPeek_18091;
  assign v_18081 = ~vout_canPeek_18082;
  pebbles_core
    pebbles_core_18082
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18083),
       .in0_consume_en(vin0_consume_en_18082),
       .out_canPeek(vout_canPeek_18082),
       .out_peek(vout_peek_18082));
  assign v_18083 = v_18084 | v_18089;
  assign v_18084 = mux_18084(v_18085);
  assign v_18085 = vout_canPeek_18082 & v_18086;
  assign v_18086 = v_18087 & 1'h1;
  assign v_18087 = v_18088 | 1'h0;
  assign v_18088 = ~v_18075;
  assign v_18089 = mux_18089(v_18090);
  assign v_18090 = ~v_18085;
  pebbles_core
    pebbles_core_18091
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18092),
       .in0_consume_en(vin0_consume_en_18091),
       .out_canPeek(vout_canPeek_18091),
       .out_peek(vout_peek_18091));
  assign v_18092 = v_18093 | v_18094;
  assign v_18093 = mux_18093(v_18079);
  assign v_18094 = mux_18094(v_18095);
  assign v_18095 = ~v_18079;
  assign v_18096 = v_18097 & 1'h1;
  assign v_18097 = v_18098 & v_18099;
  assign v_18098 = ~act_18078;
  assign v_18099 = v_18100 | v_18104;
  assign v_18100 = v_18101 | v_18102;
  assign v_18101 = mux_18101(v_18035);
  assign v_18102 = mux_18102(v_18103);
  assign v_18103 = ~v_18035;
  assign v_18104 = ~v_18075;
  assign v_18105 = v_18106 | v_18107;
  assign v_18106 = mux_18106(v_18077);
  assign v_18107 = mux_18107(v_18096);
  assign v_18108 = v_18109 & 1'h1;
  assign v_18109 = v_18110 & v_18111;
  assign v_18110 = ~act_18034;
  assign v_18111 = v_18112 | v_18120;
  assign v_18112 = v_18113 | v_18118;
  assign v_18113 = mux_18113(v_18114);
  assign v_18114 = v_18031 & v_18115;
  assign v_18115 = v_18116 & 1'h1;
  assign v_18116 = v_18117 | 1'h0;
  assign v_18117 = ~v_18024;
  assign v_18118 = mux_18118(v_18119);
  assign v_18119 = ~v_18114;
  assign v_18120 = ~v_18031;
  assign v_18121 = v_18122 | v_18123;
  assign v_18122 = mux_18122(v_18033);
  assign v_18123 = mux_18123(v_18108);
  assign v_18125 = v_18126 | v_18201;
  assign v_18126 = act_18127 & 1'h1;
  assign act_18127 = v_18128 | v_18158;
  assign v_18128 = v_18129 & v_18159;
  assign v_18129 = v_18130 & v_18168;
  assign v_18130 = ~v_18131;
  assign v_18132 = v_18133 | v_18152;
  assign v_18133 = act_18134 & 1'h1;
  assign act_18134 = v_18135 | v_18141;
  assign v_18135 = v_18136 & v_18142;
  assign v_18136 = v_18137 & vout_canPeek_18147;
  assign v_18137 = ~vout_canPeek_18138;
  pebbles_core
    pebbles_core_18138
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18139),
       .in0_consume_en(vin0_consume_en_18138),
       .out_canPeek(vout_canPeek_18138),
       .out_peek(vout_peek_18138));
  assign v_18139 = v_18140 | v_18145;
  assign v_18140 = mux_18140(v_18141);
  assign v_18141 = vout_canPeek_18138 & v_18142;
  assign v_18142 = v_18143 & 1'h1;
  assign v_18143 = v_18144 | 1'h0;
  assign v_18144 = ~v_18131;
  assign v_18145 = mux_18145(v_18146);
  assign v_18146 = ~v_18141;
  pebbles_core
    pebbles_core_18147
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18148),
       .in0_consume_en(vin0_consume_en_18147),
       .out_canPeek(vout_canPeek_18147),
       .out_peek(vout_peek_18147));
  assign v_18148 = v_18149 | v_18150;
  assign v_18149 = mux_18149(v_18135);
  assign v_18150 = mux_18150(v_18151);
  assign v_18151 = ~v_18135;
  assign v_18152 = v_18153 & 1'h1;
  assign v_18153 = v_18154 & v_18155;
  assign v_18154 = ~act_18134;
  assign v_18155 = v_18156 | v_18164;
  assign v_18156 = v_18157 | v_18162;
  assign v_18157 = mux_18157(v_18158);
  assign v_18158 = v_18131 & v_18159;
  assign v_18159 = v_18160 & 1'h1;
  assign v_18160 = v_18161 | 1'h0;
  assign v_18161 = ~v_18124;
  assign v_18162 = mux_18162(v_18163);
  assign v_18163 = ~v_18158;
  assign v_18164 = ~v_18131;
  assign v_18165 = v_18166 | v_18167;
  assign v_18166 = mux_18166(v_18133);
  assign v_18167 = mux_18167(v_18152);
  assign v_18169 = v_18170 | v_18189;
  assign v_18170 = act_18171 & 1'h1;
  assign act_18171 = v_18172 | v_18178;
  assign v_18172 = v_18173 & v_18179;
  assign v_18173 = v_18174 & vout_canPeek_18184;
  assign v_18174 = ~vout_canPeek_18175;
  pebbles_core
    pebbles_core_18175
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18176),
       .in0_consume_en(vin0_consume_en_18175),
       .out_canPeek(vout_canPeek_18175),
       .out_peek(vout_peek_18175));
  assign v_18176 = v_18177 | v_18182;
  assign v_18177 = mux_18177(v_18178);
  assign v_18178 = vout_canPeek_18175 & v_18179;
  assign v_18179 = v_18180 & 1'h1;
  assign v_18180 = v_18181 | 1'h0;
  assign v_18181 = ~v_18168;
  assign v_18182 = mux_18182(v_18183);
  assign v_18183 = ~v_18178;
  pebbles_core
    pebbles_core_18184
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18185),
       .in0_consume_en(vin0_consume_en_18184),
       .out_canPeek(vout_canPeek_18184),
       .out_peek(vout_peek_18184));
  assign v_18185 = v_18186 | v_18187;
  assign v_18186 = mux_18186(v_18172);
  assign v_18187 = mux_18187(v_18188);
  assign v_18188 = ~v_18172;
  assign v_18189 = v_18190 & 1'h1;
  assign v_18190 = v_18191 & v_18192;
  assign v_18191 = ~act_18171;
  assign v_18192 = v_18193 | v_18197;
  assign v_18193 = v_18194 | v_18195;
  assign v_18194 = mux_18194(v_18128);
  assign v_18195 = mux_18195(v_18196);
  assign v_18196 = ~v_18128;
  assign v_18197 = ~v_18168;
  assign v_18198 = v_18199 | v_18200;
  assign v_18199 = mux_18199(v_18170);
  assign v_18200 = mux_18200(v_18189);
  assign v_18201 = v_18202 & 1'h1;
  assign v_18202 = v_18203 & v_18204;
  assign v_18203 = ~act_18127;
  assign v_18204 = v_18205 | v_18209;
  assign v_18205 = v_18206 | v_18207;
  assign v_18206 = mux_18206(v_18028);
  assign v_18207 = mux_18207(v_18208);
  assign v_18208 = ~v_18028;
  assign v_18209 = ~v_18124;
  assign v_18210 = v_18211 | v_18212;
  assign v_18211 = mux_18211(v_18126);
  assign v_18212 = mux_18212(v_18201);
  assign v_18213 = v_18214 & 1'h1;
  assign v_18214 = v_18215 & v_18216;
  assign v_18215 = ~act_18027;
  assign v_18216 = v_18217 | v_18221;
  assign v_18217 = v_18218 | v_18219;
  assign v_18218 = mux_18218(v_17816);
  assign v_18219 = mux_18219(v_18220);
  assign v_18220 = ~v_17816;
  assign v_18221 = ~v_18024;
  assign v_18222 = v_18223 | v_18224;
  assign v_18223 = mux_18223(v_18026);
  assign v_18224 = mux_18224(v_18213);
  assign v_18225 = v_18226 & 1'h1;
  assign v_18226 = v_18227 & v_18228;
  assign v_18227 = ~act_17815;
  assign v_18228 = v_18229 | v_18237;
  assign v_18229 = v_18230 | v_18235;
  assign v_18230 = mux_18230(v_18231);
  assign v_18231 = v_17812 & v_18232;
  assign v_18232 = v_18233 & 1'h1;
  assign v_18233 = v_18234 | 1'h0;
  assign v_18234 = ~v_17805;
  assign v_18235 = mux_18235(v_18236);
  assign v_18236 = ~v_18231;
  assign v_18237 = ~v_17812;
  assign v_18238 = v_18239 | v_18240;
  assign v_18239 = mux_18239(v_17814);
  assign v_18240 = mux_18240(v_18225);
  assign v_18242 = v_18243 | v_18654;
  assign v_18243 = act_18244 & 1'h1;
  assign act_18244 = v_18245 | v_18443;
  assign v_18245 = v_18246 & v_18444;
  assign v_18246 = v_18247 & v_18453;
  assign v_18247 = ~v_18248;
  assign v_18249 = v_18250 | v_18437;
  assign v_18250 = act_18251 & 1'h1;
  assign act_18251 = v_18252 | v_18338;
  assign v_18252 = v_18253 & v_18339;
  assign v_18253 = v_18254 & v_18348;
  assign v_18254 = ~v_18255;
  assign v_18256 = v_18257 | v_18332;
  assign v_18257 = act_18258 & 1'h1;
  assign act_18258 = v_18259 | v_18289;
  assign v_18259 = v_18260 & v_18290;
  assign v_18260 = v_18261 & v_18299;
  assign v_18261 = ~v_18262;
  assign v_18263 = v_18264 | v_18283;
  assign v_18264 = act_18265 & 1'h1;
  assign act_18265 = v_18266 | v_18272;
  assign v_18266 = v_18267 & v_18273;
  assign v_18267 = v_18268 & vout_canPeek_18278;
  assign v_18268 = ~vout_canPeek_18269;
  pebbles_core
    pebbles_core_18269
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18270),
       .in0_consume_en(vin0_consume_en_18269),
       .out_canPeek(vout_canPeek_18269),
       .out_peek(vout_peek_18269));
  assign v_18270 = v_18271 | v_18276;
  assign v_18271 = mux_18271(v_18272);
  assign v_18272 = vout_canPeek_18269 & v_18273;
  assign v_18273 = v_18274 & 1'h1;
  assign v_18274 = v_18275 | 1'h0;
  assign v_18275 = ~v_18262;
  assign v_18276 = mux_18276(v_18277);
  assign v_18277 = ~v_18272;
  pebbles_core
    pebbles_core_18278
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18279),
       .in0_consume_en(vin0_consume_en_18278),
       .out_canPeek(vout_canPeek_18278),
       .out_peek(vout_peek_18278));
  assign v_18279 = v_18280 | v_18281;
  assign v_18280 = mux_18280(v_18266);
  assign v_18281 = mux_18281(v_18282);
  assign v_18282 = ~v_18266;
  assign v_18283 = v_18284 & 1'h1;
  assign v_18284 = v_18285 & v_18286;
  assign v_18285 = ~act_18265;
  assign v_18286 = v_18287 | v_18295;
  assign v_18287 = v_18288 | v_18293;
  assign v_18288 = mux_18288(v_18289);
  assign v_18289 = v_18262 & v_18290;
  assign v_18290 = v_18291 & 1'h1;
  assign v_18291 = v_18292 | 1'h0;
  assign v_18292 = ~v_18255;
  assign v_18293 = mux_18293(v_18294);
  assign v_18294 = ~v_18289;
  assign v_18295 = ~v_18262;
  assign v_18296 = v_18297 | v_18298;
  assign v_18297 = mux_18297(v_18264);
  assign v_18298 = mux_18298(v_18283);
  assign v_18300 = v_18301 | v_18320;
  assign v_18301 = act_18302 & 1'h1;
  assign act_18302 = v_18303 | v_18309;
  assign v_18303 = v_18304 & v_18310;
  assign v_18304 = v_18305 & vout_canPeek_18315;
  assign v_18305 = ~vout_canPeek_18306;
  pebbles_core
    pebbles_core_18306
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18307),
       .in0_consume_en(vin0_consume_en_18306),
       .out_canPeek(vout_canPeek_18306),
       .out_peek(vout_peek_18306));
  assign v_18307 = v_18308 | v_18313;
  assign v_18308 = mux_18308(v_18309);
  assign v_18309 = vout_canPeek_18306 & v_18310;
  assign v_18310 = v_18311 & 1'h1;
  assign v_18311 = v_18312 | 1'h0;
  assign v_18312 = ~v_18299;
  assign v_18313 = mux_18313(v_18314);
  assign v_18314 = ~v_18309;
  pebbles_core
    pebbles_core_18315
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18316),
       .in0_consume_en(vin0_consume_en_18315),
       .out_canPeek(vout_canPeek_18315),
       .out_peek(vout_peek_18315));
  assign v_18316 = v_18317 | v_18318;
  assign v_18317 = mux_18317(v_18303);
  assign v_18318 = mux_18318(v_18319);
  assign v_18319 = ~v_18303;
  assign v_18320 = v_18321 & 1'h1;
  assign v_18321 = v_18322 & v_18323;
  assign v_18322 = ~act_18302;
  assign v_18323 = v_18324 | v_18328;
  assign v_18324 = v_18325 | v_18326;
  assign v_18325 = mux_18325(v_18259);
  assign v_18326 = mux_18326(v_18327);
  assign v_18327 = ~v_18259;
  assign v_18328 = ~v_18299;
  assign v_18329 = v_18330 | v_18331;
  assign v_18330 = mux_18330(v_18301);
  assign v_18331 = mux_18331(v_18320);
  assign v_18332 = v_18333 & 1'h1;
  assign v_18333 = v_18334 & v_18335;
  assign v_18334 = ~act_18258;
  assign v_18335 = v_18336 | v_18344;
  assign v_18336 = v_18337 | v_18342;
  assign v_18337 = mux_18337(v_18338);
  assign v_18338 = v_18255 & v_18339;
  assign v_18339 = v_18340 & 1'h1;
  assign v_18340 = v_18341 | 1'h0;
  assign v_18341 = ~v_18248;
  assign v_18342 = mux_18342(v_18343);
  assign v_18343 = ~v_18338;
  assign v_18344 = ~v_18255;
  assign v_18345 = v_18346 | v_18347;
  assign v_18346 = mux_18346(v_18257);
  assign v_18347 = mux_18347(v_18332);
  assign v_18349 = v_18350 | v_18425;
  assign v_18350 = act_18351 & 1'h1;
  assign act_18351 = v_18352 | v_18382;
  assign v_18352 = v_18353 & v_18383;
  assign v_18353 = v_18354 & v_18392;
  assign v_18354 = ~v_18355;
  assign v_18356 = v_18357 | v_18376;
  assign v_18357 = act_18358 & 1'h1;
  assign act_18358 = v_18359 | v_18365;
  assign v_18359 = v_18360 & v_18366;
  assign v_18360 = v_18361 & vout_canPeek_18371;
  assign v_18361 = ~vout_canPeek_18362;
  pebbles_core
    pebbles_core_18362
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18363),
       .in0_consume_en(vin0_consume_en_18362),
       .out_canPeek(vout_canPeek_18362),
       .out_peek(vout_peek_18362));
  assign v_18363 = v_18364 | v_18369;
  assign v_18364 = mux_18364(v_18365);
  assign v_18365 = vout_canPeek_18362 & v_18366;
  assign v_18366 = v_18367 & 1'h1;
  assign v_18367 = v_18368 | 1'h0;
  assign v_18368 = ~v_18355;
  assign v_18369 = mux_18369(v_18370);
  assign v_18370 = ~v_18365;
  pebbles_core
    pebbles_core_18371
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18372),
       .in0_consume_en(vin0_consume_en_18371),
       .out_canPeek(vout_canPeek_18371),
       .out_peek(vout_peek_18371));
  assign v_18372 = v_18373 | v_18374;
  assign v_18373 = mux_18373(v_18359);
  assign v_18374 = mux_18374(v_18375);
  assign v_18375 = ~v_18359;
  assign v_18376 = v_18377 & 1'h1;
  assign v_18377 = v_18378 & v_18379;
  assign v_18378 = ~act_18358;
  assign v_18379 = v_18380 | v_18388;
  assign v_18380 = v_18381 | v_18386;
  assign v_18381 = mux_18381(v_18382);
  assign v_18382 = v_18355 & v_18383;
  assign v_18383 = v_18384 & 1'h1;
  assign v_18384 = v_18385 | 1'h0;
  assign v_18385 = ~v_18348;
  assign v_18386 = mux_18386(v_18387);
  assign v_18387 = ~v_18382;
  assign v_18388 = ~v_18355;
  assign v_18389 = v_18390 | v_18391;
  assign v_18390 = mux_18390(v_18357);
  assign v_18391 = mux_18391(v_18376);
  assign v_18393 = v_18394 | v_18413;
  assign v_18394 = act_18395 & 1'h1;
  assign act_18395 = v_18396 | v_18402;
  assign v_18396 = v_18397 & v_18403;
  assign v_18397 = v_18398 & vout_canPeek_18408;
  assign v_18398 = ~vout_canPeek_18399;
  pebbles_core
    pebbles_core_18399
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18400),
       .in0_consume_en(vin0_consume_en_18399),
       .out_canPeek(vout_canPeek_18399),
       .out_peek(vout_peek_18399));
  assign v_18400 = v_18401 | v_18406;
  assign v_18401 = mux_18401(v_18402);
  assign v_18402 = vout_canPeek_18399 & v_18403;
  assign v_18403 = v_18404 & 1'h1;
  assign v_18404 = v_18405 | 1'h0;
  assign v_18405 = ~v_18392;
  assign v_18406 = mux_18406(v_18407);
  assign v_18407 = ~v_18402;
  pebbles_core
    pebbles_core_18408
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18409),
       .in0_consume_en(vin0_consume_en_18408),
       .out_canPeek(vout_canPeek_18408),
       .out_peek(vout_peek_18408));
  assign v_18409 = v_18410 | v_18411;
  assign v_18410 = mux_18410(v_18396);
  assign v_18411 = mux_18411(v_18412);
  assign v_18412 = ~v_18396;
  assign v_18413 = v_18414 & 1'h1;
  assign v_18414 = v_18415 & v_18416;
  assign v_18415 = ~act_18395;
  assign v_18416 = v_18417 | v_18421;
  assign v_18417 = v_18418 | v_18419;
  assign v_18418 = mux_18418(v_18352);
  assign v_18419 = mux_18419(v_18420);
  assign v_18420 = ~v_18352;
  assign v_18421 = ~v_18392;
  assign v_18422 = v_18423 | v_18424;
  assign v_18423 = mux_18423(v_18394);
  assign v_18424 = mux_18424(v_18413);
  assign v_18425 = v_18426 & 1'h1;
  assign v_18426 = v_18427 & v_18428;
  assign v_18427 = ~act_18351;
  assign v_18428 = v_18429 | v_18433;
  assign v_18429 = v_18430 | v_18431;
  assign v_18430 = mux_18430(v_18252);
  assign v_18431 = mux_18431(v_18432);
  assign v_18432 = ~v_18252;
  assign v_18433 = ~v_18348;
  assign v_18434 = v_18435 | v_18436;
  assign v_18435 = mux_18435(v_18350);
  assign v_18436 = mux_18436(v_18425);
  assign v_18437 = v_18438 & 1'h1;
  assign v_18438 = v_18439 & v_18440;
  assign v_18439 = ~act_18251;
  assign v_18440 = v_18441 | v_18449;
  assign v_18441 = v_18442 | v_18447;
  assign v_18442 = mux_18442(v_18443);
  assign v_18443 = v_18248 & v_18444;
  assign v_18444 = v_18445 & 1'h1;
  assign v_18445 = v_18446 | 1'h0;
  assign v_18446 = ~v_18241;
  assign v_18447 = mux_18447(v_18448);
  assign v_18448 = ~v_18443;
  assign v_18449 = ~v_18248;
  assign v_18450 = v_18451 | v_18452;
  assign v_18451 = mux_18451(v_18250);
  assign v_18452 = mux_18452(v_18437);
  assign v_18454 = v_18455 | v_18642;
  assign v_18455 = act_18456 & 1'h1;
  assign act_18456 = v_18457 | v_18543;
  assign v_18457 = v_18458 & v_18544;
  assign v_18458 = v_18459 & v_18553;
  assign v_18459 = ~v_18460;
  assign v_18461 = v_18462 | v_18537;
  assign v_18462 = act_18463 & 1'h1;
  assign act_18463 = v_18464 | v_18494;
  assign v_18464 = v_18465 & v_18495;
  assign v_18465 = v_18466 & v_18504;
  assign v_18466 = ~v_18467;
  assign v_18468 = v_18469 | v_18488;
  assign v_18469 = act_18470 & 1'h1;
  assign act_18470 = v_18471 | v_18477;
  assign v_18471 = v_18472 & v_18478;
  assign v_18472 = v_18473 & vout_canPeek_18483;
  assign v_18473 = ~vout_canPeek_18474;
  pebbles_core
    pebbles_core_18474
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18475),
       .in0_consume_en(vin0_consume_en_18474),
       .out_canPeek(vout_canPeek_18474),
       .out_peek(vout_peek_18474));
  assign v_18475 = v_18476 | v_18481;
  assign v_18476 = mux_18476(v_18477);
  assign v_18477 = vout_canPeek_18474 & v_18478;
  assign v_18478 = v_18479 & 1'h1;
  assign v_18479 = v_18480 | 1'h0;
  assign v_18480 = ~v_18467;
  assign v_18481 = mux_18481(v_18482);
  assign v_18482 = ~v_18477;
  pebbles_core
    pebbles_core_18483
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18484),
       .in0_consume_en(vin0_consume_en_18483),
       .out_canPeek(vout_canPeek_18483),
       .out_peek(vout_peek_18483));
  assign v_18484 = v_18485 | v_18486;
  assign v_18485 = mux_18485(v_18471);
  assign v_18486 = mux_18486(v_18487);
  assign v_18487 = ~v_18471;
  assign v_18488 = v_18489 & 1'h1;
  assign v_18489 = v_18490 & v_18491;
  assign v_18490 = ~act_18470;
  assign v_18491 = v_18492 | v_18500;
  assign v_18492 = v_18493 | v_18498;
  assign v_18493 = mux_18493(v_18494);
  assign v_18494 = v_18467 & v_18495;
  assign v_18495 = v_18496 & 1'h1;
  assign v_18496 = v_18497 | 1'h0;
  assign v_18497 = ~v_18460;
  assign v_18498 = mux_18498(v_18499);
  assign v_18499 = ~v_18494;
  assign v_18500 = ~v_18467;
  assign v_18501 = v_18502 | v_18503;
  assign v_18502 = mux_18502(v_18469);
  assign v_18503 = mux_18503(v_18488);
  assign v_18505 = v_18506 | v_18525;
  assign v_18506 = act_18507 & 1'h1;
  assign act_18507 = v_18508 | v_18514;
  assign v_18508 = v_18509 & v_18515;
  assign v_18509 = v_18510 & vout_canPeek_18520;
  assign v_18510 = ~vout_canPeek_18511;
  pebbles_core
    pebbles_core_18511
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18512),
       .in0_consume_en(vin0_consume_en_18511),
       .out_canPeek(vout_canPeek_18511),
       .out_peek(vout_peek_18511));
  assign v_18512 = v_18513 | v_18518;
  assign v_18513 = mux_18513(v_18514);
  assign v_18514 = vout_canPeek_18511 & v_18515;
  assign v_18515 = v_18516 & 1'h1;
  assign v_18516 = v_18517 | 1'h0;
  assign v_18517 = ~v_18504;
  assign v_18518 = mux_18518(v_18519);
  assign v_18519 = ~v_18514;
  pebbles_core
    pebbles_core_18520
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18521),
       .in0_consume_en(vin0_consume_en_18520),
       .out_canPeek(vout_canPeek_18520),
       .out_peek(vout_peek_18520));
  assign v_18521 = v_18522 | v_18523;
  assign v_18522 = mux_18522(v_18508);
  assign v_18523 = mux_18523(v_18524);
  assign v_18524 = ~v_18508;
  assign v_18525 = v_18526 & 1'h1;
  assign v_18526 = v_18527 & v_18528;
  assign v_18527 = ~act_18507;
  assign v_18528 = v_18529 | v_18533;
  assign v_18529 = v_18530 | v_18531;
  assign v_18530 = mux_18530(v_18464);
  assign v_18531 = mux_18531(v_18532);
  assign v_18532 = ~v_18464;
  assign v_18533 = ~v_18504;
  assign v_18534 = v_18535 | v_18536;
  assign v_18535 = mux_18535(v_18506);
  assign v_18536 = mux_18536(v_18525);
  assign v_18537 = v_18538 & 1'h1;
  assign v_18538 = v_18539 & v_18540;
  assign v_18539 = ~act_18463;
  assign v_18540 = v_18541 | v_18549;
  assign v_18541 = v_18542 | v_18547;
  assign v_18542 = mux_18542(v_18543);
  assign v_18543 = v_18460 & v_18544;
  assign v_18544 = v_18545 & 1'h1;
  assign v_18545 = v_18546 | 1'h0;
  assign v_18546 = ~v_18453;
  assign v_18547 = mux_18547(v_18548);
  assign v_18548 = ~v_18543;
  assign v_18549 = ~v_18460;
  assign v_18550 = v_18551 | v_18552;
  assign v_18551 = mux_18551(v_18462);
  assign v_18552 = mux_18552(v_18537);
  assign v_18554 = v_18555 | v_18630;
  assign v_18555 = act_18556 & 1'h1;
  assign act_18556 = v_18557 | v_18587;
  assign v_18557 = v_18558 & v_18588;
  assign v_18558 = v_18559 & v_18597;
  assign v_18559 = ~v_18560;
  assign v_18561 = v_18562 | v_18581;
  assign v_18562 = act_18563 & 1'h1;
  assign act_18563 = v_18564 | v_18570;
  assign v_18564 = v_18565 & v_18571;
  assign v_18565 = v_18566 & vout_canPeek_18576;
  assign v_18566 = ~vout_canPeek_18567;
  pebbles_core
    pebbles_core_18567
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18568),
       .in0_consume_en(vin0_consume_en_18567),
       .out_canPeek(vout_canPeek_18567),
       .out_peek(vout_peek_18567));
  assign v_18568 = v_18569 | v_18574;
  assign v_18569 = mux_18569(v_18570);
  assign v_18570 = vout_canPeek_18567 & v_18571;
  assign v_18571 = v_18572 & 1'h1;
  assign v_18572 = v_18573 | 1'h0;
  assign v_18573 = ~v_18560;
  assign v_18574 = mux_18574(v_18575);
  assign v_18575 = ~v_18570;
  pebbles_core
    pebbles_core_18576
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18577),
       .in0_consume_en(vin0_consume_en_18576),
       .out_canPeek(vout_canPeek_18576),
       .out_peek(vout_peek_18576));
  assign v_18577 = v_18578 | v_18579;
  assign v_18578 = mux_18578(v_18564);
  assign v_18579 = mux_18579(v_18580);
  assign v_18580 = ~v_18564;
  assign v_18581 = v_18582 & 1'h1;
  assign v_18582 = v_18583 & v_18584;
  assign v_18583 = ~act_18563;
  assign v_18584 = v_18585 | v_18593;
  assign v_18585 = v_18586 | v_18591;
  assign v_18586 = mux_18586(v_18587);
  assign v_18587 = v_18560 & v_18588;
  assign v_18588 = v_18589 & 1'h1;
  assign v_18589 = v_18590 | 1'h0;
  assign v_18590 = ~v_18553;
  assign v_18591 = mux_18591(v_18592);
  assign v_18592 = ~v_18587;
  assign v_18593 = ~v_18560;
  assign v_18594 = v_18595 | v_18596;
  assign v_18595 = mux_18595(v_18562);
  assign v_18596 = mux_18596(v_18581);
  assign v_18598 = v_18599 | v_18618;
  assign v_18599 = act_18600 & 1'h1;
  assign act_18600 = v_18601 | v_18607;
  assign v_18601 = v_18602 & v_18608;
  assign v_18602 = v_18603 & vout_canPeek_18613;
  assign v_18603 = ~vout_canPeek_18604;
  pebbles_core
    pebbles_core_18604
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18605),
       .in0_consume_en(vin0_consume_en_18604),
       .out_canPeek(vout_canPeek_18604),
       .out_peek(vout_peek_18604));
  assign v_18605 = v_18606 | v_18611;
  assign v_18606 = mux_18606(v_18607);
  assign v_18607 = vout_canPeek_18604 & v_18608;
  assign v_18608 = v_18609 & 1'h1;
  assign v_18609 = v_18610 | 1'h0;
  assign v_18610 = ~v_18597;
  assign v_18611 = mux_18611(v_18612);
  assign v_18612 = ~v_18607;
  pebbles_core
    pebbles_core_18613
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18614),
       .in0_consume_en(vin0_consume_en_18613),
       .out_canPeek(vout_canPeek_18613),
       .out_peek(vout_peek_18613));
  assign v_18614 = v_18615 | v_18616;
  assign v_18615 = mux_18615(v_18601);
  assign v_18616 = mux_18616(v_18617);
  assign v_18617 = ~v_18601;
  assign v_18618 = v_18619 & 1'h1;
  assign v_18619 = v_18620 & v_18621;
  assign v_18620 = ~act_18600;
  assign v_18621 = v_18622 | v_18626;
  assign v_18622 = v_18623 | v_18624;
  assign v_18623 = mux_18623(v_18557);
  assign v_18624 = mux_18624(v_18625);
  assign v_18625 = ~v_18557;
  assign v_18626 = ~v_18597;
  assign v_18627 = v_18628 | v_18629;
  assign v_18628 = mux_18628(v_18599);
  assign v_18629 = mux_18629(v_18618);
  assign v_18630 = v_18631 & 1'h1;
  assign v_18631 = v_18632 & v_18633;
  assign v_18632 = ~act_18556;
  assign v_18633 = v_18634 | v_18638;
  assign v_18634 = v_18635 | v_18636;
  assign v_18635 = mux_18635(v_18457);
  assign v_18636 = mux_18636(v_18637);
  assign v_18637 = ~v_18457;
  assign v_18638 = ~v_18553;
  assign v_18639 = v_18640 | v_18641;
  assign v_18640 = mux_18640(v_18555);
  assign v_18641 = mux_18641(v_18630);
  assign v_18642 = v_18643 & 1'h1;
  assign v_18643 = v_18644 & v_18645;
  assign v_18644 = ~act_18456;
  assign v_18645 = v_18646 | v_18650;
  assign v_18646 = v_18647 | v_18648;
  assign v_18647 = mux_18647(v_18245);
  assign v_18648 = mux_18648(v_18649);
  assign v_18649 = ~v_18245;
  assign v_18650 = ~v_18453;
  assign v_18651 = v_18652 | v_18653;
  assign v_18652 = mux_18652(v_18455);
  assign v_18653 = mux_18653(v_18642);
  assign v_18654 = v_18655 & 1'h1;
  assign v_18655 = v_18656 & v_18657;
  assign v_18656 = ~act_18244;
  assign v_18657 = v_18658 | v_18662;
  assign v_18658 = v_18659 | v_18660;
  assign v_18659 = mux_18659(v_17809);
  assign v_18660 = mux_18660(v_18661);
  assign v_18661 = ~v_17809;
  assign v_18662 = ~v_18241;
  assign v_18663 = v_18664 | v_18665;
  assign v_18664 = mux_18664(v_18243);
  assign v_18665 = mux_18665(v_18654);
  assign v_18666 = v_18667 & 1'h1;
  assign v_18667 = v_18668 & v_18669;
  assign v_18668 = ~act_17808;
  assign v_18669 = v_18670 | v_18674;
  assign v_18670 = v_18671 | v_18672;
  assign v_18671 = mux_18671(v_16925);
  assign v_18672 = mux_18672(v_18673);
  assign v_18673 = ~v_16925;
  assign v_18674 = ~v_17805;
  assign v_18675 = v_18676 | v_18677;
  assign v_18676 = mux_18676(v_17807);
  assign v_18677 = mux_18677(v_18666);
  assign v_18678 = v_18679 & 1'h1;
  assign v_18679 = v_18680 & v_18681;
  assign v_18680 = ~act_16924;
  assign v_18681 = v_18682 | v_18686;
  assign v_18682 = v_18683 | v_18684;
  assign v_18683 = mux_18683(v_15145);
  assign v_18684 = mux_18684(v_18685);
  assign v_18685 = ~v_15145;
  assign v_18686 = ~v_16921;
  assign v_18687 = v_18688 | v_18689;
  assign v_18688 = mux_18688(v_16923);
  assign v_18689 = mux_18689(v_18678);
  assign v_18690 = v_18691 & 1'h1;
  assign v_18691 = v_18692 & v_18693;
  assign v_18692 = ~act_15144;
  assign v_18693 = v_18694 | v_18702;
  assign v_18694 = v_18695 | v_18700;
  assign v_18695 = mux_18695(v_18696);
  assign v_18696 = v_15141 & v_18697;
  assign v_18697 = v_18698 & 1'h1;
  assign v_18698 = v_18699 | 1'h0;
  assign v_18699 = ~v_15134;
  assign v_18700 = mux_18700(v_18701);
  assign v_18701 = ~v_18696;
  assign v_18702 = ~v_15141;
  assign v_18703 = v_18704 | v_18705;
  assign v_18704 = mux_18704(v_15143);
  assign v_18705 = mux_18705(v_18690);
  assign v_18707 = v_18708 | v_22255;
  assign v_18708 = act_18709 & 1'h1;
  assign act_18709 = v_18710 | v_20476;
  assign v_18710 = v_18711 & v_20477;
  assign v_18711 = v_18712 & v_20486;
  assign v_18712 = ~v_18713;
  assign v_18714 = v_18715 | v_20470;
  assign v_18715 = act_18716 & 1'h1;
  assign act_18716 = v_18717 | v_19587;
  assign v_18717 = v_18718 & v_19588;
  assign v_18718 = v_18719 & v_19597;
  assign v_18719 = ~v_18720;
  assign v_18721 = v_18722 | v_19581;
  assign v_18722 = act_18723 & 1'h1;
  assign act_18723 = v_18724 | v_19146;
  assign v_18724 = v_18725 & v_19147;
  assign v_18725 = v_18726 & v_19156;
  assign v_18726 = ~v_18727;
  assign v_18728 = v_18729 | v_19140;
  assign v_18729 = act_18730 & 1'h1;
  assign act_18730 = v_18731 | v_18929;
  assign v_18731 = v_18732 & v_18930;
  assign v_18732 = v_18733 & v_18939;
  assign v_18733 = ~v_18734;
  assign v_18735 = v_18736 | v_18923;
  assign v_18736 = act_18737 & 1'h1;
  assign act_18737 = v_18738 | v_18824;
  assign v_18738 = v_18739 & v_18825;
  assign v_18739 = v_18740 & v_18834;
  assign v_18740 = ~v_18741;
  assign v_18742 = v_18743 | v_18818;
  assign v_18743 = act_18744 & 1'h1;
  assign act_18744 = v_18745 | v_18775;
  assign v_18745 = v_18746 & v_18776;
  assign v_18746 = v_18747 & v_18785;
  assign v_18747 = ~v_18748;
  assign v_18749 = v_18750 | v_18769;
  assign v_18750 = act_18751 & 1'h1;
  assign act_18751 = v_18752 | v_18758;
  assign v_18752 = v_18753 & v_18759;
  assign v_18753 = v_18754 & vout_canPeek_18764;
  assign v_18754 = ~vout_canPeek_18755;
  pebbles_core
    pebbles_core_18755
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18756),
       .in0_consume_en(vin0_consume_en_18755),
       .out_canPeek(vout_canPeek_18755),
       .out_peek(vout_peek_18755));
  assign v_18756 = v_18757 | v_18762;
  assign v_18757 = mux_18757(v_18758);
  assign v_18758 = vout_canPeek_18755 & v_18759;
  assign v_18759 = v_18760 & 1'h1;
  assign v_18760 = v_18761 | 1'h0;
  assign v_18761 = ~v_18748;
  assign v_18762 = mux_18762(v_18763);
  assign v_18763 = ~v_18758;
  pebbles_core
    pebbles_core_18764
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18765),
       .in0_consume_en(vin0_consume_en_18764),
       .out_canPeek(vout_canPeek_18764),
       .out_peek(vout_peek_18764));
  assign v_18765 = v_18766 | v_18767;
  assign v_18766 = mux_18766(v_18752);
  assign v_18767 = mux_18767(v_18768);
  assign v_18768 = ~v_18752;
  assign v_18769 = v_18770 & 1'h1;
  assign v_18770 = v_18771 & v_18772;
  assign v_18771 = ~act_18751;
  assign v_18772 = v_18773 | v_18781;
  assign v_18773 = v_18774 | v_18779;
  assign v_18774 = mux_18774(v_18775);
  assign v_18775 = v_18748 & v_18776;
  assign v_18776 = v_18777 & 1'h1;
  assign v_18777 = v_18778 | 1'h0;
  assign v_18778 = ~v_18741;
  assign v_18779 = mux_18779(v_18780);
  assign v_18780 = ~v_18775;
  assign v_18781 = ~v_18748;
  assign v_18782 = v_18783 | v_18784;
  assign v_18783 = mux_18783(v_18750);
  assign v_18784 = mux_18784(v_18769);
  assign v_18786 = v_18787 | v_18806;
  assign v_18787 = act_18788 & 1'h1;
  assign act_18788 = v_18789 | v_18795;
  assign v_18789 = v_18790 & v_18796;
  assign v_18790 = v_18791 & vout_canPeek_18801;
  assign v_18791 = ~vout_canPeek_18792;
  pebbles_core
    pebbles_core_18792
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18793),
       .in0_consume_en(vin0_consume_en_18792),
       .out_canPeek(vout_canPeek_18792),
       .out_peek(vout_peek_18792));
  assign v_18793 = v_18794 | v_18799;
  assign v_18794 = mux_18794(v_18795);
  assign v_18795 = vout_canPeek_18792 & v_18796;
  assign v_18796 = v_18797 & 1'h1;
  assign v_18797 = v_18798 | 1'h0;
  assign v_18798 = ~v_18785;
  assign v_18799 = mux_18799(v_18800);
  assign v_18800 = ~v_18795;
  pebbles_core
    pebbles_core_18801
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18802),
       .in0_consume_en(vin0_consume_en_18801),
       .out_canPeek(vout_canPeek_18801),
       .out_peek(vout_peek_18801));
  assign v_18802 = v_18803 | v_18804;
  assign v_18803 = mux_18803(v_18789);
  assign v_18804 = mux_18804(v_18805);
  assign v_18805 = ~v_18789;
  assign v_18806 = v_18807 & 1'h1;
  assign v_18807 = v_18808 & v_18809;
  assign v_18808 = ~act_18788;
  assign v_18809 = v_18810 | v_18814;
  assign v_18810 = v_18811 | v_18812;
  assign v_18811 = mux_18811(v_18745);
  assign v_18812 = mux_18812(v_18813);
  assign v_18813 = ~v_18745;
  assign v_18814 = ~v_18785;
  assign v_18815 = v_18816 | v_18817;
  assign v_18816 = mux_18816(v_18787);
  assign v_18817 = mux_18817(v_18806);
  assign v_18818 = v_18819 & 1'h1;
  assign v_18819 = v_18820 & v_18821;
  assign v_18820 = ~act_18744;
  assign v_18821 = v_18822 | v_18830;
  assign v_18822 = v_18823 | v_18828;
  assign v_18823 = mux_18823(v_18824);
  assign v_18824 = v_18741 & v_18825;
  assign v_18825 = v_18826 & 1'h1;
  assign v_18826 = v_18827 | 1'h0;
  assign v_18827 = ~v_18734;
  assign v_18828 = mux_18828(v_18829);
  assign v_18829 = ~v_18824;
  assign v_18830 = ~v_18741;
  assign v_18831 = v_18832 | v_18833;
  assign v_18832 = mux_18832(v_18743);
  assign v_18833 = mux_18833(v_18818);
  assign v_18835 = v_18836 | v_18911;
  assign v_18836 = act_18837 & 1'h1;
  assign act_18837 = v_18838 | v_18868;
  assign v_18838 = v_18839 & v_18869;
  assign v_18839 = v_18840 & v_18878;
  assign v_18840 = ~v_18841;
  assign v_18842 = v_18843 | v_18862;
  assign v_18843 = act_18844 & 1'h1;
  assign act_18844 = v_18845 | v_18851;
  assign v_18845 = v_18846 & v_18852;
  assign v_18846 = v_18847 & vout_canPeek_18857;
  assign v_18847 = ~vout_canPeek_18848;
  pebbles_core
    pebbles_core_18848
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18849),
       .in0_consume_en(vin0_consume_en_18848),
       .out_canPeek(vout_canPeek_18848),
       .out_peek(vout_peek_18848));
  assign v_18849 = v_18850 | v_18855;
  assign v_18850 = mux_18850(v_18851);
  assign v_18851 = vout_canPeek_18848 & v_18852;
  assign v_18852 = v_18853 & 1'h1;
  assign v_18853 = v_18854 | 1'h0;
  assign v_18854 = ~v_18841;
  assign v_18855 = mux_18855(v_18856);
  assign v_18856 = ~v_18851;
  pebbles_core
    pebbles_core_18857
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18858),
       .in0_consume_en(vin0_consume_en_18857),
       .out_canPeek(vout_canPeek_18857),
       .out_peek(vout_peek_18857));
  assign v_18858 = v_18859 | v_18860;
  assign v_18859 = mux_18859(v_18845);
  assign v_18860 = mux_18860(v_18861);
  assign v_18861 = ~v_18845;
  assign v_18862 = v_18863 & 1'h1;
  assign v_18863 = v_18864 & v_18865;
  assign v_18864 = ~act_18844;
  assign v_18865 = v_18866 | v_18874;
  assign v_18866 = v_18867 | v_18872;
  assign v_18867 = mux_18867(v_18868);
  assign v_18868 = v_18841 & v_18869;
  assign v_18869 = v_18870 & 1'h1;
  assign v_18870 = v_18871 | 1'h0;
  assign v_18871 = ~v_18834;
  assign v_18872 = mux_18872(v_18873);
  assign v_18873 = ~v_18868;
  assign v_18874 = ~v_18841;
  assign v_18875 = v_18876 | v_18877;
  assign v_18876 = mux_18876(v_18843);
  assign v_18877 = mux_18877(v_18862);
  assign v_18879 = v_18880 | v_18899;
  assign v_18880 = act_18881 & 1'h1;
  assign act_18881 = v_18882 | v_18888;
  assign v_18882 = v_18883 & v_18889;
  assign v_18883 = v_18884 & vout_canPeek_18894;
  assign v_18884 = ~vout_canPeek_18885;
  pebbles_core
    pebbles_core_18885
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18886),
       .in0_consume_en(vin0_consume_en_18885),
       .out_canPeek(vout_canPeek_18885),
       .out_peek(vout_peek_18885));
  assign v_18886 = v_18887 | v_18892;
  assign v_18887 = mux_18887(v_18888);
  assign v_18888 = vout_canPeek_18885 & v_18889;
  assign v_18889 = v_18890 & 1'h1;
  assign v_18890 = v_18891 | 1'h0;
  assign v_18891 = ~v_18878;
  assign v_18892 = mux_18892(v_18893);
  assign v_18893 = ~v_18888;
  pebbles_core
    pebbles_core_18894
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18895),
       .in0_consume_en(vin0_consume_en_18894),
       .out_canPeek(vout_canPeek_18894),
       .out_peek(vout_peek_18894));
  assign v_18895 = v_18896 | v_18897;
  assign v_18896 = mux_18896(v_18882);
  assign v_18897 = mux_18897(v_18898);
  assign v_18898 = ~v_18882;
  assign v_18899 = v_18900 & 1'h1;
  assign v_18900 = v_18901 & v_18902;
  assign v_18901 = ~act_18881;
  assign v_18902 = v_18903 | v_18907;
  assign v_18903 = v_18904 | v_18905;
  assign v_18904 = mux_18904(v_18838);
  assign v_18905 = mux_18905(v_18906);
  assign v_18906 = ~v_18838;
  assign v_18907 = ~v_18878;
  assign v_18908 = v_18909 | v_18910;
  assign v_18909 = mux_18909(v_18880);
  assign v_18910 = mux_18910(v_18899);
  assign v_18911 = v_18912 & 1'h1;
  assign v_18912 = v_18913 & v_18914;
  assign v_18913 = ~act_18837;
  assign v_18914 = v_18915 | v_18919;
  assign v_18915 = v_18916 | v_18917;
  assign v_18916 = mux_18916(v_18738);
  assign v_18917 = mux_18917(v_18918);
  assign v_18918 = ~v_18738;
  assign v_18919 = ~v_18834;
  assign v_18920 = v_18921 | v_18922;
  assign v_18921 = mux_18921(v_18836);
  assign v_18922 = mux_18922(v_18911);
  assign v_18923 = v_18924 & 1'h1;
  assign v_18924 = v_18925 & v_18926;
  assign v_18925 = ~act_18737;
  assign v_18926 = v_18927 | v_18935;
  assign v_18927 = v_18928 | v_18933;
  assign v_18928 = mux_18928(v_18929);
  assign v_18929 = v_18734 & v_18930;
  assign v_18930 = v_18931 & 1'h1;
  assign v_18931 = v_18932 | 1'h0;
  assign v_18932 = ~v_18727;
  assign v_18933 = mux_18933(v_18934);
  assign v_18934 = ~v_18929;
  assign v_18935 = ~v_18734;
  assign v_18936 = v_18937 | v_18938;
  assign v_18937 = mux_18937(v_18736);
  assign v_18938 = mux_18938(v_18923);
  assign v_18940 = v_18941 | v_19128;
  assign v_18941 = act_18942 & 1'h1;
  assign act_18942 = v_18943 | v_19029;
  assign v_18943 = v_18944 & v_19030;
  assign v_18944 = v_18945 & v_19039;
  assign v_18945 = ~v_18946;
  assign v_18947 = v_18948 | v_19023;
  assign v_18948 = act_18949 & 1'h1;
  assign act_18949 = v_18950 | v_18980;
  assign v_18950 = v_18951 & v_18981;
  assign v_18951 = v_18952 & v_18990;
  assign v_18952 = ~v_18953;
  assign v_18954 = v_18955 | v_18974;
  assign v_18955 = act_18956 & 1'h1;
  assign act_18956 = v_18957 | v_18963;
  assign v_18957 = v_18958 & v_18964;
  assign v_18958 = v_18959 & vout_canPeek_18969;
  assign v_18959 = ~vout_canPeek_18960;
  pebbles_core
    pebbles_core_18960
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18961),
       .in0_consume_en(vin0_consume_en_18960),
       .out_canPeek(vout_canPeek_18960),
       .out_peek(vout_peek_18960));
  assign v_18961 = v_18962 | v_18967;
  assign v_18962 = mux_18962(v_18963);
  assign v_18963 = vout_canPeek_18960 & v_18964;
  assign v_18964 = v_18965 & 1'h1;
  assign v_18965 = v_18966 | 1'h0;
  assign v_18966 = ~v_18953;
  assign v_18967 = mux_18967(v_18968);
  assign v_18968 = ~v_18963;
  pebbles_core
    pebbles_core_18969
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18970),
       .in0_consume_en(vin0_consume_en_18969),
       .out_canPeek(vout_canPeek_18969),
       .out_peek(vout_peek_18969));
  assign v_18970 = v_18971 | v_18972;
  assign v_18971 = mux_18971(v_18957);
  assign v_18972 = mux_18972(v_18973);
  assign v_18973 = ~v_18957;
  assign v_18974 = v_18975 & 1'h1;
  assign v_18975 = v_18976 & v_18977;
  assign v_18976 = ~act_18956;
  assign v_18977 = v_18978 | v_18986;
  assign v_18978 = v_18979 | v_18984;
  assign v_18979 = mux_18979(v_18980);
  assign v_18980 = v_18953 & v_18981;
  assign v_18981 = v_18982 & 1'h1;
  assign v_18982 = v_18983 | 1'h0;
  assign v_18983 = ~v_18946;
  assign v_18984 = mux_18984(v_18985);
  assign v_18985 = ~v_18980;
  assign v_18986 = ~v_18953;
  assign v_18987 = v_18988 | v_18989;
  assign v_18988 = mux_18988(v_18955);
  assign v_18989 = mux_18989(v_18974);
  assign v_18991 = v_18992 | v_19011;
  assign v_18992 = act_18993 & 1'h1;
  assign act_18993 = v_18994 | v_19000;
  assign v_18994 = v_18995 & v_19001;
  assign v_18995 = v_18996 & vout_canPeek_19006;
  assign v_18996 = ~vout_canPeek_18997;
  pebbles_core
    pebbles_core_18997
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_18998),
       .in0_consume_en(vin0_consume_en_18997),
       .out_canPeek(vout_canPeek_18997),
       .out_peek(vout_peek_18997));
  assign v_18998 = v_18999 | v_19004;
  assign v_18999 = mux_18999(v_19000);
  assign v_19000 = vout_canPeek_18997 & v_19001;
  assign v_19001 = v_19002 & 1'h1;
  assign v_19002 = v_19003 | 1'h0;
  assign v_19003 = ~v_18990;
  assign v_19004 = mux_19004(v_19005);
  assign v_19005 = ~v_19000;
  pebbles_core
    pebbles_core_19006
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19007),
       .in0_consume_en(vin0_consume_en_19006),
       .out_canPeek(vout_canPeek_19006),
       .out_peek(vout_peek_19006));
  assign v_19007 = v_19008 | v_19009;
  assign v_19008 = mux_19008(v_18994);
  assign v_19009 = mux_19009(v_19010);
  assign v_19010 = ~v_18994;
  assign v_19011 = v_19012 & 1'h1;
  assign v_19012 = v_19013 & v_19014;
  assign v_19013 = ~act_18993;
  assign v_19014 = v_19015 | v_19019;
  assign v_19015 = v_19016 | v_19017;
  assign v_19016 = mux_19016(v_18950);
  assign v_19017 = mux_19017(v_19018);
  assign v_19018 = ~v_18950;
  assign v_19019 = ~v_18990;
  assign v_19020 = v_19021 | v_19022;
  assign v_19021 = mux_19021(v_18992);
  assign v_19022 = mux_19022(v_19011);
  assign v_19023 = v_19024 & 1'h1;
  assign v_19024 = v_19025 & v_19026;
  assign v_19025 = ~act_18949;
  assign v_19026 = v_19027 | v_19035;
  assign v_19027 = v_19028 | v_19033;
  assign v_19028 = mux_19028(v_19029);
  assign v_19029 = v_18946 & v_19030;
  assign v_19030 = v_19031 & 1'h1;
  assign v_19031 = v_19032 | 1'h0;
  assign v_19032 = ~v_18939;
  assign v_19033 = mux_19033(v_19034);
  assign v_19034 = ~v_19029;
  assign v_19035 = ~v_18946;
  assign v_19036 = v_19037 | v_19038;
  assign v_19037 = mux_19037(v_18948);
  assign v_19038 = mux_19038(v_19023);
  assign v_19040 = v_19041 | v_19116;
  assign v_19041 = act_19042 & 1'h1;
  assign act_19042 = v_19043 | v_19073;
  assign v_19043 = v_19044 & v_19074;
  assign v_19044 = v_19045 & v_19083;
  assign v_19045 = ~v_19046;
  assign v_19047 = v_19048 | v_19067;
  assign v_19048 = act_19049 & 1'h1;
  assign act_19049 = v_19050 | v_19056;
  assign v_19050 = v_19051 & v_19057;
  assign v_19051 = v_19052 & vout_canPeek_19062;
  assign v_19052 = ~vout_canPeek_19053;
  pebbles_core
    pebbles_core_19053
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19054),
       .in0_consume_en(vin0_consume_en_19053),
       .out_canPeek(vout_canPeek_19053),
       .out_peek(vout_peek_19053));
  assign v_19054 = v_19055 | v_19060;
  assign v_19055 = mux_19055(v_19056);
  assign v_19056 = vout_canPeek_19053 & v_19057;
  assign v_19057 = v_19058 & 1'h1;
  assign v_19058 = v_19059 | 1'h0;
  assign v_19059 = ~v_19046;
  assign v_19060 = mux_19060(v_19061);
  assign v_19061 = ~v_19056;
  pebbles_core
    pebbles_core_19062
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19063),
       .in0_consume_en(vin0_consume_en_19062),
       .out_canPeek(vout_canPeek_19062),
       .out_peek(vout_peek_19062));
  assign v_19063 = v_19064 | v_19065;
  assign v_19064 = mux_19064(v_19050);
  assign v_19065 = mux_19065(v_19066);
  assign v_19066 = ~v_19050;
  assign v_19067 = v_19068 & 1'h1;
  assign v_19068 = v_19069 & v_19070;
  assign v_19069 = ~act_19049;
  assign v_19070 = v_19071 | v_19079;
  assign v_19071 = v_19072 | v_19077;
  assign v_19072 = mux_19072(v_19073);
  assign v_19073 = v_19046 & v_19074;
  assign v_19074 = v_19075 & 1'h1;
  assign v_19075 = v_19076 | 1'h0;
  assign v_19076 = ~v_19039;
  assign v_19077 = mux_19077(v_19078);
  assign v_19078 = ~v_19073;
  assign v_19079 = ~v_19046;
  assign v_19080 = v_19081 | v_19082;
  assign v_19081 = mux_19081(v_19048);
  assign v_19082 = mux_19082(v_19067);
  assign v_19084 = v_19085 | v_19104;
  assign v_19085 = act_19086 & 1'h1;
  assign act_19086 = v_19087 | v_19093;
  assign v_19087 = v_19088 & v_19094;
  assign v_19088 = v_19089 & vout_canPeek_19099;
  assign v_19089 = ~vout_canPeek_19090;
  pebbles_core
    pebbles_core_19090
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19091),
       .in0_consume_en(vin0_consume_en_19090),
       .out_canPeek(vout_canPeek_19090),
       .out_peek(vout_peek_19090));
  assign v_19091 = v_19092 | v_19097;
  assign v_19092 = mux_19092(v_19093);
  assign v_19093 = vout_canPeek_19090 & v_19094;
  assign v_19094 = v_19095 & 1'h1;
  assign v_19095 = v_19096 | 1'h0;
  assign v_19096 = ~v_19083;
  assign v_19097 = mux_19097(v_19098);
  assign v_19098 = ~v_19093;
  pebbles_core
    pebbles_core_19099
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19100),
       .in0_consume_en(vin0_consume_en_19099),
       .out_canPeek(vout_canPeek_19099),
       .out_peek(vout_peek_19099));
  assign v_19100 = v_19101 | v_19102;
  assign v_19101 = mux_19101(v_19087);
  assign v_19102 = mux_19102(v_19103);
  assign v_19103 = ~v_19087;
  assign v_19104 = v_19105 & 1'h1;
  assign v_19105 = v_19106 & v_19107;
  assign v_19106 = ~act_19086;
  assign v_19107 = v_19108 | v_19112;
  assign v_19108 = v_19109 | v_19110;
  assign v_19109 = mux_19109(v_19043);
  assign v_19110 = mux_19110(v_19111);
  assign v_19111 = ~v_19043;
  assign v_19112 = ~v_19083;
  assign v_19113 = v_19114 | v_19115;
  assign v_19114 = mux_19114(v_19085);
  assign v_19115 = mux_19115(v_19104);
  assign v_19116 = v_19117 & 1'h1;
  assign v_19117 = v_19118 & v_19119;
  assign v_19118 = ~act_19042;
  assign v_19119 = v_19120 | v_19124;
  assign v_19120 = v_19121 | v_19122;
  assign v_19121 = mux_19121(v_18943);
  assign v_19122 = mux_19122(v_19123);
  assign v_19123 = ~v_18943;
  assign v_19124 = ~v_19039;
  assign v_19125 = v_19126 | v_19127;
  assign v_19126 = mux_19126(v_19041);
  assign v_19127 = mux_19127(v_19116);
  assign v_19128 = v_19129 & 1'h1;
  assign v_19129 = v_19130 & v_19131;
  assign v_19130 = ~act_18942;
  assign v_19131 = v_19132 | v_19136;
  assign v_19132 = v_19133 | v_19134;
  assign v_19133 = mux_19133(v_18731);
  assign v_19134 = mux_19134(v_19135);
  assign v_19135 = ~v_18731;
  assign v_19136 = ~v_18939;
  assign v_19137 = v_19138 | v_19139;
  assign v_19138 = mux_19138(v_18941);
  assign v_19139 = mux_19139(v_19128);
  assign v_19140 = v_19141 & 1'h1;
  assign v_19141 = v_19142 & v_19143;
  assign v_19142 = ~act_18730;
  assign v_19143 = v_19144 | v_19152;
  assign v_19144 = v_19145 | v_19150;
  assign v_19145 = mux_19145(v_19146);
  assign v_19146 = v_18727 & v_19147;
  assign v_19147 = v_19148 & 1'h1;
  assign v_19148 = v_19149 | 1'h0;
  assign v_19149 = ~v_18720;
  assign v_19150 = mux_19150(v_19151);
  assign v_19151 = ~v_19146;
  assign v_19152 = ~v_18727;
  assign v_19153 = v_19154 | v_19155;
  assign v_19154 = mux_19154(v_18729);
  assign v_19155 = mux_19155(v_19140);
  assign v_19157 = v_19158 | v_19569;
  assign v_19158 = act_19159 & 1'h1;
  assign act_19159 = v_19160 | v_19358;
  assign v_19160 = v_19161 & v_19359;
  assign v_19161 = v_19162 & v_19368;
  assign v_19162 = ~v_19163;
  assign v_19164 = v_19165 | v_19352;
  assign v_19165 = act_19166 & 1'h1;
  assign act_19166 = v_19167 | v_19253;
  assign v_19167 = v_19168 & v_19254;
  assign v_19168 = v_19169 & v_19263;
  assign v_19169 = ~v_19170;
  assign v_19171 = v_19172 | v_19247;
  assign v_19172 = act_19173 & 1'h1;
  assign act_19173 = v_19174 | v_19204;
  assign v_19174 = v_19175 & v_19205;
  assign v_19175 = v_19176 & v_19214;
  assign v_19176 = ~v_19177;
  assign v_19178 = v_19179 | v_19198;
  assign v_19179 = act_19180 & 1'h1;
  assign act_19180 = v_19181 | v_19187;
  assign v_19181 = v_19182 & v_19188;
  assign v_19182 = v_19183 & vout_canPeek_19193;
  assign v_19183 = ~vout_canPeek_19184;
  pebbles_core
    pebbles_core_19184
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19185),
       .in0_consume_en(vin0_consume_en_19184),
       .out_canPeek(vout_canPeek_19184),
       .out_peek(vout_peek_19184));
  assign v_19185 = v_19186 | v_19191;
  assign v_19186 = mux_19186(v_19187);
  assign v_19187 = vout_canPeek_19184 & v_19188;
  assign v_19188 = v_19189 & 1'h1;
  assign v_19189 = v_19190 | 1'h0;
  assign v_19190 = ~v_19177;
  assign v_19191 = mux_19191(v_19192);
  assign v_19192 = ~v_19187;
  pebbles_core
    pebbles_core_19193
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19194),
       .in0_consume_en(vin0_consume_en_19193),
       .out_canPeek(vout_canPeek_19193),
       .out_peek(vout_peek_19193));
  assign v_19194 = v_19195 | v_19196;
  assign v_19195 = mux_19195(v_19181);
  assign v_19196 = mux_19196(v_19197);
  assign v_19197 = ~v_19181;
  assign v_19198 = v_19199 & 1'h1;
  assign v_19199 = v_19200 & v_19201;
  assign v_19200 = ~act_19180;
  assign v_19201 = v_19202 | v_19210;
  assign v_19202 = v_19203 | v_19208;
  assign v_19203 = mux_19203(v_19204);
  assign v_19204 = v_19177 & v_19205;
  assign v_19205 = v_19206 & 1'h1;
  assign v_19206 = v_19207 | 1'h0;
  assign v_19207 = ~v_19170;
  assign v_19208 = mux_19208(v_19209);
  assign v_19209 = ~v_19204;
  assign v_19210 = ~v_19177;
  assign v_19211 = v_19212 | v_19213;
  assign v_19212 = mux_19212(v_19179);
  assign v_19213 = mux_19213(v_19198);
  assign v_19215 = v_19216 | v_19235;
  assign v_19216 = act_19217 & 1'h1;
  assign act_19217 = v_19218 | v_19224;
  assign v_19218 = v_19219 & v_19225;
  assign v_19219 = v_19220 & vout_canPeek_19230;
  assign v_19220 = ~vout_canPeek_19221;
  pebbles_core
    pebbles_core_19221
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19222),
       .in0_consume_en(vin0_consume_en_19221),
       .out_canPeek(vout_canPeek_19221),
       .out_peek(vout_peek_19221));
  assign v_19222 = v_19223 | v_19228;
  assign v_19223 = mux_19223(v_19224);
  assign v_19224 = vout_canPeek_19221 & v_19225;
  assign v_19225 = v_19226 & 1'h1;
  assign v_19226 = v_19227 | 1'h0;
  assign v_19227 = ~v_19214;
  assign v_19228 = mux_19228(v_19229);
  assign v_19229 = ~v_19224;
  pebbles_core
    pebbles_core_19230
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19231),
       .in0_consume_en(vin0_consume_en_19230),
       .out_canPeek(vout_canPeek_19230),
       .out_peek(vout_peek_19230));
  assign v_19231 = v_19232 | v_19233;
  assign v_19232 = mux_19232(v_19218);
  assign v_19233 = mux_19233(v_19234);
  assign v_19234 = ~v_19218;
  assign v_19235 = v_19236 & 1'h1;
  assign v_19236 = v_19237 & v_19238;
  assign v_19237 = ~act_19217;
  assign v_19238 = v_19239 | v_19243;
  assign v_19239 = v_19240 | v_19241;
  assign v_19240 = mux_19240(v_19174);
  assign v_19241 = mux_19241(v_19242);
  assign v_19242 = ~v_19174;
  assign v_19243 = ~v_19214;
  assign v_19244 = v_19245 | v_19246;
  assign v_19245 = mux_19245(v_19216);
  assign v_19246 = mux_19246(v_19235);
  assign v_19247 = v_19248 & 1'h1;
  assign v_19248 = v_19249 & v_19250;
  assign v_19249 = ~act_19173;
  assign v_19250 = v_19251 | v_19259;
  assign v_19251 = v_19252 | v_19257;
  assign v_19252 = mux_19252(v_19253);
  assign v_19253 = v_19170 & v_19254;
  assign v_19254 = v_19255 & 1'h1;
  assign v_19255 = v_19256 | 1'h0;
  assign v_19256 = ~v_19163;
  assign v_19257 = mux_19257(v_19258);
  assign v_19258 = ~v_19253;
  assign v_19259 = ~v_19170;
  assign v_19260 = v_19261 | v_19262;
  assign v_19261 = mux_19261(v_19172);
  assign v_19262 = mux_19262(v_19247);
  assign v_19264 = v_19265 | v_19340;
  assign v_19265 = act_19266 & 1'h1;
  assign act_19266 = v_19267 | v_19297;
  assign v_19267 = v_19268 & v_19298;
  assign v_19268 = v_19269 & v_19307;
  assign v_19269 = ~v_19270;
  assign v_19271 = v_19272 | v_19291;
  assign v_19272 = act_19273 & 1'h1;
  assign act_19273 = v_19274 | v_19280;
  assign v_19274 = v_19275 & v_19281;
  assign v_19275 = v_19276 & vout_canPeek_19286;
  assign v_19276 = ~vout_canPeek_19277;
  pebbles_core
    pebbles_core_19277
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19278),
       .in0_consume_en(vin0_consume_en_19277),
       .out_canPeek(vout_canPeek_19277),
       .out_peek(vout_peek_19277));
  assign v_19278 = v_19279 | v_19284;
  assign v_19279 = mux_19279(v_19280);
  assign v_19280 = vout_canPeek_19277 & v_19281;
  assign v_19281 = v_19282 & 1'h1;
  assign v_19282 = v_19283 | 1'h0;
  assign v_19283 = ~v_19270;
  assign v_19284 = mux_19284(v_19285);
  assign v_19285 = ~v_19280;
  pebbles_core
    pebbles_core_19286
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19287),
       .in0_consume_en(vin0_consume_en_19286),
       .out_canPeek(vout_canPeek_19286),
       .out_peek(vout_peek_19286));
  assign v_19287 = v_19288 | v_19289;
  assign v_19288 = mux_19288(v_19274);
  assign v_19289 = mux_19289(v_19290);
  assign v_19290 = ~v_19274;
  assign v_19291 = v_19292 & 1'h1;
  assign v_19292 = v_19293 & v_19294;
  assign v_19293 = ~act_19273;
  assign v_19294 = v_19295 | v_19303;
  assign v_19295 = v_19296 | v_19301;
  assign v_19296 = mux_19296(v_19297);
  assign v_19297 = v_19270 & v_19298;
  assign v_19298 = v_19299 & 1'h1;
  assign v_19299 = v_19300 | 1'h0;
  assign v_19300 = ~v_19263;
  assign v_19301 = mux_19301(v_19302);
  assign v_19302 = ~v_19297;
  assign v_19303 = ~v_19270;
  assign v_19304 = v_19305 | v_19306;
  assign v_19305 = mux_19305(v_19272);
  assign v_19306 = mux_19306(v_19291);
  assign v_19308 = v_19309 | v_19328;
  assign v_19309 = act_19310 & 1'h1;
  assign act_19310 = v_19311 | v_19317;
  assign v_19311 = v_19312 & v_19318;
  assign v_19312 = v_19313 & vout_canPeek_19323;
  assign v_19313 = ~vout_canPeek_19314;
  pebbles_core
    pebbles_core_19314
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19315),
       .in0_consume_en(vin0_consume_en_19314),
       .out_canPeek(vout_canPeek_19314),
       .out_peek(vout_peek_19314));
  assign v_19315 = v_19316 | v_19321;
  assign v_19316 = mux_19316(v_19317);
  assign v_19317 = vout_canPeek_19314 & v_19318;
  assign v_19318 = v_19319 & 1'h1;
  assign v_19319 = v_19320 | 1'h0;
  assign v_19320 = ~v_19307;
  assign v_19321 = mux_19321(v_19322);
  assign v_19322 = ~v_19317;
  pebbles_core
    pebbles_core_19323
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19324),
       .in0_consume_en(vin0_consume_en_19323),
       .out_canPeek(vout_canPeek_19323),
       .out_peek(vout_peek_19323));
  assign v_19324 = v_19325 | v_19326;
  assign v_19325 = mux_19325(v_19311);
  assign v_19326 = mux_19326(v_19327);
  assign v_19327 = ~v_19311;
  assign v_19328 = v_19329 & 1'h1;
  assign v_19329 = v_19330 & v_19331;
  assign v_19330 = ~act_19310;
  assign v_19331 = v_19332 | v_19336;
  assign v_19332 = v_19333 | v_19334;
  assign v_19333 = mux_19333(v_19267);
  assign v_19334 = mux_19334(v_19335);
  assign v_19335 = ~v_19267;
  assign v_19336 = ~v_19307;
  assign v_19337 = v_19338 | v_19339;
  assign v_19338 = mux_19338(v_19309);
  assign v_19339 = mux_19339(v_19328);
  assign v_19340 = v_19341 & 1'h1;
  assign v_19341 = v_19342 & v_19343;
  assign v_19342 = ~act_19266;
  assign v_19343 = v_19344 | v_19348;
  assign v_19344 = v_19345 | v_19346;
  assign v_19345 = mux_19345(v_19167);
  assign v_19346 = mux_19346(v_19347);
  assign v_19347 = ~v_19167;
  assign v_19348 = ~v_19263;
  assign v_19349 = v_19350 | v_19351;
  assign v_19350 = mux_19350(v_19265);
  assign v_19351 = mux_19351(v_19340);
  assign v_19352 = v_19353 & 1'h1;
  assign v_19353 = v_19354 & v_19355;
  assign v_19354 = ~act_19166;
  assign v_19355 = v_19356 | v_19364;
  assign v_19356 = v_19357 | v_19362;
  assign v_19357 = mux_19357(v_19358);
  assign v_19358 = v_19163 & v_19359;
  assign v_19359 = v_19360 & 1'h1;
  assign v_19360 = v_19361 | 1'h0;
  assign v_19361 = ~v_19156;
  assign v_19362 = mux_19362(v_19363);
  assign v_19363 = ~v_19358;
  assign v_19364 = ~v_19163;
  assign v_19365 = v_19366 | v_19367;
  assign v_19366 = mux_19366(v_19165);
  assign v_19367 = mux_19367(v_19352);
  assign v_19369 = v_19370 | v_19557;
  assign v_19370 = act_19371 & 1'h1;
  assign act_19371 = v_19372 | v_19458;
  assign v_19372 = v_19373 & v_19459;
  assign v_19373 = v_19374 & v_19468;
  assign v_19374 = ~v_19375;
  assign v_19376 = v_19377 | v_19452;
  assign v_19377 = act_19378 & 1'h1;
  assign act_19378 = v_19379 | v_19409;
  assign v_19379 = v_19380 & v_19410;
  assign v_19380 = v_19381 & v_19419;
  assign v_19381 = ~v_19382;
  assign v_19383 = v_19384 | v_19403;
  assign v_19384 = act_19385 & 1'h1;
  assign act_19385 = v_19386 | v_19392;
  assign v_19386 = v_19387 & v_19393;
  assign v_19387 = v_19388 & vout_canPeek_19398;
  assign v_19388 = ~vout_canPeek_19389;
  pebbles_core
    pebbles_core_19389
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19390),
       .in0_consume_en(vin0_consume_en_19389),
       .out_canPeek(vout_canPeek_19389),
       .out_peek(vout_peek_19389));
  assign v_19390 = v_19391 | v_19396;
  assign v_19391 = mux_19391(v_19392);
  assign v_19392 = vout_canPeek_19389 & v_19393;
  assign v_19393 = v_19394 & 1'h1;
  assign v_19394 = v_19395 | 1'h0;
  assign v_19395 = ~v_19382;
  assign v_19396 = mux_19396(v_19397);
  assign v_19397 = ~v_19392;
  pebbles_core
    pebbles_core_19398
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19399),
       .in0_consume_en(vin0_consume_en_19398),
       .out_canPeek(vout_canPeek_19398),
       .out_peek(vout_peek_19398));
  assign v_19399 = v_19400 | v_19401;
  assign v_19400 = mux_19400(v_19386);
  assign v_19401 = mux_19401(v_19402);
  assign v_19402 = ~v_19386;
  assign v_19403 = v_19404 & 1'h1;
  assign v_19404 = v_19405 & v_19406;
  assign v_19405 = ~act_19385;
  assign v_19406 = v_19407 | v_19415;
  assign v_19407 = v_19408 | v_19413;
  assign v_19408 = mux_19408(v_19409);
  assign v_19409 = v_19382 & v_19410;
  assign v_19410 = v_19411 & 1'h1;
  assign v_19411 = v_19412 | 1'h0;
  assign v_19412 = ~v_19375;
  assign v_19413 = mux_19413(v_19414);
  assign v_19414 = ~v_19409;
  assign v_19415 = ~v_19382;
  assign v_19416 = v_19417 | v_19418;
  assign v_19417 = mux_19417(v_19384);
  assign v_19418 = mux_19418(v_19403);
  assign v_19420 = v_19421 | v_19440;
  assign v_19421 = act_19422 & 1'h1;
  assign act_19422 = v_19423 | v_19429;
  assign v_19423 = v_19424 & v_19430;
  assign v_19424 = v_19425 & vout_canPeek_19435;
  assign v_19425 = ~vout_canPeek_19426;
  pebbles_core
    pebbles_core_19426
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19427),
       .in0_consume_en(vin0_consume_en_19426),
       .out_canPeek(vout_canPeek_19426),
       .out_peek(vout_peek_19426));
  assign v_19427 = v_19428 | v_19433;
  assign v_19428 = mux_19428(v_19429);
  assign v_19429 = vout_canPeek_19426 & v_19430;
  assign v_19430 = v_19431 & 1'h1;
  assign v_19431 = v_19432 | 1'h0;
  assign v_19432 = ~v_19419;
  assign v_19433 = mux_19433(v_19434);
  assign v_19434 = ~v_19429;
  pebbles_core
    pebbles_core_19435
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19436),
       .in0_consume_en(vin0_consume_en_19435),
       .out_canPeek(vout_canPeek_19435),
       .out_peek(vout_peek_19435));
  assign v_19436 = v_19437 | v_19438;
  assign v_19437 = mux_19437(v_19423);
  assign v_19438 = mux_19438(v_19439);
  assign v_19439 = ~v_19423;
  assign v_19440 = v_19441 & 1'h1;
  assign v_19441 = v_19442 & v_19443;
  assign v_19442 = ~act_19422;
  assign v_19443 = v_19444 | v_19448;
  assign v_19444 = v_19445 | v_19446;
  assign v_19445 = mux_19445(v_19379);
  assign v_19446 = mux_19446(v_19447);
  assign v_19447 = ~v_19379;
  assign v_19448 = ~v_19419;
  assign v_19449 = v_19450 | v_19451;
  assign v_19450 = mux_19450(v_19421);
  assign v_19451 = mux_19451(v_19440);
  assign v_19452 = v_19453 & 1'h1;
  assign v_19453 = v_19454 & v_19455;
  assign v_19454 = ~act_19378;
  assign v_19455 = v_19456 | v_19464;
  assign v_19456 = v_19457 | v_19462;
  assign v_19457 = mux_19457(v_19458);
  assign v_19458 = v_19375 & v_19459;
  assign v_19459 = v_19460 & 1'h1;
  assign v_19460 = v_19461 | 1'h0;
  assign v_19461 = ~v_19368;
  assign v_19462 = mux_19462(v_19463);
  assign v_19463 = ~v_19458;
  assign v_19464 = ~v_19375;
  assign v_19465 = v_19466 | v_19467;
  assign v_19466 = mux_19466(v_19377);
  assign v_19467 = mux_19467(v_19452);
  assign v_19469 = v_19470 | v_19545;
  assign v_19470 = act_19471 & 1'h1;
  assign act_19471 = v_19472 | v_19502;
  assign v_19472 = v_19473 & v_19503;
  assign v_19473 = v_19474 & v_19512;
  assign v_19474 = ~v_19475;
  assign v_19476 = v_19477 | v_19496;
  assign v_19477 = act_19478 & 1'h1;
  assign act_19478 = v_19479 | v_19485;
  assign v_19479 = v_19480 & v_19486;
  assign v_19480 = v_19481 & vout_canPeek_19491;
  assign v_19481 = ~vout_canPeek_19482;
  pebbles_core
    pebbles_core_19482
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19483),
       .in0_consume_en(vin0_consume_en_19482),
       .out_canPeek(vout_canPeek_19482),
       .out_peek(vout_peek_19482));
  assign v_19483 = v_19484 | v_19489;
  assign v_19484 = mux_19484(v_19485);
  assign v_19485 = vout_canPeek_19482 & v_19486;
  assign v_19486 = v_19487 & 1'h1;
  assign v_19487 = v_19488 | 1'h0;
  assign v_19488 = ~v_19475;
  assign v_19489 = mux_19489(v_19490);
  assign v_19490 = ~v_19485;
  pebbles_core
    pebbles_core_19491
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19492),
       .in0_consume_en(vin0_consume_en_19491),
       .out_canPeek(vout_canPeek_19491),
       .out_peek(vout_peek_19491));
  assign v_19492 = v_19493 | v_19494;
  assign v_19493 = mux_19493(v_19479);
  assign v_19494 = mux_19494(v_19495);
  assign v_19495 = ~v_19479;
  assign v_19496 = v_19497 & 1'h1;
  assign v_19497 = v_19498 & v_19499;
  assign v_19498 = ~act_19478;
  assign v_19499 = v_19500 | v_19508;
  assign v_19500 = v_19501 | v_19506;
  assign v_19501 = mux_19501(v_19502);
  assign v_19502 = v_19475 & v_19503;
  assign v_19503 = v_19504 & 1'h1;
  assign v_19504 = v_19505 | 1'h0;
  assign v_19505 = ~v_19468;
  assign v_19506 = mux_19506(v_19507);
  assign v_19507 = ~v_19502;
  assign v_19508 = ~v_19475;
  assign v_19509 = v_19510 | v_19511;
  assign v_19510 = mux_19510(v_19477);
  assign v_19511 = mux_19511(v_19496);
  assign v_19513 = v_19514 | v_19533;
  assign v_19514 = act_19515 & 1'h1;
  assign act_19515 = v_19516 | v_19522;
  assign v_19516 = v_19517 & v_19523;
  assign v_19517 = v_19518 & vout_canPeek_19528;
  assign v_19518 = ~vout_canPeek_19519;
  pebbles_core
    pebbles_core_19519
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19520),
       .in0_consume_en(vin0_consume_en_19519),
       .out_canPeek(vout_canPeek_19519),
       .out_peek(vout_peek_19519));
  assign v_19520 = v_19521 | v_19526;
  assign v_19521 = mux_19521(v_19522);
  assign v_19522 = vout_canPeek_19519 & v_19523;
  assign v_19523 = v_19524 & 1'h1;
  assign v_19524 = v_19525 | 1'h0;
  assign v_19525 = ~v_19512;
  assign v_19526 = mux_19526(v_19527);
  assign v_19527 = ~v_19522;
  pebbles_core
    pebbles_core_19528
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19529),
       .in0_consume_en(vin0_consume_en_19528),
       .out_canPeek(vout_canPeek_19528),
       .out_peek(vout_peek_19528));
  assign v_19529 = v_19530 | v_19531;
  assign v_19530 = mux_19530(v_19516);
  assign v_19531 = mux_19531(v_19532);
  assign v_19532 = ~v_19516;
  assign v_19533 = v_19534 & 1'h1;
  assign v_19534 = v_19535 & v_19536;
  assign v_19535 = ~act_19515;
  assign v_19536 = v_19537 | v_19541;
  assign v_19537 = v_19538 | v_19539;
  assign v_19538 = mux_19538(v_19472);
  assign v_19539 = mux_19539(v_19540);
  assign v_19540 = ~v_19472;
  assign v_19541 = ~v_19512;
  assign v_19542 = v_19543 | v_19544;
  assign v_19543 = mux_19543(v_19514);
  assign v_19544 = mux_19544(v_19533);
  assign v_19545 = v_19546 & 1'h1;
  assign v_19546 = v_19547 & v_19548;
  assign v_19547 = ~act_19471;
  assign v_19548 = v_19549 | v_19553;
  assign v_19549 = v_19550 | v_19551;
  assign v_19550 = mux_19550(v_19372);
  assign v_19551 = mux_19551(v_19552);
  assign v_19552 = ~v_19372;
  assign v_19553 = ~v_19468;
  assign v_19554 = v_19555 | v_19556;
  assign v_19555 = mux_19555(v_19470);
  assign v_19556 = mux_19556(v_19545);
  assign v_19557 = v_19558 & 1'h1;
  assign v_19558 = v_19559 & v_19560;
  assign v_19559 = ~act_19371;
  assign v_19560 = v_19561 | v_19565;
  assign v_19561 = v_19562 | v_19563;
  assign v_19562 = mux_19562(v_19160);
  assign v_19563 = mux_19563(v_19564);
  assign v_19564 = ~v_19160;
  assign v_19565 = ~v_19368;
  assign v_19566 = v_19567 | v_19568;
  assign v_19567 = mux_19567(v_19370);
  assign v_19568 = mux_19568(v_19557);
  assign v_19569 = v_19570 & 1'h1;
  assign v_19570 = v_19571 & v_19572;
  assign v_19571 = ~act_19159;
  assign v_19572 = v_19573 | v_19577;
  assign v_19573 = v_19574 | v_19575;
  assign v_19574 = mux_19574(v_18724);
  assign v_19575 = mux_19575(v_19576);
  assign v_19576 = ~v_18724;
  assign v_19577 = ~v_19156;
  assign v_19578 = v_19579 | v_19580;
  assign v_19579 = mux_19579(v_19158);
  assign v_19580 = mux_19580(v_19569);
  assign v_19581 = v_19582 & 1'h1;
  assign v_19582 = v_19583 & v_19584;
  assign v_19583 = ~act_18723;
  assign v_19584 = v_19585 | v_19593;
  assign v_19585 = v_19586 | v_19591;
  assign v_19586 = mux_19586(v_19587);
  assign v_19587 = v_18720 & v_19588;
  assign v_19588 = v_19589 & 1'h1;
  assign v_19589 = v_19590 | 1'h0;
  assign v_19590 = ~v_18713;
  assign v_19591 = mux_19591(v_19592);
  assign v_19592 = ~v_19587;
  assign v_19593 = ~v_18720;
  assign v_19594 = v_19595 | v_19596;
  assign v_19595 = mux_19595(v_18722);
  assign v_19596 = mux_19596(v_19581);
  assign v_19598 = v_19599 | v_20458;
  assign v_19599 = act_19600 & 1'h1;
  assign act_19600 = v_19601 | v_20023;
  assign v_19601 = v_19602 & v_20024;
  assign v_19602 = v_19603 & v_20033;
  assign v_19603 = ~v_19604;
  assign v_19605 = v_19606 | v_20017;
  assign v_19606 = act_19607 & 1'h1;
  assign act_19607 = v_19608 | v_19806;
  assign v_19608 = v_19609 & v_19807;
  assign v_19609 = v_19610 & v_19816;
  assign v_19610 = ~v_19611;
  assign v_19612 = v_19613 | v_19800;
  assign v_19613 = act_19614 & 1'h1;
  assign act_19614 = v_19615 | v_19701;
  assign v_19615 = v_19616 & v_19702;
  assign v_19616 = v_19617 & v_19711;
  assign v_19617 = ~v_19618;
  assign v_19619 = v_19620 | v_19695;
  assign v_19620 = act_19621 & 1'h1;
  assign act_19621 = v_19622 | v_19652;
  assign v_19622 = v_19623 & v_19653;
  assign v_19623 = v_19624 & v_19662;
  assign v_19624 = ~v_19625;
  assign v_19626 = v_19627 | v_19646;
  assign v_19627 = act_19628 & 1'h1;
  assign act_19628 = v_19629 | v_19635;
  assign v_19629 = v_19630 & v_19636;
  assign v_19630 = v_19631 & vout_canPeek_19641;
  assign v_19631 = ~vout_canPeek_19632;
  pebbles_core
    pebbles_core_19632
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19633),
       .in0_consume_en(vin0_consume_en_19632),
       .out_canPeek(vout_canPeek_19632),
       .out_peek(vout_peek_19632));
  assign v_19633 = v_19634 | v_19639;
  assign v_19634 = mux_19634(v_19635);
  assign v_19635 = vout_canPeek_19632 & v_19636;
  assign v_19636 = v_19637 & 1'h1;
  assign v_19637 = v_19638 | 1'h0;
  assign v_19638 = ~v_19625;
  assign v_19639 = mux_19639(v_19640);
  assign v_19640 = ~v_19635;
  pebbles_core
    pebbles_core_19641
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19642),
       .in0_consume_en(vin0_consume_en_19641),
       .out_canPeek(vout_canPeek_19641),
       .out_peek(vout_peek_19641));
  assign v_19642 = v_19643 | v_19644;
  assign v_19643 = mux_19643(v_19629);
  assign v_19644 = mux_19644(v_19645);
  assign v_19645 = ~v_19629;
  assign v_19646 = v_19647 & 1'h1;
  assign v_19647 = v_19648 & v_19649;
  assign v_19648 = ~act_19628;
  assign v_19649 = v_19650 | v_19658;
  assign v_19650 = v_19651 | v_19656;
  assign v_19651 = mux_19651(v_19652);
  assign v_19652 = v_19625 & v_19653;
  assign v_19653 = v_19654 & 1'h1;
  assign v_19654 = v_19655 | 1'h0;
  assign v_19655 = ~v_19618;
  assign v_19656 = mux_19656(v_19657);
  assign v_19657 = ~v_19652;
  assign v_19658 = ~v_19625;
  assign v_19659 = v_19660 | v_19661;
  assign v_19660 = mux_19660(v_19627);
  assign v_19661 = mux_19661(v_19646);
  assign v_19663 = v_19664 | v_19683;
  assign v_19664 = act_19665 & 1'h1;
  assign act_19665 = v_19666 | v_19672;
  assign v_19666 = v_19667 & v_19673;
  assign v_19667 = v_19668 & vout_canPeek_19678;
  assign v_19668 = ~vout_canPeek_19669;
  pebbles_core
    pebbles_core_19669
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19670),
       .in0_consume_en(vin0_consume_en_19669),
       .out_canPeek(vout_canPeek_19669),
       .out_peek(vout_peek_19669));
  assign v_19670 = v_19671 | v_19676;
  assign v_19671 = mux_19671(v_19672);
  assign v_19672 = vout_canPeek_19669 & v_19673;
  assign v_19673 = v_19674 & 1'h1;
  assign v_19674 = v_19675 | 1'h0;
  assign v_19675 = ~v_19662;
  assign v_19676 = mux_19676(v_19677);
  assign v_19677 = ~v_19672;
  pebbles_core
    pebbles_core_19678
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19679),
       .in0_consume_en(vin0_consume_en_19678),
       .out_canPeek(vout_canPeek_19678),
       .out_peek(vout_peek_19678));
  assign v_19679 = v_19680 | v_19681;
  assign v_19680 = mux_19680(v_19666);
  assign v_19681 = mux_19681(v_19682);
  assign v_19682 = ~v_19666;
  assign v_19683 = v_19684 & 1'h1;
  assign v_19684 = v_19685 & v_19686;
  assign v_19685 = ~act_19665;
  assign v_19686 = v_19687 | v_19691;
  assign v_19687 = v_19688 | v_19689;
  assign v_19688 = mux_19688(v_19622);
  assign v_19689 = mux_19689(v_19690);
  assign v_19690 = ~v_19622;
  assign v_19691 = ~v_19662;
  assign v_19692 = v_19693 | v_19694;
  assign v_19693 = mux_19693(v_19664);
  assign v_19694 = mux_19694(v_19683);
  assign v_19695 = v_19696 & 1'h1;
  assign v_19696 = v_19697 & v_19698;
  assign v_19697 = ~act_19621;
  assign v_19698 = v_19699 | v_19707;
  assign v_19699 = v_19700 | v_19705;
  assign v_19700 = mux_19700(v_19701);
  assign v_19701 = v_19618 & v_19702;
  assign v_19702 = v_19703 & 1'h1;
  assign v_19703 = v_19704 | 1'h0;
  assign v_19704 = ~v_19611;
  assign v_19705 = mux_19705(v_19706);
  assign v_19706 = ~v_19701;
  assign v_19707 = ~v_19618;
  assign v_19708 = v_19709 | v_19710;
  assign v_19709 = mux_19709(v_19620);
  assign v_19710 = mux_19710(v_19695);
  assign v_19712 = v_19713 | v_19788;
  assign v_19713 = act_19714 & 1'h1;
  assign act_19714 = v_19715 | v_19745;
  assign v_19715 = v_19716 & v_19746;
  assign v_19716 = v_19717 & v_19755;
  assign v_19717 = ~v_19718;
  assign v_19719 = v_19720 | v_19739;
  assign v_19720 = act_19721 & 1'h1;
  assign act_19721 = v_19722 | v_19728;
  assign v_19722 = v_19723 & v_19729;
  assign v_19723 = v_19724 & vout_canPeek_19734;
  assign v_19724 = ~vout_canPeek_19725;
  pebbles_core
    pebbles_core_19725
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19726),
       .in0_consume_en(vin0_consume_en_19725),
       .out_canPeek(vout_canPeek_19725),
       .out_peek(vout_peek_19725));
  assign v_19726 = v_19727 | v_19732;
  assign v_19727 = mux_19727(v_19728);
  assign v_19728 = vout_canPeek_19725 & v_19729;
  assign v_19729 = v_19730 & 1'h1;
  assign v_19730 = v_19731 | 1'h0;
  assign v_19731 = ~v_19718;
  assign v_19732 = mux_19732(v_19733);
  assign v_19733 = ~v_19728;
  pebbles_core
    pebbles_core_19734
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19735),
       .in0_consume_en(vin0_consume_en_19734),
       .out_canPeek(vout_canPeek_19734),
       .out_peek(vout_peek_19734));
  assign v_19735 = v_19736 | v_19737;
  assign v_19736 = mux_19736(v_19722);
  assign v_19737 = mux_19737(v_19738);
  assign v_19738 = ~v_19722;
  assign v_19739 = v_19740 & 1'h1;
  assign v_19740 = v_19741 & v_19742;
  assign v_19741 = ~act_19721;
  assign v_19742 = v_19743 | v_19751;
  assign v_19743 = v_19744 | v_19749;
  assign v_19744 = mux_19744(v_19745);
  assign v_19745 = v_19718 & v_19746;
  assign v_19746 = v_19747 & 1'h1;
  assign v_19747 = v_19748 | 1'h0;
  assign v_19748 = ~v_19711;
  assign v_19749 = mux_19749(v_19750);
  assign v_19750 = ~v_19745;
  assign v_19751 = ~v_19718;
  assign v_19752 = v_19753 | v_19754;
  assign v_19753 = mux_19753(v_19720);
  assign v_19754 = mux_19754(v_19739);
  assign v_19756 = v_19757 | v_19776;
  assign v_19757 = act_19758 & 1'h1;
  assign act_19758 = v_19759 | v_19765;
  assign v_19759 = v_19760 & v_19766;
  assign v_19760 = v_19761 & vout_canPeek_19771;
  assign v_19761 = ~vout_canPeek_19762;
  pebbles_core
    pebbles_core_19762
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19763),
       .in0_consume_en(vin0_consume_en_19762),
       .out_canPeek(vout_canPeek_19762),
       .out_peek(vout_peek_19762));
  assign v_19763 = v_19764 | v_19769;
  assign v_19764 = mux_19764(v_19765);
  assign v_19765 = vout_canPeek_19762 & v_19766;
  assign v_19766 = v_19767 & 1'h1;
  assign v_19767 = v_19768 | 1'h0;
  assign v_19768 = ~v_19755;
  assign v_19769 = mux_19769(v_19770);
  assign v_19770 = ~v_19765;
  pebbles_core
    pebbles_core_19771
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19772),
       .in0_consume_en(vin0_consume_en_19771),
       .out_canPeek(vout_canPeek_19771),
       .out_peek(vout_peek_19771));
  assign v_19772 = v_19773 | v_19774;
  assign v_19773 = mux_19773(v_19759);
  assign v_19774 = mux_19774(v_19775);
  assign v_19775 = ~v_19759;
  assign v_19776 = v_19777 & 1'h1;
  assign v_19777 = v_19778 & v_19779;
  assign v_19778 = ~act_19758;
  assign v_19779 = v_19780 | v_19784;
  assign v_19780 = v_19781 | v_19782;
  assign v_19781 = mux_19781(v_19715);
  assign v_19782 = mux_19782(v_19783);
  assign v_19783 = ~v_19715;
  assign v_19784 = ~v_19755;
  assign v_19785 = v_19786 | v_19787;
  assign v_19786 = mux_19786(v_19757);
  assign v_19787 = mux_19787(v_19776);
  assign v_19788 = v_19789 & 1'h1;
  assign v_19789 = v_19790 & v_19791;
  assign v_19790 = ~act_19714;
  assign v_19791 = v_19792 | v_19796;
  assign v_19792 = v_19793 | v_19794;
  assign v_19793 = mux_19793(v_19615);
  assign v_19794 = mux_19794(v_19795);
  assign v_19795 = ~v_19615;
  assign v_19796 = ~v_19711;
  assign v_19797 = v_19798 | v_19799;
  assign v_19798 = mux_19798(v_19713);
  assign v_19799 = mux_19799(v_19788);
  assign v_19800 = v_19801 & 1'h1;
  assign v_19801 = v_19802 & v_19803;
  assign v_19802 = ~act_19614;
  assign v_19803 = v_19804 | v_19812;
  assign v_19804 = v_19805 | v_19810;
  assign v_19805 = mux_19805(v_19806);
  assign v_19806 = v_19611 & v_19807;
  assign v_19807 = v_19808 & 1'h1;
  assign v_19808 = v_19809 | 1'h0;
  assign v_19809 = ~v_19604;
  assign v_19810 = mux_19810(v_19811);
  assign v_19811 = ~v_19806;
  assign v_19812 = ~v_19611;
  assign v_19813 = v_19814 | v_19815;
  assign v_19814 = mux_19814(v_19613);
  assign v_19815 = mux_19815(v_19800);
  assign v_19817 = v_19818 | v_20005;
  assign v_19818 = act_19819 & 1'h1;
  assign act_19819 = v_19820 | v_19906;
  assign v_19820 = v_19821 & v_19907;
  assign v_19821 = v_19822 & v_19916;
  assign v_19822 = ~v_19823;
  assign v_19824 = v_19825 | v_19900;
  assign v_19825 = act_19826 & 1'h1;
  assign act_19826 = v_19827 | v_19857;
  assign v_19827 = v_19828 & v_19858;
  assign v_19828 = v_19829 & v_19867;
  assign v_19829 = ~v_19830;
  assign v_19831 = v_19832 | v_19851;
  assign v_19832 = act_19833 & 1'h1;
  assign act_19833 = v_19834 | v_19840;
  assign v_19834 = v_19835 & v_19841;
  assign v_19835 = v_19836 & vout_canPeek_19846;
  assign v_19836 = ~vout_canPeek_19837;
  pebbles_core
    pebbles_core_19837
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19838),
       .in0_consume_en(vin0_consume_en_19837),
       .out_canPeek(vout_canPeek_19837),
       .out_peek(vout_peek_19837));
  assign v_19838 = v_19839 | v_19844;
  assign v_19839 = mux_19839(v_19840);
  assign v_19840 = vout_canPeek_19837 & v_19841;
  assign v_19841 = v_19842 & 1'h1;
  assign v_19842 = v_19843 | 1'h0;
  assign v_19843 = ~v_19830;
  assign v_19844 = mux_19844(v_19845);
  assign v_19845 = ~v_19840;
  pebbles_core
    pebbles_core_19846
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19847),
       .in0_consume_en(vin0_consume_en_19846),
       .out_canPeek(vout_canPeek_19846),
       .out_peek(vout_peek_19846));
  assign v_19847 = v_19848 | v_19849;
  assign v_19848 = mux_19848(v_19834);
  assign v_19849 = mux_19849(v_19850);
  assign v_19850 = ~v_19834;
  assign v_19851 = v_19852 & 1'h1;
  assign v_19852 = v_19853 & v_19854;
  assign v_19853 = ~act_19833;
  assign v_19854 = v_19855 | v_19863;
  assign v_19855 = v_19856 | v_19861;
  assign v_19856 = mux_19856(v_19857);
  assign v_19857 = v_19830 & v_19858;
  assign v_19858 = v_19859 & 1'h1;
  assign v_19859 = v_19860 | 1'h0;
  assign v_19860 = ~v_19823;
  assign v_19861 = mux_19861(v_19862);
  assign v_19862 = ~v_19857;
  assign v_19863 = ~v_19830;
  assign v_19864 = v_19865 | v_19866;
  assign v_19865 = mux_19865(v_19832);
  assign v_19866 = mux_19866(v_19851);
  assign v_19868 = v_19869 | v_19888;
  assign v_19869 = act_19870 & 1'h1;
  assign act_19870 = v_19871 | v_19877;
  assign v_19871 = v_19872 & v_19878;
  assign v_19872 = v_19873 & vout_canPeek_19883;
  assign v_19873 = ~vout_canPeek_19874;
  pebbles_core
    pebbles_core_19874
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19875),
       .in0_consume_en(vin0_consume_en_19874),
       .out_canPeek(vout_canPeek_19874),
       .out_peek(vout_peek_19874));
  assign v_19875 = v_19876 | v_19881;
  assign v_19876 = mux_19876(v_19877);
  assign v_19877 = vout_canPeek_19874 & v_19878;
  assign v_19878 = v_19879 & 1'h1;
  assign v_19879 = v_19880 | 1'h0;
  assign v_19880 = ~v_19867;
  assign v_19881 = mux_19881(v_19882);
  assign v_19882 = ~v_19877;
  pebbles_core
    pebbles_core_19883
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19884),
       .in0_consume_en(vin0_consume_en_19883),
       .out_canPeek(vout_canPeek_19883),
       .out_peek(vout_peek_19883));
  assign v_19884 = v_19885 | v_19886;
  assign v_19885 = mux_19885(v_19871);
  assign v_19886 = mux_19886(v_19887);
  assign v_19887 = ~v_19871;
  assign v_19888 = v_19889 & 1'h1;
  assign v_19889 = v_19890 & v_19891;
  assign v_19890 = ~act_19870;
  assign v_19891 = v_19892 | v_19896;
  assign v_19892 = v_19893 | v_19894;
  assign v_19893 = mux_19893(v_19827);
  assign v_19894 = mux_19894(v_19895);
  assign v_19895 = ~v_19827;
  assign v_19896 = ~v_19867;
  assign v_19897 = v_19898 | v_19899;
  assign v_19898 = mux_19898(v_19869);
  assign v_19899 = mux_19899(v_19888);
  assign v_19900 = v_19901 & 1'h1;
  assign v_19901 = v_19902 & v_19903;
  assign v_19902 = ~act_19826;
  assign v_19903 = v_19904 | v_19912;
  assign v_19904 = v_19905 | v_19910;
  assign v_19905 = mux_19905(v_19906);
  assign v_19906 = v_19823 & v_19907;
  assign v_19907 = v_19908 & 1'h1;
  assign v_19908 = v_19909 | 1'h0;
  assign v_19909 = ~v_19816;
  assign v_19910 = mux_19910(v_19911);
  assign v_19911 = ~v_19906;
  assign v_19912 = ~v_19823;
  assign v_19913 = v_19914 | v_19915;
  assign v_19914 = mux_19914(v_19825);
  assign v_19915 = mux_19915(v_19900);
  assign v_19917 = v_19918 | v_19993;
  assign v_19918 = act_19919 & 1'h1;
  assign act_19919 = v_19920 | v_19950;
  assign v_19920 = v_19921 & v_19951;
  assign v_19921 = v_19922 & v_19960;
  assign v_19922 = ~v_19923;
  assign v_19924 = v_19925 | v_19944;
  assign v_19925 = act_19926 & 1'h1;
  assign act_19926 = v_19927 | v_19933;
  assign v_19927 = v_19928 & v_19934;
  assign v_19928 = v_19929 & vout_canPeek_19939;
  assign v_19929 = ~vout_canPeek_19930;
  pebbles_core
    pebbles_core_19930
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19931),
       .in0_consume_en(vin0_consume_en_19930),
       .out_canPeek(vout_canPeek_19930),
       .out_peek(vout_peek_19930));
  assign v_19931 = v_19932 | v_19937;
  assign v_19932 = mux_19932(v_19933);
  assign v_19933 = vout_canPeek_19930 & v_19934;
  assign v_19934 = v_19935 & 1'h1;
  assign v_19935 = v_19936 | 1'h0;
  assign v_19936 = ~v_19923;
  assign v_19937 = mux_19937(v_19938);
  assign v_19938 = ~v_19933;
  pebbles_core
    pebbles_core_19939
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19940),
       .in0_consume_en(vin0_consume_en_19939),
       .out_canPeek(vout_canPeek_19939),
       .out_peek(vout_peek_19939));
  assign v_19940 = v_19941 | v_19942;
  assign v_19941 = mux_19941(v_19927);
  assign v_19942 = mux_19942(v_19943);
  assign v_19943 = ~v_19927;
  assign v_19944 = v_19945 & 1'h1;
  assign v_19945 = v_19946 & v_19947;
  assign v_19946 = ~act_19926;
  assign v_19947 = v_19948 | v_19956;
  assign v_19948 = v_19949 | v_19954;
  assign v_19949 = mux_19949(v_19950);
  assign v_19950 = v_19923 & v_19951;
  assign v_19951 = v_19952 & 1'h1;
  assign v_19952 = v_19953 | 1'h0;
  assign v_19953 = ~v_19916;
  assign v_19954 = mux_19954(v_19955);
  assign v_19955 = ~v_19950;
  assign v_19956 = ~v_19923;
  assign v_19957 = v_19958 | v_19959;
  assign v_19958 = mux_19958(v_19925);
  assign v_19959 = mux_19959(v_19944);
  assign v_19961 = v_19962 | v_19981;
  assign v_19962 = act_19963 & 1'h1;
  assign act_19963 = v_19964 | v_19970;
  assign v_19964 = v_19965 & v_19971;
  assign v_19965 = v_19966 & vout_canPeek_19976;
  assign v_19966 = ~vout_canPeek_19967;
  pebbles_core
    pebbles_core_19967
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19968),
       .in0_consume_en(vin0_consume_en_19967),
       .out_canPeek(vout_canPeek_19967),
       .out_peek(vout_peek_19967));
  assign v_19968 = v_19969 | v_19974;
  assign v_19969 = mux_19969(v_19970);
  assign v_19970 = vout_canPeek_19967 & v_19971;
  assign v_19971 = v_19972 & 1'h1;
  assign v_19972 = v_19973 | 1'h0;
  assign v_19973 = ~v_19960;
  assign v_19974 = mux_19974(v_19975);
  assign v_19975 = ~v_19970;
  pebbles_core
    pebbles_core_19976
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_19977),
       .in0_consume_en(vin0_consume_en_19976),
       .out_canPeek(vout_canPeek_19976),
       .out_peek(vout_peek_19976));
  assign v_19977 = v_19978 | v_19979;
  assign v_19978 = mux_19978(v_19964);
  assign v_19979 = mux_19979(v_19980);
  assign v_19980 = ~v_19964;
  assign v_19981 = v_19982 & 1'h1;
  assign v_19982 = v_19983 & v_19984;
  assign v_19983 = ~act_19963;
  assign v_19984 = v_19985 | v_19989;
  assign v_19985 = v_19986 | v_19987;
  assign v_19986 = mux_19986(v_19920);
  assign v_19987 = mux_19987(v_19988);
  assign v_19988 = ~v_19920;
  assign v_19989 = ~v_19960;
  assign v_19990 = v_19991 | v_19992;
  assign v_19991 = mux_19991(v_19962);
  assign v_19992 = mux_19992(v_19981);
  assign v_19993 = v_19994 & 1'h1;
  assign v_19994 = v_19995 & v_19996;
  assign v_19995 = ~act_19919;
  assign v_19996 = v_19997 | v_20001;
  assign v_19997 = v_19998 | v_19999;
  assign v_19998 = mux_19998(v_19820);
  assign v_19999 = mux_19999(v_20000);
  assign v_20000 = ~v_19820;
  assign v_20001 = ~v_19916;
  assign v_20002 = v_20003 | v_20004;
  assign v_20003 = mux_20003(v_19918);
  assign v_20004 = mux_20004(v_19993);
  assign v_20005 = v_20006 & 1'h1;
  assign v_20006 = v_20007 & v_20008;
  assign v_20007 = ~act_19819;
  assign v_20008 = v_20009 | v_20013;
  assign v_20009 = v_20010 | v_20011;
  assign v_20010 = mux_20010(v_19608);
  assign v_20011 = mux_20011(v_20012);
  assign v_20012 = ~v_19608;
  assign v_20013 = ~v_19816;
  assign v_20014 = v_20015 | v_20016;
  assign v_20015 = mux_20015(v_19818);
  assign v_20016 = mux_20016(v_20005);
  assign v_20017 = v_20018 & 1'h1;
  assign v_20018 = v_20019 & v_20020;
  assign v_20019 = ~act_19607;
  assign v_20020 = v_20021 | v_20029;
  assign v_20021 = v_20022 | v_20027;
  assign v_20022 = mux_20022(v_20023);
  assign v_20023 = v_19604 & v_20024;
  assign v_20024 = v_20025 & 1'h1;
  assign v_20025 = v_20026 | 1'h0;
  assign v_20026 = ~v_19597;
  assign v_20027 = mux_20027(v_20028);
  assign v_20028 = ~v_20023;
  assign v_20029 = ~v_19604;
  assign v_20030 = v_20031 | v_20032;
  assign v_20031 = mux_20031(v_19606);
  assign v_20032 = mux_20032(v_20017);
  assign v_20034 = v_20035 | v_20446;
  assign v_20035 = act_20036 & 1'h1;
  assign act_20036 = v_20037 | v_20235;
  assign v_20037 = v_20038 & v_20236;
  assign v_20038 = v_20039 & v_20245;
  assign v_20039 = ~v_20040;
  assign v_20041 = v_20042 | v_20229;
  assign v_20042 = act_20043 & 1'h1;
  assign act_20043 = v_20044 | v_20130;
  assign v_20044 = v_20045 & v_20131;
  assign v_20045 = v_20046 & v_20140;
  assign v_20046 = ~v_20047;
  assign v_20048 = v_20049 | v_20124;
  assign v_20049 = act_20050 & 1'h1;
  assign act_20050 = v_20051 | v_20081;
  assign v_20051 = v_20052 & v_20082;
  assign v_20052 = v_20053 & v_20091;
  assign v_20053 = ~v_20054;
  assign v_20055 = v_20056 | v_20075;
  assign v_20056 = act_20057 & 1'h1;
  assign act_20057 = v_20058 | v_20064;
  assign v_20058 = v_20059 & v_20065;
  assign v_20059 = v_20060 & vout_canPeek_20070;
  assign v_20060 = ~vout_canPeek_20061;
  pebbles_core
    pebbles_core_20061
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20062),
       .in0_consume_en(vin0_consume_en_20061),
       .out_canPeek(vout_canPeek_20061),
       .out_peek(vout_peek_20061));
  assign v_20062 = v_20063 | v_20068;
  assign v_20063 = mux_20063(v_20064);
  assign v_20064 = vout_canPeek_20061 & v_20065;
  assign v_20065 = v_20066 & 1'h1;
  assign v_20066 = v_20067 | 1'h0;
  assign v_20067 = ~v_20054;
  assign v_20068 = mux_20068(v_20069);
  assign v_20069 = ~v_20064;
  pebbles_core
    pebbles_core_20070
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20071),
       .in0_consume_en(vin0_consume_en_20070),
       .out_canPeek(vout_canPeek_20070),
       .out_peek(vout_peek_20070));
  assign v_20071 = v_20072 | v_20073;
  assign v_20072 = mux_20072(v_20058);
  assign v_20073 = mux_20073(v_20074);
  assign v_20074 = ~v_20058;
  assign v_20075 = v_20076 & 1'h1;
  assign v_20076 = v_20077 & v_20078;
  assign v_20077 = ~act_20057;
  assign v_20078 = v_20079 | v_20087;
  assign v_20079 = v_20080 | v_20085;
  assign v_20080 = mux_20080(v_20081);
  assign v_20081 = v_20054 & v_20082;
  assign v_20082 = v_20083 & 1'h1;
  assign v_20083 = v_20084 | 1'h0;
  assign v_20084 = ~v_20047;
  assign v_20085 = mux_20085(v_20086);
  assign v_20086 = ~v_20081;
  assign v_20087 = ~v_20054;
  assign v_20088 = v_20089 | v_20090;
  assign v_20089 = mux_20089(v_20056);
  assign v_20090 = mux_20090(v_20075);
  assign v_20092 = v_20093 | v_20112;
  assign v_20093 = act_20094 & 1'h1;
  assign act_20094 = v_20095 | v_20101;
  assign v_20095 = v_20096 & v_20102;
  assign v_20096 = v_20097 & vout_canPeek_20107;
  assign v_20097 = ~vout_canPeek_20098;
  pebbles_core
    pebbles_core_20098
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20099),
       .in0_consume_en(vin0_consume_en_20098),
       .out_canPeek(vout_canPeek_20098),
       .out_peek(vout_peek_20098));
  assign v_20099 = v_20100 | v_20105;
  assign v_20100 = mux_20100(v_20101);
  assign v_20101 = vout_canPeek_20098 & v_20102;
  assign v_20102 = v_20103 & 1'h1;
  assign v_20103 = v_20104 | 1'h0;
  assign v_20104 = ~v_20091;
  assign v_20105 = mux_20105(v_20106);
  assign v_20106 = ~v_20101;
  pebbles_core
    pebbles_core_20107
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20108),
       .in0_consume_en(vin0_consume_en_20107),
       .out_canPeek(vout_canPeek_20107),
       .out_peek(vout_peek_20107));
  assign v_20108 = v_20109 | v_20110;
  assign v_20109 = mux_20109(v_20095);
  assign v_20110 = mux_20110(v_20111);
  assign v_20111 = ~v_20095;
  assign v_20112 = v_20113 & 1'h1;
  assign v_20113 = v_20114 & v_20115;
  assign v_20114 = ~act_20094;
  assign v_20115 = v_20116 | v_20120;
  assign v_20116 = v_20117 | v_20118;
  assign v_20117 = mux_20117(v_20051);
  assign v_20118 = mux_20118(v_20119);
  assign v_20119 = ~v_20051;
  assign v_20120 = ~v_20091;
  assign v_20121 = v_20122 | v_20123;
  assign v_20122 = mux_20122(v_20093);
  assign v_20123 = mux_20123(v_20112);
  assign v_20124 = v_20125 & 1'h1;
  assign v_20125 = v_20126 & v_20127;
  assign v_20126 = ~act_20050;
  assign v_20127 = v_20128 | v_20136;
  assign v_20128 = v_20129 | v_20134;
  assign v_20129 = mux_20129(v_20130);
  assign v_20130 = v_20047 & v_20131;
  assign v_20131 = v_20132 & 1'h1;
  assign v_20132 = v_20133 | 1'h0;
  assign v_20133 = ~v_20040;
  assign v_20134 = mux_20134(v_20135);
  assign v_20135 = ~v_20130;
  assign v_20136 = ~v_20047;
  assign v_20137 = v_20138 | v_20139;
  assign v_20138 = mux_20138(v_20049);
  assign v_20139 = mux_20139(v_20124);
  assign v_20141 = v_20142 | v_20217;
  assign v_20142 = act_20143 & 1'h1;
  assign act_20143 = v_20144 | v_20174;
  assign v_20144 = v_20145 & v_20175;
  assign v_20145 = v_20146 & v_20184;
  assign v_20146 = ~v_20147;
  assign v_20148 = v_20149 | v_20168;
  assign v_20149 = act_20150 & 1'h1;
  assign act_20150 = v_20151 | v_20157;
  assign v_20151 = v_20152 & v_20158;
  assign v_20152 = v_20153 & vout_canPeek_20163;
  assign v_20153 = ~vout_canPeek_20154;
  pebbles_core
    pebbles_core_20154
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20155),
       .in0_consume_en(vin0_consume_en_20154),
       .out_canPeek(vout_canPeek_20154),
       .out_peek(vout_peek_20154));
  assign v_20155 = v_20156 | v_20161;
  assign v_20156 = mux_20156(v_20157);
  assign v_20157 = vout_canPeek_20154 & v_20158;
  assign v_20158 = v_20159 & 1'h1;
  assign v_20159 = v_20160 | 1'h0;
  assign v_20160 = ~v_20147;
  assign v_20161 = mux_20161(v_20162);
  assign v_20162 = ~v_20157;
  pebbles_core
    pebbles_core_20163
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20164),
       .in0_consume_en(vin0_consume_en_20163),
       .out_canPeek(vout_canPeek_20163),
       .out_peek(vout_peek_20163));
  assign v_20164 = v_20165 | v_20166;
  assign v_20165 = mux_20165(v_20151);
  assign v_20166 = mux_20166(v_20167);
  assign v_20167 = ~v_20151;
  assign v_20168 = v_20169 & 1'h1;
  assign v_20169 = v_20170 & v_20171;
  assign v_20170 = ~act_20150;
  assign v_20171 = v_20172 | v_20180;
  assign v_20172 = v_20173 | v_20178;
  assign v_20173 = mux_20173(v_20174);
  assign v_20174 = v_20147 & v_20175;
  assign v_20175 = v_20176 & 1'h1;
  assign v_20176 = v_20177 | 1'h0;
  assign v_20177 = ~v_20140;
  assign v_20178 = mux_20178(v_20179);
  assign v_20179 = ~v_20174;
  assign v_20180 = ~v_20147;
  assign v_20181 = v_20182 | v_20183;
  assign v_20182 = mux_20182(v_20149);
  assign v_20183 = mux_20183(v_20168);
  assign v_20185 = v_20186 | v_20205;
  assign v_20186 = act_20187 & 1'h1;
  assign act_20187 = v_20188 | v_20194;
  assign v_20188 = v_20189 & v_20195;
  assign v_20189 = v_20190 & vout_canPeek_20200;
  assign v_20190 = ~vout_canPeek_20191;
  pebbles_core
    pebbles_core_20191
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20192),
       .in0_consume_en(vin0_consume_en_20191),
       .out_canPeek(vout_canPeek_20191),
       .out_peek(vout_peek_20191));
  assign v_20192 = v_20193 | v_20198;
  assign v_20193 = mux_20193(v_20194);
  assign v_20194 = vout_canPeek_20191 & v_20195;
  assign v_20195 = v_20196 & 1'h1;
  assign v_20196 = v_20197 | 1'h0;
  assign v_20197 = ~v_20184;
  assign v_20198 = mux_20198(v_20199);
  assign v_20199 = ~v_20194;
  pebbles_core
    pebbles_core_20200
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20201),
       .in0_consume_en(vin0_consume_en_20200),
       .out_canPeek(vout_canPeek_20200),
       .out_peek(vout_peek_20200));
  assign v_20201 = v_20202 | v_20203;
  assign v_20202 = mux_20202(v_20188);
  assign v_20203 = mux_20203(v_20204);
  assign v_20204 = ~v_20188;
  assign v_20205 = v_20206 & 1'h1;
  assign v_20206 = v_20207 & v_20208;
  assign v_20207 = ~act_20187;
  assign v_20208 = v_20209 | v_20213;
  assign v_20209 = v_20210 | v_20211;
  assign v_20210 = mux_20210(v_20144);
  assign v_20211 = mux_20211(v_20212);
  assign v_20212 = ~v_20144;
  assign v_20213 = ~v_20184;
  assign v_20214 = v_20215 | v_20216;
  assign v_20215 = mux_20215(v_20186);
  assign v_20216 = mux_20216(v_20205);
  assign v_20217 = v_20218 & 1'h1;
  assign v_20218 = v_20219 & v_20220;
  assign v_20219 = ~act_20143;
  assign v_20220 = v_20221 | v_20225;
  assign v_20221 = v_20222 | v_20223;
  assign v_20222 = mux_20222(v_20044);
  assign v_20223 = mux_20223(v_20224);
  assign v_20224 = ~v_20044;
  assign v_20225 = ~v_20140;
  assign v_20226 = v_20227 | v_20228;
  assign v_20227 = mux_20227(v_20142);
  assign v_20228 = mux_20228(v_20217);
  assign v_20229 = v_20230 & 1'h1;
  assign v_20230 = v_20231 & v_20232;
  assign v_20231 = ~act_20043;
  assign v_20232 = v_20233 | v_20241;
  assign v_20233 = v_20234 | v_20239;
  assign v_20234 = mux_20234(v_20235);
  assign v_20235 = v_20040 & v_20236;
  assign v_20236 = v_20237 & 1'h1;
  assign v_20237 = v_20238 | 1'h0;
  assign v_20238 = ~v_20033;
  assign v_20239 = mux_20239(v_20240);
  assign v_20240 = ~v_20235;
  assign v_20241 = ~v_20040;
  assign v_20242 = v_20243 | v_20244;
  assign v_20243 = mux_20243(v_20042);
  assign v_20244 = mux_20244(v_20229);
  assign v_20246 = v_20247 | v_20434;
  assign v_20247 = act_20248 & 1'h1;
  assign act_20248 = v_20249 | v_20335;
  assign v_20249 = v_20250 & v_20336;
  assign v_20250 = v_20251 & v_20345;
  assign v_20251 = ~v_20252;
  assign v_20253 = v_20254 | v_20329;
  assign v_20254 = act_20255 & 1'h1;
  assign act_20255 = v_20256 | v_20286;
  assign v_20256 = v_20257 & v_20287;
  assign v_20257 = v_20258 & v_20296;
  assign v_20258 = ~v_20259;
  assign v_20260 = v_20261 | v_20280;
  assign v_20261 = act_20262 & 1'h1;
  assign act_20262 = v_20263 | v_20269;
  assign v_20263 = v_20264 & v_20270;
  assign v_20264 = v_20265 & vout_canPeek_20275;
  assign v_20265 = ~vout_canPeek_20266;
  pebbles_core
    pebbles_core_20266
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20267),
       .in0_consume_en(vin0_consume_en_20266),
       .out_canPeek(vout_canPeek_20266),
       .out_peek(vout_peek_20266));
  assign v_20267 = v_20268 | v_20273;
  assign v_20268 = mux_20268(v_20269);
  assign v_20269 = vout_canPeek_20266 & v_20270;
  assign v_20270 = v_20271 & 1'h1;
  assign v_20271 = v_20272 | 1'h0;
  assign v_20272 = ~v_20259;
  assign v_20273 = mux_20273(v_20274);
  assign v_20274 = ~v_20269;
  pebbles_core
    pebbles_core_20275
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20276),
       .in0_consume_en(vin0_consume_en_20275),
       .out_canPeek(vout_canPeek_20275),
       .out_peek(vout_peek_20275));
  assign v_20276 = v_20277 | v_20278;
  assign v_20277 = mux_20277(v_20263);
  assign v_20278 = mux_20278(v_20279);
  assign v_20279 = ~v_20263;
  assign v_20280 = v_20281 & 1'h1;
  assign v_20281 = v_20282 & v_20283;
  assign v_20282 = ~act_20262;
  assign v_20283 = v_20284 | v_20292;
  assign v_20284 = v_20285 | v_20290;
  assign v_20285 = mux_20285(v_20286);
  assign v_20286 = v_20259 & v_20287;
  assign v_20287 = v_20288 & 1'h1;
  assign v_20288 = v_20289 | 1'h0;
  assign v_20289 = ~v_20252;
  assign v_20290 = mux_20290(v_20291);
  assign v_20291 = ~v_20286;
  assign v_20292 = ~v_20259;
  assign v_20293 = v_20294 | v_20295;
  assign v_20294 = mux_20294(v_20261);
  assign v_20295 = mux_20295(v_20280);
  assign v_20297 = v_20298 | v_20317;
  assign v_20298 = act_20299 & 1'h1;
  assign act_20299 = v_20300 | v_20306;
  assign v_20300 = v_20301 & v_20307;
  assign v_20301 = v_20302 & vout_canPeek_20312;
  assign v_20302 = ~vout_canPeek_20303;
  pebbles_core
    pebbles_core_20303
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20304),
       .in0_consume_en(vin0_consume_en_20303),
       .out_canPeek(vout_canPeek_20303),
       .out_peek(vout_peek_20303));
  assign v_20304 = v_20305 | v_20310;
  assign v_20305 = mux_20305(v_20306);
  assign v_20306 = vout_canPeek_20303 & v_20307;
  assign v_20307 = v_20308 & 1'h1;
  assign v_20308 = v_20309 | 1'h0;
  assign v_20309 = ~v_20296;
  assign v_20310 = mux_20310(v_20311);
  assign v_20311 = ~v_20306;
  pebbles_core
    pebbles_core_20312
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20313),
       .in0_consume_en(vin0_consume_en_20312),
       .out_canPeek(vout_canPeek_20312),
       .out_peek(vout_peek_20312));
  assign v_20313 = v_20314 | v_20315;
  assign v_20314 = mux_20314(v_20300);
  assign v_20315 = mux_20315(v_20316);
  assign v_20316 = ~v_20300;
  assign v_20317 = v_20318 & 1'h1;
  assign v_20318 = v_20319 & v_20320;
  assign v_20319 = ~act_20299;
  assign v_20320 = v_20321 | v_20325;
  assign v_20321 = v_20322 | v_20323;
  assign v_20322 = mux_20322(v_20256);
  assign v_20323 = mux_20323(v_20324);
  assign v_20324 = ~v_20256;
  assign v_20325 = ~v_20296;
  assign v_20326 = v_20327 | v_20328;
  assign v_20327 = mux_20327(v_20298);
  assign v_20328 = mux_20328(v_20317);
  assign v_20329 = v_20330 & 1'h1;
  assign v_20330 = v_20331 & v_20332;
  assign v_20331 = ~act_20255;
  assign v_20332 = v_20333 | v_20341;
  assign v_20333 = v_20334 | v_20339;
  assign v_20334 = mux_20334(v_20335);
  assign v_20335 = v_20252 & v_20336;
  assign v_20336 = v_20337 & 1'h1;
  assign v_20337 = v_20338 | 1'h0;
  assign v_20338 = ~v_20245;
  assign v_20339 = mux_20339(v_20340);
  assign v_20340 = ~v_20335;
  assign v_20341 = ~v_20252;
  assign v_20342 = v_20343 | v_20344;
  assign v_20343 = mux_20343(v_20254);
  assign v_20344 = mux_20344(v_20329);
  assign v_20346 = v_20347 | v_20422;
  assign v_20347 = act_20348 & 1'h1;
  assign act_20348 = v_20349 | v_20379;
  assign v_20349 = v_20350 & v_20380;
  assign v_20350 = v_20351 & v_20389;
  assign v_20351 = ~v_20352;
  assign v_20353 = v_20354 | v_20373;
  assign v_20354 = act_20355 & 1'h1;
  assign act_20355 = v_20356 | v_20362;
  assign v_20356 = v_20357 & v_20363;
  assign v_20357 = v_20358 & vout_canPeek_20368;
  assign v_20358 = ~vout_canPeek_20359;
  pebbles_core
    pebbles_core_20359
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20360),
       .in0_consume_en(vin0_consume_en_20359),
       .out_canPeek(vout_canPeek_20359),
       .out_peek(vout_peek_20359));
  assign v_20360 = v_20361 | v_20366;
  assign v_20361 = mux_20361(v_20362);
  assign v_20362 = vout_canPeek_20359 & v_20363;
  assign v_20363 = v_20364 & 1'h1;
  assign v_20364 = v_20365 | 1'h0;
  assign v_20365 = ~v_20352;
  assign v_20366 = mux_20366(v_20367);
  assign v_20367 = ~v_20362;
  pebbles_core
    pebbles_core_20368
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20369),
       .in0_consume_en(vin0_consume_en_20368),
       .out_canPeek(vout_canPeek_20368),
       .out_peek(vout_peek_20368));
  assign v_20369 = v_20370 | v_20371;
  assign v_20370 = mux_20370(v_20356);
  assign v_20371 = mux_20371(v_20372);
  assign v_20372 = ~v_20356;
  assign v_20373 = v_20374 & 1'h1;
  assign v_20374 = v_20375 & v_20376;
  assign v_20375 = ~act_20355;
  assign v_20376 = v_20377 | v_20385;
  assign v_20377 = v_20378 | v_20383;
  assign v_20378 = mux_20378(v_20379);
  assign v_20379 = v_20352 & v_20380;
  assign v_20380 = v_20381 & 1'h1;
  assign v_20381 = v_20382 | 1'h0;
  assign v_20382 = ~v_20345;
  assign v_20383 = mux_20383(v_20384);
  assign v_20384 = ~v_20379;
  assign v_20385 = ~v_20352;
  assign v_20386 = v_20387 | v_20388;
  assign v_20387 = mux_20387(v_20354);
  assign v_20388 = mux_20388(v_20373);
  assign v_20390 = v_20391 | v_20410;
  assign v_20391 = act_20392 & 1'h1;
  assign act_20392 = v_20393 | v_20399;
  assign v_20393 = v_20394 & v_20400;
  assign v_20394 = v_20395 & vout_canPeek_20405;
  assign v_20395 = ~vout_canPeek_20396;
  pebbles_core
    pebbles_core_20396
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20397),
       .in0_consume_en(vin0_consume_en_20396),
       .out_canPeek(vout_canPeek_20396),
       .out_peek(vout_peek_20396));
  assign v_20397 = v_20398 | v_20403;
  assign v_20398 = mux_20398(v_20399);
  assign v_20399 = vout_canPeek_20396 & v_20400;
  assign v_20400 = v_20401 & 1'h1;
  assign v_20401 = v_20402 | 1'h0;
  assign v_20402 = ~v_20389;
  assign v_20403 = mux_20403(v_20404);
  assign v_20404 = ~v_20399;
  pebbles_core
    pebbles_core_20405
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20406),
       .in0_consume_en(vin0_consume_en_20405),
       .out_canPeek(vout_canPeek_20405),
       .out_peek(vout_peek_20405));
  assign v_20406 = v_20407 | v_20408;
  assign v_20407 = mux_20407(v_20393);
  assign v_20408 = mux_20408(v_20409);
  assign v_20409 = ~v_20393;
  assign v_20410 = v_20411 & 1'h1;
  assign v_20411 = v_20412 & v_20413;
  assign v_20412 = ~act_20392;
  assign v_20413 = v_20414 | v_20418;
  assign v_20414 = v_20415 | v_20416;
  assign v_20415 = mux_20415(v_20349);
  assign v_20416 = mux_20416(v_20417);
  assign v_20417 = ~v_20349;
  assign v_20418 = ~v_20389;
  assign v_20419 = v_20420 | v_20421;
  assign v_20420 = mux_20420(v_20391);
  assign v_20421 = mux_20421(v_20410);
  assign v_20422 = v_20423 & 1'h1;
  assign v_20423 = v_20424 & v_20425;
  assign v_20424 = ~act_20348;
  assign v_20425 = v_20426 | v_20430;
  assign v_20426 = v_20427 | v_20428;
  assign v_20427 = mux_20427(v_20249);
  assign v_20428 = mux_20428(v_20429);
  assign v_20429 = ~v_20249;
  assign v_20430 = ~v_20345;
  assign v_20431 = v_20432 | v_20433;
  assign v_20432 = mux_20432(v_20347);
  assign v_20433 = mux_20433(v_20422);
  assign v_20434 = v_20435 & 1'h1;
  assign v_20435 = v_20436 & v_20437;
  assign v_20436 = ~act_20248;
  assign v_20437 = v_20438 | v_20442;
  assign v_20438 = v_20439 | v_20440;
  assign v_20439 = mux_20439(v_20037);
  assign v_20440 = mux_20440(v_20441);
  assign v_20441 = ~v_20037;
  assign v_20442 = ~v_20245;
  assign v_20443 = v_20444 | v_20445;
  assign v_20444 = mux_20444(v_20247);
  assign v_20445 = mux_20445(v_20434);
  assign v_20446 = v_20447 & 1'h1;
  assign v_20447 = v_20448 & v_20449;
  assign v_20448 = ~act_20036;
  assign v_20449 = v_20450 | v_20454;
  assign v_20450 = v_20451 | v_20452;
  assign v_20451 = mux_20451(v_19601);
  assign v_20452 = mux_20452(v_20453);
  assign v_20453 = ~v_19601;
  assign v_20454 = ~v_20033;
  assign v_20455 = v_20456 | v_20457;
  assign v_20456 = mux_20456(v_20035);
  assign v_20457 = mux_20457(v_20446);
  assign v_20458 = v_20459 & 1'h1;
  assign v_20459 = v_20460 & v_20461;
  assign v_20460 = ~act_19600;
  assign v_20461 = v_20462 | v_20466;
  assign v_20462 = v_20463 | v_20464;
  assign v_20463 = mux_20463(v_18717);
  assign v_20464 = mux_20464(v_20465);
  assign v_20465 = ~v_18717;
  assign v_20466 = ~v_19597;
  assign v_20467 = v_20468 | v_20469;
  assign v_20468 = mux_20468(v_19599);
  assign v_20469 = mux_20469(v_20458);
  assign v_20470 = v_20471 & 1'h1;
  assign v_20471 = v_20472 & v_20473;
  assign v_20472 = ~act_18716;
  assign v_20473 = v_20474 | v_20482;
  assign v_20474 = v_20475 | v_20480;
  assign v_20475 = mux_20475(v_20476);
  assign v_20476 = v_18713 & v_20477;
  assign v_20477 = v_20478 & 1'h1;
  assign v_20478 = v_20479 | 1'h0;
  assign v_20479 = ~v_18706;
  assign v_20480 = mux_20480(v_20481);
  assign v_20481 = ~v_20476;
  assign v_20482 = ~v_18713;
  assign v_20483 = v_20484 | v_20485;
  assign v_20484 = mux_20484(v_18715);
  assign v_20485 = mux_20485(v_20470);
  assign v_20487 = v_20488 | v_22243;
  assign v_20488 = act_20489 & 1'h1;
  assign act_20489 = v_20490 | v_21360;
  assign v_20490 = v_20491 & v_21361;
  assign v_20491 = v_20492 & v_21370;
  assign v_20492 = ~v_20493;
  assign v_20494 = v_20495 | v_21354;
  assign v_20495 = act_20496 & 1'h1;
  assign act_20496 = v_20497 | v_20919;
  assign v_20497 = v_20498 & v_20920;
  assign v_20498 = v_20499 & v_20929;
  assign v_20499 = ~v_20500;
  assign v_20501 = v_20502 | v_20913;
  assign v_20502 = act_20503 & 1'h1;
  assign act_20503 = v_20504 | v_20702;
  assign v_20504 = v_20505 & v_20703;
  assign v_20505 = v_20506 & v_20712;
  assign v_20506 = ~v_20507;
  assign v_20508 = v_20509 | v_20696;
  assign v_20509 = act_20510 & 1'h1;
  assign act_20510 = v_20511 | v_20597;
  assign v_20511 = v_20512 & v_20598;
  assign v_20512 = v_20513 & v_20607;
  assign v_20513 = ~v_20514;
  assign v_20515 = v_20516 | v_20591;
  assign v_20516 = act_20517 & 1'h1;
  assign act_20517 = v_20518 | v_20548;
  assign v_20518 = v_20519 & v_20549;
  assign v_20519 = v_20520 & v_20558;
  assign v_20520 = ~v_20521;
  assign v_20522 = v_20523 | v_20542;
  assign v_20523 = act_20524 & 1'h1;
  assign act_20524 = v_20525 | v_20531;
  assign v_20525 = v_20526 & v_20532;
  assign v_20526 = v_20527 & vout_canPeek_20537;
  assign v_20527 = ~vout_canPeek_20528;
  pebbles_core
    pebbles_core_20528
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20529),
       .in0_consume_en(vin0_consume_en_20528),
       .out_canPeek(vout_canPeek_20528),
       .out_peek(vout_peek_20528));
  assign v_20529 = v_20530 | v_20535;
  assign v_20530 = mux_20530(v_20531);
  assign v_20531 = vout_canPeek_20528 & v_20532;
  assign v_20532 = v_20533 & 1'h1;
  assign v_20533 = v_20534 | 1'h0;
  assign v_20534 = ~v_20521;
  assign v_20535 = mux_20535(v_20536);
  assign v_20536 = ~v_20531;
  pebbles_core
    pebbles_core_20537
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20538),
       .in0_consume_en(vin0_consume_en_20537),
       .out_canPeek(vout_canPeek_20537),
       .out_peek(vout_peek_20537));
  assign v_20538 = v_20539 | v_20540;
  assign v_20539 = mux_20539(v_20525);
  assign v_20540 = mux_20540(v_20541);
  assign v_20541 = ~v_20525;
  assign v_20542 = v_20543 & 1'h1;
  assign v_20543 = v_20544 & v_20545;
  assign v_20544 = ~act_20524;
  assign v_20545 = v_20546 | v_20554;
  assign v_20546 = v_20547 | v_20552;
  assign v_20547 = mux_20547(v_20548);
  assign v_20548 = v_20521 & v_20549;
  assign v_20549 = v_20550 & 1'h1;
  assign v_20550 = v_20551 | 1'h0;
  assign v_20551 = ~v_20514;
  assign v_20552 = mux_20552(v_20553);
  assign v_20553 = ~v_20548;
  assign v_20554 = ~v_20521;
  assign v_20555 = v_20556 | v_20557;
  assign v_20556 = mux_20556(v_20523);
  assign v_20557 = mux_20557(v_20542);
  assign v_20559 = v_20560 | v_20579;
  assign v_20560 = act_20561 & 1'h1;
  assign act_20561 = v_20562 | v_20568;
  assign v_20562 = v_20563 & v_20569;
  assign v_20563 = v_20564 & vout_canPeek_20574;
  assign v_20564 = ~vout_canPeek_20565;
  pebbles_core
    pebbles_core_20565
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20566),
       .in0_consume_en(vin0_consume_en_20565),
       .out_canPeek(vout_canPeek_20565),
       .out_peek(vout_peek_20565));
  assign v_20566 = v_20567 | v_20572;
  assign v_20567 = mux_20567(v_20568);
  assign v_20568 = vout_canPeek_20565 & v_20569;
  assign v_20569 = v_20570 & 1'h1;
  assign v_20570 = v_20571 | 1'h0;
  assign v_20571 = ~v_20558;
  assign v_20572 = mux_20572(v_20573);
  assign v_20573 = ~v_20568;
  pebbles_core
    pebbles_core_20574
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20575),
       .in0_consume_en(vin0_consume_en_20574),
       .out_canPeek(vout_canPeek_20574),
       .out_peek(vout_peek_20574));
  assign v_20575 = v_20576 | v_20577;
  assign v_20576 = mux_20576(v_20562);
  assign v_20577 = mux_20577(v_20578);
  assign v_20578 = ~v_20562;
  assign v_20579 = v_20580 & 1'h1;
  assign v_20580 = v_20581 & v_20582;
  assign v_20581 = ~act_20561;
  assign v_20582 = v_20583 | v_20587;
  assign v_20583 = v_20584 | v_20585;
  assign v_20584 = mux_20584(v_20518);
  assign v_20585 = mux_20585(v_20586);
  assign v_20586 = ~v_20518;
  assign v_20587 = ~v_20558;
  assign v_20588 = v_20589 | v_20590;
  assign v_20589 = mux_20589(v_20560);
  assign v_20590 = mux_20590(v_20579);
  assign v_20591 = v_20592 & 1'h1;
  assign v_20592 = v_20593 & v_20594;
  assign v_20593 = ~act_20517;
  assign v_20594 = v_20595 | v_20603;
  assign v_20595 = v_20596 | v_20601;
  assign v_20596 = mux_20596(v_20597);
  assign v_20597 = v_20514 & v_20598;
  assign v_20598 = v_20599 & 1'h1;
  assign v_20599 = v_20600 | 1'h0;
  assign v_20600 = ~v_20507;
  assign v_20601 = mux_20601(v_20602);
  assign v_20602 = ~v_20597;
  assign v_20603 = ~v_20514;
  assign v_20604 = v_20605 | v_20606;
  assign v_20605 = mux_20605(v_20516);
  assign v_20606 = mux_20606(v_20591);
  assign v_20608 = v_20609 | v_20684;
  assign v_20609 = act_20610 & 1'h1;
  assign act_20610 = v_20611 | v_20641;
  assign v_20611 = v_20612 & v_20642;
  assign v_20612 = v_20613 & v_20651;
  assign v_20613 = ~v_20614;
  assign v_20615 = v_20616 | v_20635;
  assign v_20616 = act_20617 & 1'h1;
  assign act_20617 = v_20618 | v_20624;
  assign v_20618 = v_20619 & v_20625;
  assign v_20619 = v_20620 & vout_canPeek_20630;
  assign v_20620 = ~vout_canPeek_20621;
  pebbles_core
    pebbles_core_20621
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20622),
       .in0_consume_en(vin0_consume_en_20621),
       .out_canPeek(vout_canPeek_20621),
       .out_peek(vout_peek_20621));
  assign v_20622 = v_20623 | v_20628;
  assign v_20623 = mux_20623(v_20624);
  assign v_20624 = vout_canPeek_20621 & v_20625;
  assign v_20625 = v_20626 & 1'h1;
  assign v_20626 = v_20627 | 1'h0;
  assign v_20627 = ~v_20614;
  assign v_20628 = mux_20628(v_20629);
  assign v_20629 = ~v_20624;
  pebbles_core
    pebbles_core_20630
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20631),
       .in0_consume_en(vin0_consume_en_20630),
       .out_canPeek(vout_canPeek_20630),
       .out_peek(vout_peek_20630));
  assign v_20631 = v_20632 | v_20633;
  assign v_20632 = mux_20632(v_20618);
  assign v_20633 = mux_20633(v_20634);
  assign v_20634 = ~v_20618;
  assign v_20635 = v_20636 & 1'h1;
  assign v_20636 = v_20637 & v_20638;
  assign v_20637 = ~act_20617;
  assign v_20638 = v_20639 | v_20647;
  assign v_20639 = v_20640 | v_20645;
  assign v_20640 = mux_20640(v_20641);
  assign v_20641 = v_20614 & v_20642;
  assign v_20642 = v_20643 & 1'h1;
  assign v_20643 = v_20644 | 1'h0;
  assign v_20644 = ~v_20607;
  assign v_20645 = mux_20645(v_20646);
  assign v_20646 = ~v_20641;
  assign v_20647 = ~v_20614;
  assign v_20648 = v_20649 | v_20650;
  assign v_20649 = mux_20649(v_20616);
  assign v_20650 = mux_20650(v_20635);
  assign v_20652 = v_20653 | v_20672;
  assign v_20653 = act_20654 & 1'h1;
  assign act_20654 = v_20655 | v_20661;
  assign v_20655 = v_20656 & v_20662;
  assign v_20656 = v_20657 & vout_canPeek_20667;
  assign v_20657 = ~vout_canPeek_20658;
  pebbles_core
    pebbles_core_20658
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20659),
       .in0_consume_en(vin0_consume_en_20658),
       .out_canPeek(vout_canPeek_20658),
       .out_peek(vout_peek_20658));
  assign v_20659 = v_20660 | v_20665;
  assign v_20660 = mux_20660(v_20661);
  assign v_20661 = vout_canPeek_20658 & v_20662;
  assign v_20662 = v_20663 & 1'h1;
  assign v_20663 = v_20664 | 1'h0;
  assign v_20664 = ~v_20651;
  assign v_20665 = mux_20665(v_20666);
  assign v_20666 = ~v_20661;
  pebbles_core
    pebbles_core_20667
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20668),
       .in0_consume_en(vin0_consume_en_20667),
       .out_canPeek(vout_canPeek_20667),
       .out_peek(vout_peek_20667));
  assign v_20668 = v_20669 | v_20670;
  assign v_20669 = mux_20669(v_20655);
  assign v_20670 = mux_20670(v_20671);
  assign v_20671 = ~v_20655;
  assign v_20672 = v_20673 & 1'h1;
  assign v_20673 = v_20674 & v_20675;
  assign v_20674 = ~act_20654;
  assign v_20675 = v_20676 | v_20680;
  assign v_20676 = v_20677 | v_20678;
  assign v_20677 = mux_20677(v_20611);
  assign v_20678 = mux_20678(v_20679);
  assign v_20679 = ~v_20611;
  assign v_20680 = ~v_20651;
  assign v_20681 = v_20682 | v_20683;
  assign v_20682 = mux_20682(v_20653);
  assign v_20683 = mux_20683(v_20672);
  assign v_20684 = v_20685 & 1'h1;
  assign v_20685 = v_20686 & v_20687;
  assign v_20686 = ~act_20610;
  assign v_20687 = v_20688 | v_20692;
  assign v_20688 = v_20689 | v_20690;
  assign v_20689 = mux_20689(v_20511);
  assign v_20690 = mux_20690(v_20691);
  assign v_20691 = ~v_20511;
  assign v_20692 = ~v_20607;
  assign v_20693 = v_20694 | v_20695;
  assign v_20694 = mux_20694(v_20609);
  assign v_20695 = mux_20695(v_20684);
  assign v_20696 = v_20697 & 1'h1;
  assign v_20697 = v_20698 & v_20699;
  assign v_20698 = ~act_20510;
  assign v_20699 = v_20700 | v_20708;
  assign v_20700 = v_20701 | v_20706;
  assign v_20701 = mux_20701(v_20702);
  assign v_20702 = v_20507 & v_20703;
  assign v_20703 = v_20704 & 1'h1;
  assign v_20704 = v_20705 | 1'h0;
  assign v_20705 = ~v_20500;
  assign v_20706 = mux_20706(v_20707);
  assign v_20707 = ~v_20702;
  assign v_20708 = ~v_20507;
  assign v_20709 = v_20710 | v_20711;
  assign v_20710 = mux_20710(v_20509);
  assign v_20711 = mux_20711(v_20696);
  assign v_20713 = v_20714 | v_20901;
  assign v_20714 = act_20715 & 1'h1;
  assign act_20715 = v_20716 | v_20802;
  assign v_20716 = v_20717 & v_20803;
  assign v_20717 = v_20718 & v_20812;
  assign v_20718 = ~v_20719;
  assign v_20720 = v_20721 | v_20796;
  assign v_20721 = act_20722 & 1'h1;
  assign act_20722 = v_20723 | v_20753;
  assign v_20723 = v_20724 & v_20754;
  assign v_20724 = v_20725 & v_20763;
  assign v_20725 = ~v_20726;
  assign v_20727 = v_20728 | v_20747;
  assign v_20728 = act_20729 & 1'h1;
  assign act_20729 = v_20730 | v_20736;
  assign v_20730 = v_20731 & v_20737;
  assign v_20731 = v_20732 & vout_canPeek_20742;
  assign v_20732 = ~vout_canPeek_20733;
  pebbles_core
    pebbles_core_20733
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20734),
       .in0_consume_en(vin0_consume_en_20733),
       .out_canPeek(vout_canPeek_20733),
       .out_peek(vout_peek_20733));
  assign v_20734 = v_20735 | v_20740;
  assign v_20735 = mux_20735(v_20736);
  assign v_20736 = vout_canPeek_20733 & v_20737;
  assign v_20737 = v_20738 & 1'h1;
  assign v_20738 = v_20739 | 1'h0;
  assign v_20739 = ~v_20726;
  assign v_20740 = mux_20740(v_20741);
  assign v_20741 = ~v_20736;
  pebbles_core
    pebbles_core_20742
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20743),
       .in0_consume_en(vin0_consume_en_20742),
       .out_canPeek(vout_canPeek_20742),
       .out_peek(vout_peek_20742));
  assign v_20743 = v_20744 | v_20745;
  assign v_20744 = mux_20744(v_20730);
  assign v_20745 = mux_20745(v_20746);
  assign v_20746 = ~v_20730;
  assign v_20747 = v_20748 & 1'h1;
  assign v_20748 = v_20749 & v_20750;
  assign v_20749 = ~act_20729;
  assign v_20750 = v_20751 | v_20759;
  assign v_20751 = v_20752 | v_20757;
  assign v_20752 = mux_20752(v_20753);
  assign v_20753 = v_20726 & v_20754;
  assign v_20754 = v_20755 & 1'h1;
  assign v_20755 = v_20756 | 1'h0;
  assign v_20756 = ~v_20719;
  assign v_20757 = mux_20757(v_20758);
  assign v_20758 = ~v_20753;
  assign v_20759 = ~v_20726;
  assign v_20760 = v_20761 | v_20762;
  assign v_20761 = mux_20761(v_20728);
  assign v_20762 = mux_20762(v_20747);
  assign v_20764 = v_20765 | v_20784;
  assign v_20765 = act_20766 & 1'h1;
  assign act_20766 = v_20767 | v_20773;
  assign v_20767 = v_20768 & v_20774;
  assign v_20768 = v_20769 & vout_canPeek_20779;
  assign v_20769 = ~vout_canPeek_20770;
  pebbles_core
    pebbles_core_20770
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20771),
       .in0_consume_en(vin0_consume_en_20770),
       .out_canPeek(vout_canPeek_20770),
       .out_peek(vout_peek_20770));
  assign v_20771 = v_20772 | v_20777;
  assign v_20772 = mux_20772(v_20773);
  assign v_20773 = vout_canPeek_20770 & v_20774;
  assign v_20774 = v_20775 & 1'h1;
  assign v_20775 = v_20776 | 1'h0;
  assign v_20776 = ~v_20763;
  assign v_20777 = mux_20777(v_20778);
  assign v_20778 = ~v_20773;
  pebbles_core
    pebbles_core_20779
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20780),
       .in0_consume_en(vin0_consume_en_20779),
       .out_canPeek(vout_canPeek_20779),
       .out_peek(vout_peek_20779));
  assign v_20780 = v_20781 | v_20782;
  assign v_20781 = mux_20781(v_20767);
  assign v_20782 = mux_20782(v_20783);
  assign v_20783 = ~v_20767;
  assign v_20784 = v_20785 & 1'h1;
  assign v_20785 = v_20786 & v_20787;
  assign v_20786 = ~act_20766;
  assign v_20787 = v_20788 | v_20792;
  assign v_20788 = v_20789 | v_20790;
  assign v_20789 = mux_20789(v_20723);
  assign v_20790 = mux_20790(v_20791);
  assign v_20791 = ~v_20723;
  assign v_20792 = ~v_20763;
  assign v_20793 = v_20794 | v_20795;
  assign v_20794 = mux_20794(v_20765);
  assign v_20795 = mux_20795(v_20784);
  assign v_20796 = v_20797 & 1'h1;
  assign v_20797 = v_20798 & v_20799;
  assign v_20798 = ~act_20722;
  assign v_20799 = v_20800 | v_20808;
  assign v_20800 = v_20801 | v_20806;
  assign v_20801 = mux_20801(v_20802);
  assign v_20802 = v_20719 & v_20803;
  assign v_20803 = v_20804 & 1'h1;
  assign v_20804 = v_20805 | 1'h0;
  assign v_20805 = ~v_20712;
  assign v_20806 = mux_20806(v_20807);
  assign v_20807 = ~v_20802;
  assign v_20808 = ~v_20719;
  assign v_20809 = v_20810 | v_20811;
  assign v_20810 = mux_20810(v_20721);
  assign v_20811 = mux_20811(v_20796);
  assign v_20813 = v_20814 | v_20889;
  assign v_20814 = act_20815 & 1'h1;
  assign act_20815 = v_20816 | v_20846;
  assign v_20816 = v_20817 & v_20847;
  assign v_20817 = v_20818 & v_20856;
  assign v_20818 = ~v_20819;
  assign v_20820 = v_20821 | v_20840;
  assign v_20821 = act_20822 & 1'h1;
  assign act_20822 = v_20823 | v_20829;
  assign v_20823 = v_20824 & v_20830;
  assign v_20824 = v_20825 & vout_canPeek_20835;
  assign v_20825 = ~vout_canPeek_20826;
  pebbles_core
    pebbles_core_20826
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20827),
       .in0_consume_en(vin0_consume_en_20826),
       .out_canPeek(vout_canPeek_20826),
       .out_peek(vout_peek_20826));
  assign v_20827 = v_20828 | v_20833;
  assign v_20828 = mux_20828(v_20829);
  assign v_20829 = vout_canPeek_20826 & v_20830;
  assign v_20830 = v_20831 & 1'h1;
  assign v_20831 = v_20832 | 1'h0;
  assign v_20832 = ~v_20819;
  assign v_20833 = mux_20833(v_20834);
  assign v_20834 = ~v_20829;
  pebbles_core
    pebbles_core_20835
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20836),
       .in0_consume_en(vin0_consume_en_20835),
       .out_canPeek(vout_canPeek_20835),
       .out_peek(vout_peek_20835));
  assign v_20836 = v_20837 | v_20838;
  assign v_20837 = mux_20837(v_20823);
  assign v_20838 = mux_20838(v_20839);
  assign v_20839 = ~v_20823;
  assign v_20840 = v_20841 & 1'h1;
  assign v_20841 = v_20842 & v_20843;
  assign v_20842 = ~act_20822;
  assign v_20843 = v_20844 | v_20852;
  assign v_20844 = v_20845 | v_20850;
  assign v_20845 = mux_20845(v_20846);
  assign v_20846 = v_20819 & v_20847;
  assign v_20847 = v_20848 & 1'h1;
  assign v_20848 = v_20849 | 1'h0;
  assign v_20849 = ~v_20812;
  assign v_20850 = mux_20850(v_20851);
  assign v_20851 = ~v_20846;
  assign v_20852 = ~v_20819;
  assign v_20853 = v_20854 | v_20855;
  assign v_20854 = mux_20854(v_20821);
  assign v_20855 = mux_20855(v_20840);
  assign v_20857 = v_20858 | v_20877;
  assign v_20858 = act_20859 & 1'h1;
  assign act_20859 = v_20860 | v_20866;
  assign v_20860 = v_20861 & v_20867;
  assign v_20861 = v_20862 & vout_canPeek_20872;
  assign v_20862 = ~vout_canPeek_20863;
  pebbles_core
    pebbles_core_20863
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20864),
       .in0_consume_en(vin0_consume_en_20863),
       .out_canPeek(vout_canPeek_20863),
       .out_peek(vout_peek_20863));
  assign v_20864 = v_20865 | v_20870;
  assign v_20865 = mux_20865(v_20866);
  assign v_20866 = vout_canPeek_20863 & v_20867;
  assign v_20867 = v_20868 & 1'h1;
  assign v_20868 = v_20869 | 1'h0;
  assign v_20869 = ~v_20856;
  assign v_20870 = mux_20870(v_20871);
  assign v_20871 = ~v_20866;
  pebbles_core
    pebbles_core_20872
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20873),
       .in0_consume_en(vin0_consume_en_20872),
       .out_canPeek(vout_canPeek_20872),
       .out_peek(vout_peek_20872));
  assign v_20873 = v_20874 | v_20875;
  assign v_20874 = mux_20874(v_20860);
  assign v_20875 = mux_20875(v_20876);
  assign v_20876 = ~v_20860;
  assign v_20877 = v_20878 & 1'h1;
  assign v_20878 = v_20879 & v_20880;
  assign v_20879 = ~act_20859;
  assign v_20880 = v_20881 | v_20885;
  assign v_20881 = v_20882 | v_20883;
  assign v_20882 = mux_20882(v_20816);
  assign v_20883 = mux_20883(v_20884);
  assign v_20884 = ~v_20816;
  assign v_20885 = ~v_20856;
  assign v_20886 = v_20887 | v_20888;
  assign v_20887 = mux_20887(v_20858);
  assign v_20888 = mux_20888(v_20877);
  assign v_20889 = v_20890 & 1'h1;
  assign v_20890 = v_20891 & v_20892;
  assign v_20891 = ~act_20815;
  assign v_20892 = v_20893 | v_20897;
  assign v_20893 = v_20894 | v_20895;
  assign v_20894 = mux_20894(v_20716);
  assign v_20895 = mux_20895(v_20896);
  assign v_20896 = ~v_20716;
  assign v_20897 = ~v_20812;
  assign v_20898 = v_20899 | v_20900;
  assign v_20899 = mux_20899(v_20814);
  assign v_20900 = mux_20900(v_20889);
  assign v_20901 = v_20902 & 1'h1;
  assign v_20902 = v_20903 & v_20904;
  assign v_20903 = ~act_20715;
  assign v_20904 = v_20905 | v_20909;
  assign v_20905 = v_20906 | v_20907;
  assign v_20906 = mux_20906(v_20504);
  assign v_20907 = mux_20907(v_20908);
  assign v_20908 = ~v_20504;
  assign v_20909 = ~v_20712;
  assign v_20910 = v_20911 | v_20912;
  assign v_20911 = mux_20911(v_20714);
  assign v_20912 = mux_20912(v_20901);
  assign v_20913 = v_20914 & 1'h1;
  assign v_20914 = v_20915 & v_20916;
  assign v_20915 = ~act_20503;
  assign v_20916 = v_20917 | v_20925;
  assign v_20917 = v_20918 | v_20923;
  assign v_20918 = mux_20918(v_20919);
  assign v_20919 = v_20500 & v_20920;
  assign v_20920 = v_20921 & 1'h1;
  assign v_20921 = v_20922 | 1'h0;
  assign v_20922 = ~v_20493;
  assign v_20923 = mux_20923(v_20924);
  assign v_20924 = ~v_20919;
  assign v_20925 = ~v_20500;
  assign v_20926 = v_20927 | v_20928;
  assign v_20927 = mux_20927(v_20502);
  assign v_20928 = mux_20928(v_20913);
  assign v_20930 = v_20931 | v_21342;
  assign v_20931 = act_20932 & 1'h1;
  assign act_20932 = v_20933 | v_21131;
  assign v_20933 = v_20934 & v_21132;
  assign v_20934 = v_20935 & v_21141;
  assign v_20935 = ~v_20936;
  assign v_20937 = v_20938 | v_21125;
  assign v_20938 = act_20939 & 1'h1;
  assign act_20939 = v_20940 | v_21026;
  assign v_20940 = v_20941 & v_21027;
  assign v_20941 = v_20942 & v_21036;
  assign v_20942 = ~v_20943;
  assign v_20944 = v_20945 | v_21020;
  assign v_20945 = act_20946 & 1'h1;
  assign act_20946 = v_20947 | v_20977;
  assign v_20947 = v_20948 & v_20978;
  assign v_20948 = v_20949 & v_20987;
  assign v_20949 = ~v_20950;
  assign v_20951 = v_20952 | v_20971;
  assign v_20952 = act_20953 & 1'h1;
  assign act_20953 = v_20954 | v_20960;
  assign v_20954 = v_20955 & v_20961;
  assign v_20955 = v_20956 & vout_canPeek_20966;
  assign v_20956 = ~vout_canPeek_20957;
  pebbles_core
    pebbles_core_20957
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20958),
       .in0_consume_en(vin0_consume_en_20957),
       .out_canPeek(vout_canPeek_20957),
       .out_peek(vout_peek_20957));
  assign v_20958 = v_20959 | v_20964;
  assign v_20959 = mux_20959(v_20960);
  assign v_20960 = vout_canPeek_20957 & v_20961;
  assign v_20961 = v_20962 & 1'h1;
  assign v_20962 = v_20963 | 1'h0;
  assign v_20963 = ~v_20950;
  assign v_20964 = mux_20964(v_20965);
  assign v_20965 = ~v_20960;
  pebbles_core
    pebbles_core_20966
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20967),
       .in0_consume_en(vin0_consume_en_20966),
       .out_canPeek(vout_canPeek_20966),
       .out_peek(vout_peek_20966));
  assign v_20967 = v_20968 | v_20969;
  assign v_20968 = mux_20968(v_20954);
  assign v_20969 = mux_20969(v_20970);
  assign v_20970 = ~v_20954;
  assign v_20971 = v_20972 & 1'h1;
  assign v_20972 = v_20973 & v_20974;
  assign v_20973 = ~act_20953;
  assign v_20974 = v_20975 | v_20983;
  assign v_20975 = v_20976 | v_20981;
  assign v_20976 = mux_20976(v_20977);
  assign v_20977 = v_20950 & v_20978;
  assign v_20978 = v_20979 & 1'h1;
  assign v_20979 = v_20980 | 1'h0;
  assign v_20980 = ~v_20943;
  assign v_20981 = mux_20981(v_20982);
  assign v_20982 = ~v_20977;
  assign v_20983 = ~v_20950;
  assign v_20984 = v_20985 | v_20986;
  assign v_20985 = mux_20985(v_20952);
  assign v_20986 = mux_20986(v_20971);
  assign v_20988 = v_20989 | v_21008;
  assign v_20989 = act_20990 & 1'h1;
  assign act_20990 = v_20991 | v_20997;
  assign v_20991 = v_20992 & v_20998;
  assign v_20992 = v_20993 & vout_canPeek_21003;
  assign v_20993 = ~vout_canPeek_20994;
  pebbles_core
    pebbles_core_20994
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20995),
       .in0_consume_en(vin0_consume_en_20994),
       .out_canPeek(vout_canPeek_20994),
       .out_peek(vout_peek_20994));
  assign v_20995 = v_20996 | v_21001;
  assign v_20996 = mux_20996(v_20997);
  assign v_20997 = vout_canPeek_20994 & v_20998;
  assign v_20998 = v_20999 & 1'h1;
  assign v_20999 = v_21000 | 1'h0;
  assign v_21000 = ~v_20987;
  assign v_21001 = mux_21001(v_21002);
  assign v_21002 = ~v_20997;
  pebbles_core
    pebbles_core_21003
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21004),
       .in0_consume_en(vin0_consume_en_21003),
       .out_canPeek(vout_canPeek_21003),
       .out_peek(vout_peek_21003));
  assign v_21004 = v_21005 | v_21006;
  assign v_21005 = mux_21005(v_20991);
  assign v_21006 = mux_21006(v_21007);
  assign v_21007 = ~v_20991;
  assign v_21008 = v_21009 & 1'h1;
  assign v_21009 = v_21010 & v_21011;
  assign v_21010 = ~act_20990;
  assign v_21011 = v_21012 | v_21016;
  assign v_21012 = v_21013 | v_21014;
  assign v_21013 = mux_21013(v_20947);
  assign v_21014 = mux_21014(v_21015);
  assign v_21015 = ~v_20947;
  assign v_21016 = ~v_20987;
  assign v_21017 = v_21018 | v_21019;
  assign v_21018 = mux_21018(v_20989);
  assign v_21019 = mux_21019(v_21008);
  assign v_21020 = v_21021 & 1'h1;
  assign v_21021 = v_21022 & v_21023;
  assign v_21022 = ~act_20946;
  assign v_21023 = v_21024 | v_21032;
  assign v_21024 = v_21025 | v_21030;
  assign v_21025 = mux_21025(v_21026);
  assign v_21026 = v_20943 & v_21027;
  assign v_21027 = v_21028 & 1'h1;
  assign v_21028 = v_21029 | 1'h0;
  assign v_21029 = ~v_20936;
  assign v_21030 = mux_21030(v_21031);
  assign v_21031 = ~v_21026;
  assign v_21032 = ~v_20943;
  assign v_21033 = v_21034 | v_21035;
  assign v_21034 = mux_21034(v_20945);
  assign v_21035 = mux_21035(v_21020);
  assign v_21037 = v_21038 | v_21113;
  assign v_21038 = act_21039 & 1'h1;
  assign act_21039 = v_21040 | v_21070;
  assign v_21040 = v_21041 & v_21071;
  assign v_21041 = v_21042 & v_21080;
  assign v_21042 = ~v_21043;
  assign v_21044 = v_21045 | v_21064;
  assign v_21045 = act_21046 & 1'h1;
  assign act_21046 = v_21047 | v_21053;
  assign v_21047 = v_21048 & v_21054;
  assign v_21048 = v_21049 & vout_canPeek_21059;
  assign v_21049 = ~vout_canPeek_21050;
  pebbles_core
    pebbles_core_21050
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21051),
       .in0_consume_en(vin0_consume_en_21050),
       .out_canPeek(vout_canPeek_21050),
       .out_peek(vout_peek_21050));
  assign v_21051 = v_21052 | v_21057;
  assign v_21052 = mux_21052(v_21053);
  assign v_21053 = vout_canPeek_21050 & v_21054;
  assign v_21054 = v_21055 & 1'h1;
  assign v_21055 = v_21056 | 1'h0;
  assign v_21056 = ~v_21043;
  assign v_21057 = mux_21057(v_21058);
  assign v_21058 = ~v_21053;
  pebbles_core
    pebbles_core_21059
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21060),
       .in0_consume_en(vin0_consume_en_21059),
       .out_canPeek(vout_canPeek_21059),
       .out_peek(vout_peek_21059));
  assign v_21060 = v_21061 | v_21062;
  assign v_21061 = mux_21061(v_21047);
  assign v_21062 = mux_21062(v_21063);
  assign v_21063 = ~v_21047;
  assign v_21064 = v_21065 & 1'h1;
  assign v_21065 = v_21066 & v_21067;
  assign v_21066 = ~act_21046;
  assign v_21067 = v_21068 | v_21076;
  assign v_21068 = v_21069 | v_21074;
  assign v_21069 = mux_21069(v_21070);
  assign v_21070 = v_21043 & v_21071;
  assign v_21071 = v_21072 & 1'h1;
  assign v_21072 = v_21073 | 1'h0;
  assign v_21073 = ~v_21036;
  assign v_21074 = mux_21074(v_21075);
  assign v_21075 = ~v_21070;
  assign v_21076 = ~v_21043;
  assign v_21077 = v_21078 | v_21079;
  assign v_21078 = mux_21078(v_21045);
  assign v_21079 = mux_21079(v_21064);
  assign v_21081 = v_21082 | v_21101;
  assign v_21082 = act_21083 & 1'h1;
  assign act_21083 = v_21084 | v_21090;
  assign v_21084 = v_21085 & v_21091;
  assign v_21085 = v_21086 & vout_canPeek_21096;
  assign v_21086 = ~vout_canPeek_21087;
  pebbles_core
    pebbles_core_21087
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21088),
       .in0_consume_en(vin0_consume_en_21087),
       .out_canPeek(vout_canPeek_21087),
       .out_peek(vout_peek_21087));
  assign v_21088 = v_21089 | v_21094;
  assign v_21089 = mux_21089(v_21090);
  assign v_21090 = vout_canPeek_21087 & v_21091;
  assign v_21091 = v_21092 & 1'h1;
  assign v_21092 = v_21093 | 1'h0;
  assign v_21093 = ~v_21080;
  assign v_21094 = mux_21094(v_21095);
  assign v_21095 = ~v_21090;
  pebbles_core
    pebbles_core_21096
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21097),
       .in0_consume_en(vin0_consume_en_21096),
       .out_canPeek(vout_canPeek_21096),
       .out_peek(vout_peek_21096));
  assign v_21097 = v_21098 | v_21099;
  assign v_21098 = mux_21098(v_21084);
  assign v_21099 = mux_21099(v_21100);
  assign v_21100 = ~v_21084;
  assign v_21101 = v_21102 & 1'h1;
  assign v_21102 = v_21103 & v_21104;
  assign v_21103 = ~act_21083;
  assign v_21104 = v_21105 | v_21109;
  assign v_21105 = v_21106 | v_21107;
  assign v_21106 = mux_21106(v_21040);
  assign v_21107 = mux_21107(v_21108);
  assign v_21108 = ~v_21040;
  assign v_21109 = ~v_21080;
  assign v_21110 = v_21111 | v_21112;
  assign v_21111 = mux_21111(v_21082);
  assign v_21112 = mux_21112(v_21101);
  assign v_21113 = v_21114 & 1'h1;
  assign v_21114 = v_21115 & v_21116;
  assign v_21115 = ~act_21039;
  assign v_21116 = v_21117 | v_21121;
  assign v_21117 = v_21118 | v_21119;
  assign v_21118 = mux_21118(v_20940);
  assign v_21119 = mux_21119(v_21120);
  assign v_21120 = ~v_20940;
  assign v_21121 = ~v_21036;
  assign v_21122 = v_21123 | v_21124;
  assign v_21123 = mux_21123(v_21038);
  assign v_21124 = mux_21124(v_21113);
  assign v_21125 = v_21126 & 1'h1;
  assign v_21126 = v_21127 & v_21128;
  assign v_21127 = ~act_20939;
  assign v_21128 = v_21129 | v_21137;
  assign v_21129 = v_21130 | v_21135;
  assign v_21130 = mux_21130(v_21131);
  assign v_21131 = v_20936 & v_21132;
  assign v_21132 = v_21133 & 1'h1;
  assign v_21133 = v_21134 | 1'h0;
  assign v_21134 = ~v_20929;
  assign v_21135 = mux_21135(v_21136);
  assign v_21136 = ~v_21131;
  assign v_21137 = ~v_20936;
  assign v_21138 = v_21139 | v_21140;
  assign v_21139 = mux_21139(v_20938);
  assign v_21140 = mux_21140(v_21125);
  assign v_21142 = v_21143 | v_21330;
  assign v_21143 = act_21144 & 1'h1;
  assign act_21144 = v_21145 | v_21231;
  assign v_21145 = v_21146 & v_21232;
  assign v_21146 = v_21147 & v_21241;
  assign v_21147 = ~v_21148;
  assign v_21149 = v_21150 | v_21225;
  assign v_21150 = act_21151 & 1'h1;
  assign act_21151 = v_21152 | v_21182;
  assign v_21152 = v_21153 & v_21183;
  assign v_21153 = v_21154 & v_21192;
  assign v_21154 = ~v_21155;
  assign v_21156 = v_21157 | v_21176;
  assign v_21157 = act_21158 & 1'h1;
  assign act_21158 = v_21159 | v_21165;
  assign v_21159 = v_21160 & v_21166;
  assign v_21160 = v_21161 & vout_canPeek_21171;
  assign v_21161 = ~vout_canPeek_21162;
  pebbles_core
    pebbles_core_21162
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21163),
       .in0_consume_en(vin0_consume_en_21162),
       .out_canPeek(vout_canPeek_21162),
       .out_peek(vout_peek_21162));
  assign v_21163 = v_21164 | v_21169;
  assign v_21164 = mux_21164(v_21165);
  assign v_21165 = vout_canPeek_21162 & v_21166;
  assign v_21166 = v_21167 & 1'h1;
  assign v_21167 = v_21168 | 1'h0;
  assign v_21168 = ~v_21155;
  assign v_21169 = mux_21169(v_21170);
  assign v_21170 = ~v_21165;
  pebbles_core
    pebbles_core_21171
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21172),
       .in0_consume_en(vin0_consume_en_21171),
       .out_canPeek(vout_canPeek_21171),
       .out_peek(vout_peek_21171));
  assign v_21172 = v_21173 | v_21174;
  assign v_21173 = mux_21173(v_21159);
  assign v_21174 = mux_21174(v_21175);
  assign v_21175 = ~v_21159;
  assign v_21176 = v_21177 & 1'h1;
  assign v_21177 = v_21178 & v_21179;
  assign v_21178 = ~act_21158;
  assign v_21179 = v_21180 | v_21188;
  assign v_21180 = v_21181 | v_21186;
  assign v_21181 = mux_21181(v_21182);
  assign v_21182 = v_21155 & v_21183;
  assign v_21183 = v_21184 & 1'h1;
  assign v_21184 = v_21185 | 1'h0;
  assign v_21185 = ~v_21148;
  assign v_21186 = mux_21186(v_21187);
  assign v_21187 = ~v_21182;
  assign v_21188 = ~v_21155;
  assign v_21189 = v_21190 | v_21191;
  assign v_21190 = mux_21190(v_21157);
  assign v_21191 = mux_21191(v_21176);
  assign v_21193 = v_21194 | v_21213;
  assign v_21194 = act_21195 & 1'h1;
  assign act_21195 = v_21196 | v_21202;
  assign v_21196 = v_21197 & v_21203;
  assign v_21197 = v_21198 & vout_canPeek_21208;
  assign v_21198 = ~vout_canPeek_21199;
  pebbles_core
    pebbles_core_21199
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21200),
       .in0_consume_en(vin0_consume_en_21199),
       .out_canPeek(vout_canPeek_21199),
       .out_peek(vout_peek_21199));
  assign v_21200 = v_21201 | v_21206;
  assign v_21201 = mux_21201(v_21202);
  assign v_21202 = vout_canPeek_21199 & v_21203;
  assign v_21203 = v_21204 & 1'h1;
  assign v_21204 = v_21205 | 1'h0;
  assign v_21205 = ~v_21192;
  assign v_21206 = mux_21206(v_21207);
  assign v_21207 = ~v_21202;
  pebbles_core
    pebbles_core_21208
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21209),
       .in0_consume_en(vin0_consume_en_21208),
       .out_canPeek(vout_canPeek_21208),
       .out_peek(vout_peek_21208));
  assign v_21209 = v_21210 | v_21211;
  assign v_21210 = mux_21210(v_21196);
  assign v_21211 = mux_21211(v_21212);
  assign v_21212 = ~v_21196;
  assign v_21213 = v_21214 & 1'h1;
  assign v_21214 = v_21215 & v_21216;
  assign v_21215 = ~act_21195;
  assign v_21216 = v_21217 | v_21221;
  assign v_21217 = v_21218 | v_21219;
  assign v_21218 = mux_21218(v_21152);
  assign v_21219 = mux_21219(v_21220);
  assign v_21220 = ~v_21152;
  assign v_21221 = ~v_21192;
  assign v_21222 = v_21223 | v_21224;
  assign v_21223 = mux_21223(v_21194);
  assign v_21224 = mux_21224(v_21213);
  assign v_21225 = v_21226 & 1'h1;
  assign v_21226 = v_21227 & v_21228;
  assign v_21227 = ~act_21151;
  assign v_21228 = v_21229 | v_21237;
  assign v_21229 = v_21230 | v_21235;
  assign v_21230 = mux_21230(v_21231);
  assign v_21231 = v_21148 & v_21232;
  assign v_21232 = v_21233 & 1'h1;
  assign v_21233 = v_21234 | 1'h0;
  assign v_21234 = ~v_21141;
  assign v_21235 = mux_21235(v_21236);
  assign v_21236 = ~v_21231;
  assign v_21237 = ~v_21148;
  assign v_21238 = v_21239 | v_21240;
  assign v_21239 = mux_21239(v_21150);
  assign v_21240 = mux_21240(v_21225);
  assign v_21242 = v_21243 | v_21318;
  assign v_21243 = act_21244 & 1'h1;
  assign act_21244 = v_21245 | v_21275;
  assign v_21245 = v_21246 & v_21276;
  assign v_21246 = v_21247 & v_21285;
  assign v_21247 = ~v_21248;
  assign v_21249 = v_21250 | v_21269;
  assign v_21250 = act_21251 & 1'h1;
  assign act_21251 = v_21252 | v_21258;
  assign v_21252 = v_21253 & v_21259;
  assign v_21253 = v_21254 & vout_canPeek_21264;
  assign v_21254 = ~vout_canPeek_21255;
  pebbles_core
    pebbles_core_21255
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21256),
       .in0_consume_en(vin0_consume_en_21255),
       .out_canPeek(vout_canPeek_21255),
       .out_peek(vout_peek_21255));
  assign v_21256 = v_21257 | v_21262;
  assign v_21257 = mux_21257(v_21258);
  assign v_21258 = vout_canPeek_21255 & v_21259;
  assign v_21259 = v_21260 & 1'h1;
  assign v_21260 = v_21261 | 1'h0;
  assign v_21261 = ~v_21248;
  assign v_21262 = mux_21262(v_21263);
  assign v_21263 = ~v_21258;
  pebbles_core
    pebbles_core_21264
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21265),
       .in0_consume_en(vin0_consume_en_21264),
       .out_canPeek(vout_canPeek_21264),
       .out_peek(vout_peek_21264));
  assign v_21265 = v_21266 | v_21267;
  assign v_21266 = mux_21266(v_21252);
  assign v_21267 = mux_21267(v_21268);
  assign v_21268 = ~v_21252;
  assign v_21269 = v_21270 & 1'h1;
  assign v_21270 = v_21271 & v_21272;
  assign v_21271 = ~act_21251;
  assign v_21272 = v_21273 | v_21281;
  assign v_21273 = v_21274 | v_21279;
  assign v_21274 = mux_21274(v_21275);
  assign v_21275 = v_21248 & v_21276;
  assign v_21276 = v_21277 & 1'h1;
  assign v_21277 = v_21278 | 1'h0;
  assign v_21278 = ~v_21241;
  assign v_21279 = mux_21279(v_21280);
  assign v_21280 = ~v_21275;
  assign v_21281 = ~v_21248;
  assign v_21282 = v_21283 | v_21284;
  assign v_21283 = mux_21283(v_21250);
  assign v_21284 = mux_21284(v_21269);
  assign v_21286 = v_21287 | v_21306;
  assign v_21287 = act_21288 & 1'h1;
  assign act_21288 = v_21289 | v_21295;
  assign v_21289 = v_21290 & v_21296;
  assign v_21290 = v_21291 & vout_canPeek_21301;
  assign v_21291 = ~vout_canPeek_21292;
  pebbles_core
    pebbles_core_21292
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21293),
       .in0_consume_en(vin0_consume_en_21292),
       .out_canPeek(vout_canPeek_21292),
       .out_peek(vout_peek_21292));
  assign v_21293 = v_21294 | v_21299;
  assign v_21294 = mux_21294(v_21295);
  assign v_21295 = vout_canPeek_21292 & v_21296;
  assign v_21296 = v_21297 & 1'h1;
  assign v_21297 = v_21298 | 1'h0;
  assign v_21298 = ~v_21285;
  assign v_21299 = mux_21299(v_21300);
  assign v_21300 = ~v_21295;
  pebbles_core
    pebbles_core_21301
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21302),
       .in0_consume_en(vin0_consume_en_21301),
       .out_canPeek(vout_canPeek_21301),
       .out_peek(vout_peek_21301));
  assign v_21302 = v_21303 | v_21304;
  assign v_21303 = mux_21303(v_21289);
  assign v_21304 = mux_21304(v_21305);
  assign v_21305 = ~v_21289;
  assign v_21306 = v_21307 & 1'h1;
  assign v_21307 = v_21308 & v_21309;
  assign v_21308 = ~act_21288;
  assign v_21309 = v_21310 | v_21314;
  assign v_21310 = v_21311 | v_21312;
  assign v_21311 = mux_21311(v_21245);
  assign v_21312 = mux_21312(v_21313);
  assign v_21313 = ~v_21245;
  assign v_21314 = ~v_21285;
  assign v_21315 = v_21316 | v_21317;
  assign v_21316 = mux_21316(v_21287);
  assign v_21317 = mux_21317(v_21306);
  assign v_21318 = v_21319 & 1'h1;
  assign v_21319 = v_21320 & v_21321;
  assign v_21320 = ~act_21244;
  assign v_21321 = v_21322 | v_21326;
  assign v_21322 = v_21323 | v_21324;
  assign v_21323 = mux_21323(v_21145);
  assign v_21324 = mux_21324(v_21325);
  assign v_21325 = ~v_21145;
  assign v_21326 = ~v_21241;
  assign v_21327 = v_21328 | v_21329;
  assign v_21328 = mux_21328(v_21243);
  assign v_21329 = mux_21329(v_21318);
  assign v_21330 = v_21331 & 1'h1;
  assign v_21331 = v_21332 & v_21333;
  assign v_21332 = ~act_21144;
  assign v_21333 = v_21334 | v_21338;
  assign v_21334 = v_21335 | v_21336;
  assign v_21335 = mux_21335(v_20933);
  assign v_21336 = mux_21336(v_21337);
  assign v_21337 = ~v_20933;
  assign v_21338 = ~v_21141;
  assign v_21339 = v_21340 | v_21341;
  assign v_21340 = mux_21340(v_21143);
  assign v_21341 = mux_21341(v_21330);
  assign v_21342 = v_21343 & 1'h1;
  assign v_21343 = v_21344 & v_21345;
  assign v_21344 = ~act_20932;
  assign v_21345 = v_21346 | v_21350;
  assign v_21346 = v_21347 | v_21348;
  assign v_21347 = mux_21347(v_20497);
  assign v_21348 = mux_21348(v_21349);
  assign v_21349 = ~v_20497;
  assign v_21350 = ~v_20929;
  assign v_21351 = v_21352 | v_21353;
  assign v_21352 = mux_21352(v_20931);
  assign v_21353 = mux_21353(v_21342);
  assign v_21354 = v_21355 & 1'h1;
  assign v_21355 = v_21356 & v_21357;
  assign v_21356 = ~act_20496;
  assign v_21357 = v_21358 | v_21366;
  assign v_21358 = v_21359 | v_21364;
  assign v_21359 = mux_21359(v_21360);
  assign v_21360 = v_20493 & v_21361;
  assign v_21361 = v_21362 & 1'h1;
  assign v_21362 = v_21363 | 1'h0;
  assign v_21363 = ~v_20486;
  assign v_21364 = mux_21364(v_21365);
  assign v_21365 = ~v_21360;
  assign v_21366 = ~v_20493;
  assign v_21367 = v_21368 | v_21369;
  assign v_21368 = mux_21368(v_20495);
  assign v_21369 = mux_21369(v_21354);
  assign v_21371 = v_21372 | v_22231;
  assign v_21372 = act_21373 & 1'h1;
  assign act_21373 = v_21374 | v_21796;
  assign v_21374 = v_21375 & v_21797;
  assign v_21375 = v_21376 & v_21806;
  assign v_21376 = ~v_21377;
  assign v_21378 = v_21379 | v_21790;
  assign v_21379 = act_21380 & 1'h1;
  assign act_21380 = v_21381 | v_21579;
  assign v_21381 = v_21382 & v_21580;
  assign v_21382 = v_21383 & v_21589;
  assign v_21383 = ~v_21384;
  assign v_21385 = v_21386 | v_21573;
  assign v_21386 = act_21387 & 1'h1;
  assign act_21387 = v_21388 | v_21474;
  assign v_21388 = v_21389 & v_21475;
  assign v_21389 = v_21390 & v_21484;
  assign v_21390 = ~v_21391;
  assign v_21392 = v_21393 | v_21468;
  assign v_21393 = act_21394 & 1'h1;
  assign act_21394 = v_21395 | v_21425;
  assign v_21395 = v_21396 & v_21426;
  assign v_21396 = v_21397 & v_21435;
  assign v_21397 = ~v_21398;
  assign v_21399 = v_21400 | v_21419;
  assign v_21400 = act_21401 & 1'h1;
  assign act_21401 = v_21402 | v_21408;
  assign v_21402 = v_21403 & v_21409;
  assign v_21403 = v_21404 & vout_canPeek_21414;
  assign v_21404 = ~vout_canPeek_21405;
  pebbles_core
    pebbles_core_21405
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21406),
       .in0_consume_en(vin0_consume_en_21405),
       .out_canPeek(vout_canPeek_21405),
       .out_peek(vout_peek_21405));
  assign v_21406 = v_21407 | v_21412;
  assign v_21407 = mux_21407(v_21408);
  assign v_21408 = vout_canPeek_21405 & v_21409;
  assign v_21409 = v_21410 & 1'h1;
  assign v_21410 = v_21411 | 1'h0;
  assign v_21411 = ~v_21398;
  assign v_21412 = mux_21412(v_21413);
  assign v_21413 = ~v_21408;
  pebbles_core
    pebbles_core_21414
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21415),
       .in0_consume_en(vin0_consume_en_21414),
       .out_canPeek(vout_canPeek_21414),
       .out_peek(vout_peek_21414));
  assign v_21415 = v_21416 | v_21417;
  assign v_21416 = mux_21416(v_21402);
  assign v_21417 = mux_21417(v_21418);
  assign v_21418 = ~v_21402;
  assign v_21419 = v_21420 & 1'h1;
  assign v_21420 = v_21421 & v_21422;
  assign v_21421 = ~act_21401;
  assign v_21422 = v_21423 | v_21431;
  assign v_21423 = v_21424 | v_21429;
  assign v_21424 = mux_21424(v_21425);
  assign v_21425 = v_21398 & v_21426;
  assign v_21426 = v_21427 & 1'h1;
  assign v_21427 = v_21428 | 1'h0;
  assign v_21428 = ~v_21391;
  assign v_21429 = mux_21429(v_21430);
  assign v_21430 = ~v_21425;
  assign v_21431 = ~v_21398;
  assign v_21432 = v_21433 | v_21434;
  assign v_21433 = mux_21433(v_21400);
  assign v_21434 = mux_21434(v_21419);
  assign v_21436 = v_21437 | v_21456;
  assign v_21437 = act_21438 & 1'h1;
  assign act_21438 = v_21439 | v_21445;
  assign v_21439 = v_21440 & v_21446;
  assign v_21440 = v_21441 & vout_canPeek_21451;
  assign v_21441 = ~vout_canPeek_21442;
  pebbles_core
    pebbles_core_21442
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21443),
       .in0_consume_en(vin0_consume_en_21442),
       .out_canPeek(vout_canPeek_21442),
       .out_peek(vout_peek_21442));
  assign v_21443 = v_21444 | v_21449;
  assign v_21444 = mux_21444(v_21445);
  assign v_21445 = vout_canPeek_21442 & v_21446;
  assign v_21446 = v_21447 & 1'h1;
  assign v_21447 = v_21448 | 1'h0;
  assign v_21448 = ~v_21435;
  assign v_21449 = mux_21449(v_21450);
  assign v_21450 = ~v_21445;
  pebbles_core
    pebbles_core_21451
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21452),
       .in0_consume_en(vin0_consume_en_21451),
       .out_canPeek(vout_canPeek_21451),
       .out_peek(vout_peek_21451));
  assign v_21452 = v_21453 | v_21454;
  assign v_21453 = mux_21453(v_21439);
  assign v_21454 = mux_21454(v_21455);
  assign v_21455 = ~v_21439;
  assign v_21456 = v_21457 & 1'h1;
  assign v_21457 = v_21458 & v_21459;
  assign v_21458 = ~act_21438;
  assign v_21459 = v_21460 | v_21464;
  assign v_21460 = v_21461 | v_21462;
  assign v_21461 = mux_21461(v_21395);
  assign v_21462 = mux_21462(v_21463);
  assign v_21463 = ~v_21395;
  assign v_21464 = ~v_21435;
  assign v_21465 = v_21466 | v_21467;
  assign v_21466 = mux_21466(v_21437);
  assign v_21467 = mux_21467(v_21456);
  assign v_21468 = v_21469 & 1'h1;
  assign v_21469 = v_21470 & v_21471;
  assign v_21470 = ~act_21394;
  assign v_21471 = v_21472 | v_21480;
  assign v_21472 = v_21473 | v_21478;
  assign v_21473 = mux_21473(v_21474);
  assign v_21474 = v_21391 & v_21475;
  assign v_21475 = v_21476 & 1'h1;
  assign v_21476 = v_21477 | 1'h0;
  assign v_21477 = ~v_21384;
  assign v_21478 = mux_21478(v_21479);
  assign v_21479 = ~v_21474;
  assign v_21480 = ~v_21391;
  assign v_21481 = v_21482 | v_21483;
  assign v_21482 = mux_21482(v_21393);
  assign v_21483 = mux_21483(v_21468);
  assign v_21485 = v_21486 | v_21561;
  assign v_21486 = act_21487 & 1'h1;
  assign act_21487 = v_21488 | v_21518;
  assign v_21488 = v_21489 & v_21519;
  assign v_21489 = v_21490 & v_21528;
  assign v_21490 = ~v_21491;
  assign v_21492 = v_21493 | v_21512;
  assign v_21493 = act_21494 & 1'h1;
  assign act_21494 = v_21495 | v_21501;
  assign v_21495 = v_21496 & v_21502;
  assign v_21496 = v_21497 & vout_canPeek_21507;
  assign v_21497 = ~vout_canPeek_21498;
  pebbles_core
    pebbles_core_21498
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21499),
       .in0_consume_en(vin0_consume_en_21498),
       .out_canPeek(vout_canPeek_21498),
       .out_peek(vout_peek_21498));
  assign v_21499 = v_21500 | v_21505;
  assign v_21500 = mux_21500(v_21501);
  assign v_21501 = vout_canPeek_21498 & v_21502;
  assign v_21502 = v_21503 & 1'h1;
  assign v_21503 = v_21504 | 1'h0;
  assign v_21504 = ~v_21491;
  assign v_21505 = mux_21505(v_21506);
  assign v_21506 = ~v_21501;
  pebbles_core
    pebbles_core_21507
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21508),
       .in0_consume_en(vin0_consume_en_21507),
       .out_canPeek(vout_canPeek_21507),
       .out_peek(vout_peek_21507));
  assign v_21508 = v_21509 | v_21510;
  assign v_21509 = mux_21509(v_21495);
  assign v_21510 = mux_21510(v_21511);
  assign v_21511 = ~v_21495;
  assign v_21512 = v_21513 & 1'h1;
  assign v_21513 = v_21514 & v_21515;
  assign v_21514 = ~act_21494;
  assign v_21515 = v_21516 | v_21524;
  assign v_21516 = v_21517 | v_21522;
  assign v_21517 = mux_21517(v_21518);
  assign v_21518 = v_21491 & v_21519;
  assign v_21519 = v_21520 & 1'h1;
  assign v_21520 = v_21521 | 1'h0;
  assign v_21521 = ~v_21484;
  assign v_21522 = mux_21522(v_21523);
  assign v_21523 = ~v_21518;
  assign v_21524 = ~v_21491;
  assign v_21525 = v_21526 | v_21527;
  assign v_21526 = mux_21526(v_21493);
  assign v_21527 = mux_21527(v_21512);
  assign v_21529 = v_21530 | v_21549;
  assign v_21530 = act_21531 & 1'h1;
  assign act_21531 = v_21532 | v_21538;
  assign v_21532 = v_21533 & v_21539;
  assign v_21533 = v_21534 & vout_canPeek_21544;
  assign v_21534 = ~vout_canPeek_21535;
  pebbles_core
    pebbles_core_21535
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21536),
       .in0_consume_en(vin0_consume_en_21535),
       .out_canPeek(vout_canPeek_21535),
       .out_peek(vout_peek_21535));
  assign v_21536 = v_21537 | v_21542;
  assign v_21537 = mux_21537(v_21538);
  assign v_21538 = vout_canPeek_21535 & v_21539;
  assign v_21539 = v_21540 & 1'h1;
  assign v_21540 = v_21541 | 1'h0;
  assign v_21541 = ~v_21528;
  assign v_21542 = mux_21542(v_21543);
  assign v_21543 = ~v_21538;
  pebbles_core
    pebbles_core_21544
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21545),
       .in0_consume_en(vin0_consume_en_21544),
       .out_canPeek(vout_canPeek_21544),
       .out_peek(vout_peek_21544));
  assign v_21545 = v_21546 | v_21547;
  assign v_21546 = mux_21546(v_21532);
  assign v_21547 = mux_21547(v_21548);
  assign v_21548 = ~v_21532;
  assign v_21549 = v_21550 & 1'h1;
  assign v_21550 = v_21551 & v_21552;
  assign v_21551 = ~act_21531;
  assign v_21552 = v_21553 | v_21557;
  assign v_21553 = v_21554 | v_21555;
  assign v_21554 = mux_21554(v_21488);
  assign v_21555 = mux_21555(v_21556);
  assign v_21556 = ~v_21488;
  assign v_21557 = ~v_21528;
  assign v_21558 = v_21559 | v_21560;
  assign v_21559 = mux_21559(v_21530);
  assign v_21560 = mux_21560(v_21549);
  assign v_21561 = v_21562 & 1'h1;
  assign v_21562 = v_21563 & v_21564;
  assign v_21563 = ~act_21487;
  assign v_21564 = v_21565 | v_21569;
  assign v_21565 = v_21566 | v_21567;
  assign v_21566 = mux_21566(v_21388);
  assign v_21567 = mux_21567(v_21568);
  assign v_21568 = ~v_21388;
  assign v_21569 = ~v_21484;
  assign v_21570 = v_21571 | v_21572;
  assign v_21571 = mux_21571(v_21486);
  assign v_21572 = mux_21572(v_21561);
  assign v_21573 = v_21574 & 1'h1;
  assign v_21574 = v_21575 & v_21576;
  assign v_21575 = ~act_21387;
  assign v_21576 = v_21577 | v_21585;
  assign v_21577 = v_21578 | v_21583;
  assign v_21578 = mux_21578(v_21579);
  assign v_21579 = v_21384 & v_21580;
  assign v_21580 = v_21581 & 1'h1;
  assign v_21581 = v_21582 | 1'h0;
  assign v_21582 = ~v_21377;
  assign v_21583 = mux_21583(v_21584);
  assign v_21584 = ~v_21579;
  assign v_21585 = ~v_21384;
  assign v_21586 = v_21587 | v_21588;
  assign v_21587 = mux_21587(v_21386);
  assign v_21588 = mux_21588(v_21573);
  assign v_21590 = v_21591 | v_21778;
  assign v_21591 = act_21592 & 1'h1;
  assign act_21592 = v_21593 | v_21679;
  assign v_21593 = v_21594 & v_21680;
  assign v_21594 = v_21595 & v_21689;
  assign v_21595 = ~v_21596;
  assign v_21597 = v_21598 | v_21673;
  assign v_21598 = act_21599 & 1'h1;
  assign act_21599 = v_21600 | v_21630;
  assign v_21600 = v_21601 & v_21631;
  assign v_21601 = v_21602 & v_21640;
  assign v_21602 = ~v_21603;
  assign v_21604 = v_21605 | v_21624;
  assign v_21605 = act_21606 & 1'h1;
  assign act_21606 = v_21607 | v_21613;
  assign v_21607 = v_21608 & v_21614;
  assign v_21608 = v_21609 & vout_canPeek_21619;
  assign v_21609 = ~vout_canPeek_21610;
  pebbles_core
    pebbles_core_21610
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21611),
       .in0_consume_en(vin0_consume_en_21610),
       .out_canPeek(vout_canPeek_21610),
       .out_peek(vout_peek_21610));
  assign v_21611 = v_21612 | v_21617;
  assign v_21612 = mux_21612(v_21613);
  assign v_21613 = vout_canPeek_21610 & v_21614;
  assign v_21614 = v_21615 & 1'h1;
  assign v_21615 = v_21616 | 1'h0;
  assign v_21616 = ~v_21603;
  assign v_21617 = mux_21617(v_21618);
  assign v_21618 = ~v_21613;
  pebbles_core
    pebbles_core_21619
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21620),
       .in0_consume_en(vin0_consume_en_21619),
       .out_canPeek(vout_canPeek_21619),
       .out_peek(vout_peek_21619));
  assign v_21620 = v_21621 | v_21622;
  assign v_21621 = mux_21621(v_21607);
  assign v_21622 = mux_21622(v_21623);
  assign v_21623 = ~v_21607;
  assign v_21624 = v_21625 & 1'h1;
  assign v_21625 = v_21626 & v_21627;
  assign v_21626 = ~act_21606;
  assign v_21627 = v_21628 | v_21636;
  assign v_21628 = v_21629 | v_21634;
  assign v_21629 = mux_21629(v_21630);
  assign v_21630 = v_21603 & v_21631;
  assign v_21631 = v_21632 & 1'h1;
  assign v_21632 = v_21633 | 1'h0;
  assign v_21633 = ~v_21596;
  assign v_21634 = mux_21634(v_21635);
  assign v_21635 = ~v_21630;
  assign v_21636 = ~v_21603;
  assign v_21637 = v_21638 | v_21639;
  assign v_21638 = mux_21638(v_21605);
  assign v_21639 = mux_21639(v_21624);
  assign v_21641 = v_21642 | v_21661;
  assign v_21642 = act_21643 & 1'h1;
  assign act_21643 = v_21644 | v_21650;
  assign v_21644 = v_21645 & v_21651;
  assign v_21645 = v_21646 & vout_canPeek_21656;
  assign v_21646 = ~vout_canPeek_21647;
  pebbles_core
    pebbles_core_21647
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21648),
       .in0_consume_en(vin0_consume_en_21647),
       .out_canPeek(vout_canPeek_21647),
       .out_peek(vout_peek_21647));
  assign v_21648 = v_21649 | v_21654;
  assign v_21649 = mux_21649(v_21650);
  assign v_21650 = vout_canPeek_21647 & v_21651;
  assign v_21651 = v_21652 & 1'h1;
  assign v_21652 = v_21653 | 1'h0;
  assign v_21653 = ~v_21640;
  assign v_21654 = mux_21654(v_21655);
  assign v_21655 = ~v_21650;
  pebbles_core
    pebbles_core_21656
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21657),
       .in0_consume_en(vin0_consume_en_21656),
       .out_canPeek(vout_canPeek_21656),
       .out_peek(vout_peek_21656));
  assign v_21657 = v_21658 | v_21659;
  assign v_21658 = mux_21658(v_21644);
  assign v_21659 = mux_21659(v_21660);
  assign v_21660 = ~v_21644;
  assign v_21661 = v_21662 & 1'h1;
  assign v_21662 = v_21663 & v_21664;
  assign v_21663 = ~act_21643;
  assign v_21664 = v_21665 | v_21669;
  assign v_21665 = v_21666 | v_21667;
  assign v_21666 = mux_21666(v_21600);
  assign v_21667 = mux_21667(v_21668);
  assign v_21668 = ~v_21600;
  assign v_21669 = ~v_21640;
  assign v_21670 = v_21671 | v_21672;
  assign v_21671 = mux_21671(v_21642);
  assign v_21672 = mux_21672(v_21661);
  assign v_21673 = v_21674 & 1'h1;
  assign v_21674 = v_21675 & v_21676;
  assign v_21675 = ~act_21599;
  assign v_21676 = v_21677 | v_21685;
  assign v_21677 = v_21678 | v_21683;
  assign v_21678 = mux_21678(v_21679);
  assign v_21679 = v_21596 & v_21680;
  assign v_21680 = v_21681 & 1'h1;
  assign v_21681 = v_21682 | 1'h0;
  assign v_21682 = ~v_21589;
  assign v_21683 = mux_21683(v_21684);
  assign v_21684 = ~v_21679;
  assign v_21685 = ~v_21596;
  assign v_21686 = v_21687 | v_21688;
  assign v_21687 = mux_21687(v_21598);
  assign v_21688 = mux_21688(v_21673);
  assign v_21690 = v_21691 | v_21766;
  assign v_21691 = act_21692 & 1'h1;
  assign act_21692 = v_21693 | v_21723;
  assign v_21693 = v_21694 & v_21724;
  assign v_21694 = v_21695 & v_21733;
  assign v_21695 = ~v_21696;
  assign v_21697 = v_21698 | v_21717;
  assign v_21698 = act_21699 & 1'h1;
  assign act_21699 = v_21700 | v_21706;
  assign v_21700 = v_21701 & v_21707;
  assign v_21701 = v_21702 & vout_canPeek_21712;
  assign v_21702 = ~vout_canPeek_21703;
  pebbles_core
    pebbles_core_21703
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21704),
       .in0_consume_en(vin0_consume_en_21703),
       .out_canPeek(vout_canPeek_21703),
       .out_peek(vout_peek_21703));
  assign v_21704 = v_21705 | v_21710;
  assign v_21705 = mux_21705(v_21706);
  assign v_21706 = vout_canPeek_21703 & v_21707;
  assign v_21707 = v_21708 & 1'h1;
  assign v_21708 = v_21709 | 1'h0;
  assign v_21709 = ~v_21696;
  assign v_21710 = mux_21710(v_21711);
  assign v_21711 = ~v_21706;
  pebbles_core
    pebbles_core_21712
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21713),
       .in0_consume_en(vin0_consume_en_21712),
       .out_canPeek(vout_canPeek_21712),
       .out_peek(vout_peek_21712));
  assign v_21713 = v_21714 | v_21715;
  assign v_21714 = mux_21714(v_21700);
  assign v_21715 = mux_21715(v_21716);
  assign v_21716 = ~v_21700;
  assign v_21717 = v_21718 & 1'h1;
  assign v_21718 = v_21719 & v_21720;
  assign v_21719 = ~act_21699;
  assign v_21720 = v_21721 | v_21729;
  assign v_21721 = v_21722 | v_21727;
  assign v_21722 = mux_21722(v_21723);
  assign v_21723 = v_21696 & v_21724;
  assign v_21724 = v_21725 & 1'h1;
  assign v_21725 = v_21726 | 1'h0;
  assign v_21726 = ~v_21689;
  assign v_21727 = mux_21727(v_21728);
  assign v_21728 = ~v_21723;
  assign v_21729 = ~v_21696;
  assign v_21730 = v_21731 | v_21732;
  assign v_21731 = mux_21731(v_21698);
  assign v_21732 = mux_21732(v_21717);
  assign v_21734 = v_21735 | v_21754;
  assign v_21735 = act_21736 & 1'h1;
  assign act_21736 = v_21737 | v_21743;
  assign v_21737 = v_21738 & v_21744;
  assign v_21738 = v_21739 & vout_canPeek_21749;
  assign v_21739 = ~vout_canPeek_21740;
  pebbles_core
    pebbles_core_21740
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21741),
       .in0_consume_en(vin0_consume_en_21740),
       .out_canPeek(vout_canPeek_21740),
       .out_peek(vout_peek_21740));
  assign v_21741 = v_21742 | v_21747;
  assign v_21742 = mux_21742(v_21743);
  assign v_21743 = vout_canPeek_21740 & v_21744;
  assign v_21744 = v_21745 & 1'h1;
  assign v_21745 = v_21746 | 1'h0;
  assign v_21746 = ~v_21733;
  assign v_21747 = mux_21747(v_21748);
  assign v_21748 = ~v_21743;
  pebbles_core
    pebbles_core_21749
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21750),
       .in0_consume_en(vin0_consume_en_21749),
       .out_canPeek(vout_canPeek_21749),
       .out_peek(vout_peek_21749));
  assign v_21750 = v_21751 | v_21752;
  assign v_21751 = mux_21751(v_21737);
  assign v_21752 = mux_21752(v_21753);
  assign v_21753 = ~v_21737;
  assign v_21754 = v_21755 & 1'h1;
  assign v_21755 = v_21756 & v_21757;
  assign v_21756 = ~act_21736;
  assign v_21757 = v_21758 | v_21762;
  assign v_21758 = v_21759 | v_21760;
  assign v_21759 = mux_21759(v_21693);
  assign v_21760 = mux_21760(v_21761);
  assign v_21761 = ~v_21693;
  assign v_21762 = ~v_21733;
  assign v_21763 = v_21764 | v_21765;
  assign v_21764 = mux_21764(v_21735);
  assign v_21765 = mux_21765(v_21754);
  assign v_21766 = v_21767 & 1'h1;
  assign v_21767 = v_21768 & v_21769;
  assign v_21768 = ~act_21692;
  assign v_21769 = v_21770 | v_21774;
  assign v_21770 = v_21771 | v_21772;
  assign v_21771 = mux_21771(v_21593);
  assign v_21772 = mux_21772(v_21773);
  assign v_21773 = ~v_21593;
  assign v_21774 = ~v_21689;
  assign v_21775 = v_21776 | v_21777;
  assign v_21776 = mux_21776(v_21691);
  assign v_21777 = mux_21777(v_21766);
  assign v_21778 = v_21779 & 1'h1;
  assign v_21779 = v_21780 & v_21781;
  assign v_21780 = ~act_21592;
  assign v_21781 = v_21782 | v_21786;
  assign v_21782 = v_21783 | v_21784;
  assign v_21783 = mux_21783(v_21381);
  assign v_21784 = mux_21784(v_21785);
  assign v_21785 = ~v_21381;
  assign v_21786 = ~v_21589;
  assign v_21787 = v_21788 | v_21789;
  assign v_21788 = mux_21788(v_21591);
  assign v_21789 = mux_21789(v_21778);
  assign v_21790 = v_21791 & 1'h1;
  assign v_21791 = v_21792 & v_21793;
  assign v_21792 = ~act_21380;
  assign v_21793 = v_21794 | v_21802;
  assign v_21794 = v_21795 | v_21800;
  assign v_21795 = mux_21795(v_21796);
  assign v_21796 = v_21377 & v_21797;
  assign v_21797 = v_21798 & 1'h1;
  assign v_21798 = v_21799 | 1'h0;
  assign v_21799 = ~v_21370;
  assign v_21800 = mux_21800(v_21801);
  assign v_21801 = ~v_21796;
  assign v_21802 = ~v_21377;
  assign v_21803 = v_21804 | v_21805;
  assign v_21804 = mux_21804(v_21379);
  assign v_21805 = mux_21805(v_21790);
  assign v_21807 = v_21808 | v_22219;
  assign v_21808 = act_21809 & 1'h1;
  assign act_21809 = v_21810 | v_22008;
  assign v_21810 = v_21811 & v_22009;
  assign v_21811 = v_21812 & v_22018;
  assign v_21812 = ~v_21813;
  assign v_21814 = v_21815 | v_22002;
  assign v_21815 = act_21816 & 1'h1;
  assign act_21816 = v_21817 | v_21903;
  assign v_21817 = v_21818 & v_21904;
  assign v_21818 = v_21819 & v_21913;
  assign v_21819 = ~v_21820;
  assign v_21821 = v_21822 | v_21897;
  assign v_21822 = act_21823 & 1'h1;
  assign act_21823 = v_21824 | v_21854;
  assign v_21824 = v_21825 & v_21855;
  assign v_21825 = v_21826 & v_21864;
  assign v_21826 = ~v_21827;
  assign v_21828 = v_21829 | v_21848;
  assign v_21829 = act_21830 & 1'h1;
  assign act_21830 = v_21831 | v_21837;
  assign v_21831 = v_21832 & v_21838;
  assign v_21832 = v_21833 & vout_canPeek_21843;
  assign v_21833 = ~vout_canPeek_21834;
  pebbles_core
    pebbles_core_21834
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21835),
       .in0_consume_en(vin0_consume_en_21834),
       .out_canPeek(vout_canPeek_21834),
       .out_peek(vout_peek_21834));
  assign v_21835 = v_21836 | v_21841;
  assign v_21836 = mux_21836(v_21837);
  assign v_21837 = vout_canPeek_21834 & v_21838;
  assign v_21838 = v_21839 & 1'h1;
  assign v_21839 = v_21840 | 1'h0;
  assign v_21840 = ~v_21827;
  assign v_21841 = mux_21841(v_21842);
  assign v_21842 = ~v_21837;
  pebbles_core
    pebbles_core_21843
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21844),
       .in0_consume_en(vin0_consume_en_21843),
       .out_canPeek(vout_canPeek_21843),
       .out_peek(vout_peek_21843));
  assign v_21844 = v_21845 | v_21846;
  assign v_21845 = mux_21845(v_21831);
  assign v_21846 = mux_21846(v_21847);
  assign v_21847 = ~v_21831;
  assign v_21848 = v_21849 & 1'h1;
  assign v_21849 = v_21850 & v_21851;
  assign v_21850 = ~act_21830;
  assign v_21851 = v_21852 | v_21860;
  assign v_21852 = v_21853 | v_21858;
  assign v_21853 = mux_21853(v_21854);
  assign v_21854 = v_21827 & v_21855;
  assign v_21855 = v_21856 & 1'h1;
  assign v_21856 = v_21857 | 1'h0;
  assign v_21857 = ~v_21820;
  assign v_21858 = mux_21858(v_21859);
  assign v_21859 = ~v_21854;
  assign v_21860 = ~v_21827;
  assign v_21861 = v_21862 | v_21863;
  assign v_21862 = mux_21862(v_21829);
  assign v_21863 = mux_21863(v_21848);
  assign v_21865 = v_21866 | v_21885;
  assign v_21866 = act_21867 & 1'h1;
  assign act_21867 = v_21868 | v_21874;
  assign v_21868 = v_21869 & v_21875;
  assign v_21869 = v_21870 & vout_canPeek_21880;
  assign v_21870 = ~vout_canPeek_21871;
  pebbles_core
    pebbles_core_21871
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21872),
       .in0_consume_en(vin0_consume_en_21871),
       .out_canPeek(vout_canPeek_21871),
       .out_peek(vout_peek_21871));
  assign v_21872 = v_21873 | v_21878;
  assign v_21873 = mux_21873(v_21874);
  assign v_21874 = vout_canPeek_21871 & v_21875;
  assign v_21875 = v_21876 & 1'h1;
  assign v_21876 = v_21877 | 1'h0;
  assign v_21877 = ~v_21864;
  assign v_21878 = mux_21878(v_21879);
  assign v_21879 = ~v_21874;
  pebbles_core
    pebbles_core_21880
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21881),
       .in0_consume_en(vin0_consume_en_21880),
       .out_canPeek(vout_canPeek_21880),
       .out_peek(vout_peek_21880));
  assign v_21881 = v_21882 | v_21883;
  assign v_21882 = mux_21882(v_21868);
  assign v_21883 = mux_21883(v_21884);
  assign v_21884 = ~v_21868;
  assign v_21885 = v_21886 & 1'h1;
  assign v_21886 = v_21887 & v_21888;
  assign v_21887 = ~act_21867;
  assign v_21888 = v_21889 | v_21893;
  assign v_21889 = v_21890 | v_21891;
  assign v_21890 = mux_21890(v_21824);
  assign v_21891 = mux_21891(v_21892);
  assign v_21892 = ~v_21824;
  assign v_21893 = ~v_21864;
  assign v_21894 = v_21895 | v_21896;
  assign v_21895 = mux_21895(v_21866);
  assign v_21896 = mux_21896(v_21885);
  assign v_21897 = v_21898 & 1'h1;
  assign v_21898 = v_21899 & v_21900;
  assign v_21899 = ~act_21823;
  assign v_21900 = v_21901 | v_21909;
  assign v_21901 = v_21902 | v_21907;
  assign v_21902 = mux_21902(v_21903);
  assign v_21903 = v_21820 & v_21904;
  assign v_21904 = v_21905 & 1'h1;
  assign v_21905 = v_21906 | 1'h0;
  assign v_21906 = ~v_21813;
  assign v_21907 = mux_21907(v_21908);
  assign v_21908 = ~v_21903;
  assign v_21909 = ~v_21820;
  assign v_21910 = v_21911 | v_21912;
  assign v_21911 = mux_21911(v_21822);
  assign v_21912 = mux_21912(v_21897);
  assign v_21914 = v_21915 | v_21990;
  assign v_21915 = act_21916 & 1'h1;
  assign act_21916 = v_21917 | v_21947;
  assign v_21917 = v_21918 & v_21948;
  assign v_21918 = v_21919 & v_21957;
  assign v_21919 = ~v_21920;
  assign v_21921 = v_21922 | v_21941;
  assign v_21922 = act_21923 & 1'h1;
  assign act_21923 = v_21924 | v_21930;
  assign v_21924 = v_21925 & v_21931;
  assign v_21925 = v_21926 & vout_canPeek_21936;
  assign v_21926 = ~vout_canPeek_21927;
  pebbles_core
    pebbles_core_21927
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21928),
       .in0_consume_en(vin0_consume_en_21927),
       .out_canPeek(vout_canPeek_21927),
       .out_peek(vout_peek_21927));
  assign v_21928 = v_21929 | v_21934;
  assign v_21929 = mux_21929(v_21930);
  assign v_21930 = vout_canPeek_21927 & v_21931;
  assign v_21931 = v_21932 & 1'h1;
  assign v_21932 = v_21933 | 1'h0;
  assign v_21933 = ~v_21920;
  assign v_21934 = mux_21934(v_21935);
  assign v_21935 = ~v_21930;
  pebbles_core
    pebbles_core_21936
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21937),
       .in0_consume_en(vin0_consume_en_21936),
       .out_canPeek(vout_canPeek_21936),
       .out_peek(vout_peek_21936));
  assign v_21937 = v_21938 | v_21939;
  assign v_21938 = mux_21938(v_21924);
  assign v_21939 = mux_21939(v_21940);
  assign v_21940 = ~v_21924;
  assign v_21941 = v_21942 & 1'h1;
  assign v_21942 = v_21943 & v_21944;
  assign v_21943 = ~act_21923;
  assign v_21944 = v_21945 | v_21953;
  assign v_21945 = v_21946 | v_21951;
  assign v_21946 = mux_21946(v_21947);
  assign v_21947 = v_21920 & v_21948;
  assign v_21948 = v_21949 & 1'h1;
  assign v_21949 = v_21950 | 1'h0;
  assign v_21950 = ~v_21913;
  assign v_21951 = mux_21951(v_21952);
  assign v_21952 = ~v_21947;
  assign v_21953 = ~v_21920;
  assign v_21954 = v_21955 | v_21956;
  assign v_21955 = mux_21955(v_21922);
  assign v_21956 = mux_21956(v_21941);
  assign v_21958 = v_21959 | v_21978;
  assign v_21959 = act_21960 & 1'h1;
  assign act_21960 = v_21961 | v_21967;
  assign v_21961 = v_21962 & v_21968;
  assign v_21962 = v_21963 & vout_canPeek_21973;
  assign v_21963 = ~vout_canPeek_21964;
  pebbles_core
    pebbles_core_21964
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21965),
       .in0_consume_en(vin0_consume_en_21964),
       .out_canPeek(vout_canPeek_21964),
       .out_peek(vout_peek_21964));
  assign v_21965 = v_21966 | v_21971;
  assign v_21966 = mux_21966(v_21967);
  assign v_21967 = vout_canPeek_21964 & v_21968;
  assign v_21968 = v_21969 & 1'h1;
  assign v_21969 = v_21970 | 1'h0;
  assign v_21970 = ~v_21957;
  assign v_21971 = mux_21971(v_21972);
  assign v_21972 = ~v_21967;
  pebbles_core
    pebbles_core_21973
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_21974),
       .in0_consume_en(vin0_consume_en_21973),
       .out_canPeek(vout_canPeek_21973),
       .out_peek(vout_peek_21973));
  assign v_21974 = v_21975 | v_21976;
  assign v_21975 = mux_21975(v_21961);
  assign v_21976 = mux_21976(v_21977);
  assign v_21977 = ~v_21961;
  assign v_21978 = v_21979 & 1'h1;
  assign v_21979 = v_21980 & v_21981;
  assign v_21980 = ~act_21960;
  assign v_21981 = v_21982 | v_21986;
  assign v_21982 = v_21983 | v_21984;
  assign v_21983 = mux_21983(v_21917);
  assign v_21984 = mux_21984(v_21985);
  assign v_21985 = ~v_21917;
  assign v_21986 = ~v_21957;
  assign v_21987 = v_21988 | v_21989;
  assign v_21988 = mux_21988(v_21959);
  assign v_21989 = mux_21989(v_21978);
  assign v_21990 = v_21991 & 1'h1;
  assign v_21991 = v_21992 & v_21993;
  assign v_21992 = ~act_21916;
  assign v_21993 = v_21994 | v_21998;
  assign v_21994 = v_21995 | v_21996;
  assign v_21995 = mux_21995(v_21817);
  assign v_21996 = mux_21996(v_21997);
  assign v_21997 = ~v_21817;
  assign v_21998 = ~v_21913;
  assign v_21999 = v_22000 | v_22001;
  assign v_22000 = mux_22000(v_21915);
  assign v_22001 = mux_22001(v_21990);
  assign v_22002 = v_22003 & 1'h1;
  assign v_22003 = v_22004 & v_22005;
  assign v_22004 = ~act_21816;
  assign v_22005 = v_22006 | v_22014;
  assign v_22006 = v_22007 | v_22012;
  assign v_22007 = mux_22007(v_22008);
  assign v_22008 = v_21813 & v_22009;
  assign v_22009 = v_22010 & 1'h1;
  assign v_22010 = v_22011 | 1'h0;
  assign v_22011 = ~v_21806;
  assign v_22012 = mux_22012(v_22013);
  assign v_22013 = ~v_22008;
  assign v_22014 = ~v_21813;
  assign v_22015 = v_22016 | v_22017;
  assign v_22016 = mux_22016(v_21815);
  assign v_22017 = mux_22017(v_22002);
  assign v_22019 = v_22020 | v_22207;
  assign v_22020 = act_22021 & 1'h1;
  assign act_22021 = v_22022 | v_22108;
  assign v_22022 = v_22023 & v_22109;
  assign v_22023 = v_22024 & v_22118;
  assign v_22024 = ~v_22025;
  assign v_22026 = v_22027 | v_22102;
  assign v_22027 = act_22028 & 1'h1;
  assign act_22028 = v_22029 | v_22059;
  assign v_22029 = v_22030 & v_22060;
  assign v_22030 = v_22031 & v_22069;
  assign v_22031 = ~v_22032;
  assign v_22033 = v_22034 | v_22053;
  assign v_22034 = act_22035 & 1'h1;
  assign act_22035 = v_22036 | v_22042;
  assign v_22036 = v_22037 & v_22043;
  assign v_22037 = v_22038 & vout_canPeek_22048;
  assign v_22038 = ~vout_canPeek_22039;
  pebbles_core
    pebbles_core_22039
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_22040),
       .in0_consume_en(vin0_consume_en_22039),
       .out_canPeek(vout_canPeek_22039),
       .out_peek(vout_peek_22039));
  assign v_22040 = v_22041 | v_22046;
  assign v_22041 = mux_22041(v_22042);
  assign v_22042 = vout_canPeek_22039 & v_22043;
  assign v_22043 = v_22044 & 1'h1;
  assign v_22044 = v_22045 | 1'h0;
  assign v_22045 = ~v_22032;
  assign v_22046 = mux_22046(v_22047);
  assign v_22047 = ~v_22042;
  pebbles_core
    pebbles_core_22048
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_22049),
       .in0_consume_en(vin0_consume_en_22048),
       .out_canPeek(vout_canPeek_22048),
       .out_peek(vout_peek_22048));
  assign v_22049 = v_22050 | v_22051;
  assign v_22050 = mux_22050(v_22036);
  assign v_22051 = mux_22051(v_22052);
  assign v_22052 = ~v_22036;
  assign v_22053 = v_22054 & 1'h1;
  assign v_22054 = v_22055 & v_22056;
  assign v_22055 = ~act_22035;
  assign v_22056 = v_22057 | v_22065;
  assign v_22057 = v_22058 | v_22063;
  assign v_22058 = mux_22058(v_22059);
  assign v_22059 = v_22032 & v_22060;
  assign v_22060 = v_22061 & 1'h1;
  assign v_22061 = v_22062 | 1'h0;
  assign v_22062 = ~v_22025;
  assign v_22063 = mux_22063(v_22064);
  assign v_22064 = ~v_22059;
  assign v_22065 = ~v_22032;
  assign v_22066 = v_22067 | v_22068;
  assign v_22067 = mux_22067(v_22034);
  assign v_22068 = mux_22068(v_22053);
  assign v_22070 = v_22071 | v_22090;
  assign v_22071 = act_22072 & 1'h1;
  assign act_22072 = v_22073 | v_22079;
  assign v_22073 = v_22074 & v_22080;
  assign v_22074 = v_22075 & vout_canPeek_22085;
  assign v_22075 = ~vout_canPeek_22076;
  pebbles_core
    pebbles_core_22076
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_22077),
       .in0_consume_en(vin0_consume_en_22076),
       .out_canPeek(vout_canPeek_22076),
       .out_peek(vout_peek_22076));
  assign v_22077 = v_22078 | v_22083;
  assign v_22078 = mux_22078(v_22079);
  assign v_22079 = vout_canPeek_22076 & v_22080;
  assign v_22080 = v_22081 & 1'h1;
  assign v_22081 = v_22082 | 1'h0;
  assign v_22082 = ~v_22069;
  assign v_22083 = mux_22083(v_22084);
  assign v_22084 = ~v_22079;
  pebbles_core
    pebbles_core_22085
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_22086),
       .in0_consume_en(vin0_consume_en_22085),
       .out_canPeek(vout_canPeek_22085),
       .out_peek(vout_peek_22085));
  assign v_22086 = v_22087 | v_22088;
  assign v_22087 = mux_22087(v_22073);
  assign v_22088 = mux_22088(v_22089);
  assign v_22089 = ~v_22073;
  assign v_22090 = v_22091 & 1'h1;
  assign v_22091 = v_22092 & v_22093;
  assign v_22092 = ~act_22072;
  assign v_22093 = v_22094 | v_22098;
  assign v_22094 = v_22095 | v_22096;
  assign v_22095 = mux_22095(v_22029);
  assign v_22096 = mux_22096(v_22097);
  assign v_22097 = ~v_22029;
  assign v_22098 = ~v_22069;
  assign v_22099 = v_22100 | v_22101;
  assign v_22100 = mux_22100(v_22071);
  assign v_22101 = mux_22101(v_22090);
  assign v_22102 = v_22103 & 1'h1;
  assign v_22103 = v_22104 & v_22105;
  assign v_22104 = ~act_22028;
  assign v_22105 = v_22106 | v_22114;
  assign v_22106 = v_22107 | v_22112;
  assign v_22107 = mux_22107(v_22108);
  assign v_22108 = v_22025 & v_22109;
  assign v_22109 = v_22110 & 1'h1;
  assign v_22110 = v_22111 | 1'h0;
  assign v_22111 = ~v_22018;
  assign v_22112 = mux_22112(v_22113);
  assign v_22113 = ~v_22108;
  assign v_22114 = ~v_22025;
  assign v_22115 = v_22116 | v_22117;
  assign v_22116 = mux_22116(v_22027);
  assign v_22117 = mux_22117(v_22102);
  assign v_22119 = v_22120 | v_22195;
  assign v_22120 = act_22121 & 1'h1;
  assign act_22121 = v_22122 | v_22152;
  assign v_22122 = v_22123 & v_22153;
  assign v_22123 = v_22124 & v_22162;
  assign v_22124 = ~v_22125;
  assign v_22126 = v_22127 | v_22146;
  assign v_22127 = act_22128 & 1'h1;
  assign act_22128 = v_22129 | v_22135;
  assign v_22129 = v_22130 & v_22136;
  assign v_22130 = v_22131 & vout_canPeek_22141;
  assign v_22131 = ~vout_canPeek_22132;
  pebbles_core
    pebbles_core_22132
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_22133),
       .in0_consume_en(vin0_consume_en_22132),
       .out_canPeek(vout_canPeek_22132),
       .out_peek(vout_peek_22132));
  assign v_22133 = v_22134 | v_22139;
  assign v_22134 = mux_22134(v_22135);
  assign v_22135 = vout_canPeek_22132 & v_22136;
  assign v_22136 = v_22137 & 1'h1;
  assign v_22137 = v_22138 | 1'h0;
  assign v_22138 = ~v_22125;
  assign v_22139 = mux_22139(v_22140);
  assign v_22140 = ~v_22135;
  pebbles_core
    pebbles_core_22141
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_22142),
       .in0_consume_en(vin0_consume_en_22141),
       .out_canPeek(vout_canPeek_22141),
       .out_peek(vout_peek_22141));
  assign v_22142 = v_22143 | v_22144;
  assign v_22143 = mux_22143(v_22129);
  assign v_22144 = mux_22144(v_22145);
  assign v_22145 = ~v_22129;
  assign v_22146 = v_22147 & 1'h1;
  assign v_22147 = v_22148 & v_22149;
  assign v_22148 = ~act_22128;
  assign v_22149 = v_22150 | v_22158;
  assign v_22150 = v_22151 | v_22156;
  assign v_22151 = mux_22151(v_22152);
  assign v_22152 = v_22125 & v_22153;
  assign v_22153 = v_22154 & 1'h1;
  assign v_22154 = v_22155 | 1'h0;
  assign v_22155 = ~v_22118;
  assign v_22156 = mux_22156(v_22157);
  assign v_22157 = ~v_22152;
  assign v_22158 = ~v_22125;
  assign v_22159 = v_22160 | v_22161;
  assign v_22160 = mux_22160(v_22127);
  assign v_22161 = mux_22161(v_22146);
  assign v_22163 = v_22164 | v_22183;
  assign v_22164 = act_22165 & 1'h1;
  assign act_22165 = v_22166 | v_22172;
  assign v_22166 = v_22167 & v_22173;
  assign v_22167 = v_22168 & vout_canPeek_22178;
  assign v_22168 = ~vout_canPeek_22169;
  pebbles_core
    pebbles_core_22169
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_22170),
       .in0_consume_en(vin0_consume_en_22169),
       .out_canPeek(vout_canPeek_22169),
       .out_peek(vout_peek_22169));
  assign v_22170 = v_22171 | v_22176;
  assign v_22171 = mux_22171(v_22172);
  assign v_22172 = vout_canPeek_22169 & v_22173;
  assign v_22173 = v_22174 & 1'h1;
  assign v_22174 = v_22175 | 1'h0;
  assign v_22175 = ~v_22162;
  assign v_22176 = mux_22176(v_22177);
  assign v_22177 = ~v_22172;
  pebbles_core
    pebbles_core_22178
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_22179),
       .in0_consume_en(vin0_consume_en_22178),
       .out_canPeek(vout_canPeek_22178),
       .out_peek(vout_peek_22178));
  assign v_22179 = v_22180 | v_22181;
  assign v_22180 = mux_22180(v_22166);
  assign v_22181 = mux_22181(v_22182);
  assign v_22182 = ~v_22166;
  assign v_22183 = v_22184 & 1'h1;
  assign v_22184 = v_22185 & v_22186;
  assign v_22185 = ~act_22165;
  assign v_22186 = v_22187 | v_22191;
  assign v_22187 = v_22188 | v_22189;
  assign v_22188 = mux_22188(v_22122);
  assign v_22189 = mux_22189(v_22190);
  assign v_22190 = ~v_22122;
  assign v_22191 = ~v_22162;
  assign v_22192 = v_22193 | v_22194;
  assign v_22193 = mux_22193(v_22164);
  assign v_22194 = mux_22194(v_22183);
  assign v_22195 = v_22196 & 1'h1;
  assign v_22196 = v_22197 & v_22198;
  assign v_22197 = ~act_22121;
  assign v_22198 = v_22199 | v_22203;
  assign v_22199 = v_22200 | v_22201;
  assign v_22200 = mux_22200(v_22022);
  assign v_22201 = mux_22201(v_22202);
  assign v_22202 = ~v_22022;
  assign v_22203 = ~v_22118;
  assign v_22204 = v_22205 | v_22206;
  assign v_22205 = mux_22205(v_22120);
  assign v_22206 = mux_22206(v_22195);
  assign v_22207 = v_22208 & 1'h1;
  assign v_22208 = v_22209 & v_22210;
  assign v_22209 = ~act_22021;
  assign v_22210 = v_22211 | v_22215;
  assign v_22211 = v_22212 | v_22213;
  assign v_22212 = mux_22212(v_21810);
  assign v_22213 = mux_22213(v_22214);
  assign v_22214 = ~v_21810;
  assign v_22215 = ~v_22018;
  assign v_22216 = v_22217 | v_22218;
  assign v_22217 = mux_22217(v_22020);
  assign v_22218 = mux_22218(v_22207);
  assign v_22219 = v_22220 & 1'h1;
  assign v_22220 = v_22221 & v_22222;
  assign v_22221 = ~act_21809;
  assign v_22222 = v_22223 | v_22227;
  assign v_22223 = v_22224 | v_22225;
  assign v_22224 = mux_22224(v_21374);
  assign v_22225 = mux_22225(v_22226);
  assign v_22226 = ~v_21374;
  assign v_22227 = ~v_21806;
  assign v_22228 = v_22229 | v_22230;
  assign v_22229 = mux_22229(v_21808);
  assign v_22230 = mux_22230(v_22219);
  assign v_22231 = v_22232 & 1'h1;
  assign v_22232 = v_22233 & v_22234;
  assign v_22233 = ~act_21373;
  assign v_22234 = v_22235 | v_22239;
  assign v_22235 = v_22236 | v_22237;
  assign v_22236 = mux_22236(v_20490);
  assign v_22237 = mux_22237(v_22238);
  assign v_22238 = ~v_20490;
  assign v_22239 = ~v_21370;
  assign v_22240 = v_22241 | v_22242;
  assign v_22241 = mux_22241(v_21372);
  assign v_22242 = mux_22242(v_22231);
  assign v_22243 = v_22244 & 1'h1;
  assign v_22244 = v_22245 & v_22246;
  assign v_22245 = ~act_20489;
  assign v_22246 = v_22247 | v_22251;
  assign v_22247 = v_22248 | v_22249;
  assign v_22248 = mux_22248(v_18710);
  assign v_22249 = mux_22249(v_22250);
  assign v_22250 = ~v_18710;
  assign v_22251 = ~v_20486;
  assign v_22252 = v_22253 | v_22254;
  assign v_22253 = mux_22253(v_20488);
  assign v_22254 = mux_22254(v_22243);
  assign v_22255 = v_22256 & 1'h1;
  assign v_22256 = v_22257 & v_22258;
  assign v_22257 = ~act_18709;
  assign v_22258 = v_22259 | v_22263;
  assign v_22259 = v_22260 | v_22261;
  assign v_22260 = mux_22260(v_15138);
  assign v_22261 = mux_22261(v_22262);
  assign v_22262 = ~v_15138;
  assign v_22263 = ~v_18706;
  assign v_22264 = v_22265 | v_22266;
  assign v_22265 = mux_22265(v_18708);
  assign v_22266 = mux_22266(v_22255);
  assign v_22267 = v_22268 & 1'h1;
  assign v_22268 = v_22269 & v_22270;
  assign v_22269 = ~act_15137;
  assign v_22270 = v_22271 | v_22275;
  assign v_22271 = v_22272 | v_22273;
  assign v_22272 = mux_22272(v_7982);
  assign v_22273 = mux_22273(v_22274);
  assign v_22274 = ~v_7982;
  assign v_22275 = ~v_15134;
  assign v_22276 = v_22277 | v_22278;
  assign v_22277 = mux_22277(v_15136);
  assign v_22278 = mux_22278(v_22267);
  assign v_22279 = v_22280 & 1'h1;
  assign v_22280 = v_22281 & v_22282;
  assign v_22281 = ~act_7981;
  assign v_22282 = v_22283 | v_22287;
  assign v_22283 = v_22284 | v_22285;
  assign v_22284 = mux_22284(v_7975);
  assign v_22285 = mux_22285(v_22286);
  assign v_22286 = ~v_7975;
  assign v_22287 = ~v_7978;
  assign v_22288 = v_22289 | v_22290;
  assign v_22289 = mux_22289(v_7980);
  assign v_22290 = mux_22290(v_22279);
  assign v_22291 = v_22292 & 1'h1;
  assign v_22292 = v_22293 & v_22294;
  assign v_22293 = ~act_7974;
  assign v_22294 = v_22295 | v_22301;
  assign v_22295 = v_22296 | v_22299;
  assign v_22296 = mux_22296(v_22297);
  assign v_22297 = v_22298 & 1'h1;
  assign v_22298 = out_consume_en;
  assign v_22299 = mux_22299(v_22300);
  assign v_22300 = ~v_22297;
  assign v_22301 = ~v_7971;
  assign v_22302 = v_22303 | v_22304;
  assign v_22303 = mux_22303(v_7973);
  assign v_22304 = mux_22304(v_22291);
  assign v_22305 = mux_22305(v_22306);
  assign v_22306 = ~v_7967;
  assign v_22307 = ~v_7957;
  assign v_22308 = v_22309 | v_22310;
  assign v_22309 = mux_22309(v_7959);
  assign v_22310 = mux_22310(v_7961);
  assign v_22311 = mux_22311(v_22312);
  assign v_22312 = ~v_7953;
  assign v_22313 = ~v_4398;
  assign v_22314 = v_22315 | v_22316;
  assign v_22315 = mux_22315(v_4400);
  assign v_22316 = mux_22316(v_7947);
  assign v_22317 = mux_22317(v_22318);
  assign v_22318 = ~v_4395;
  assign v_22319 = ~v_4385;
  assign v_22320 = v_22321 | v_22322;
  assign v_22321 = mux_22321(v_4387);
  assign v_22322 = mux_22322(v_4389);
  assign v_22323 = mux_22323(v_22324);
  assign v_22324 = ~v_4381;
  assign v_22325 = ~v_2618;
  assign v_22326 = v_22327 | v_22328;
  assign v_22327 = mux_22327(v_2620);
  assign v_22328 = mux_22328(v_4375);
  assign v_22329 = mux_22329(v_22330);
  assign v_22330 = ~v_2615;
  assign v_22331 = ~v_2605;
  assign v_22332 = v_22333 | v_22334;
  assign v_22333 = mux_22333(v_2607);
  assign v_22334 = mux_22334(v_2609);
  assign v_22335 = mux_22335(v_22336);
  assign v_22336 = ~v_2601;
  assign v_22337 = ~v_1734;
  assign v_22338 = v_22339 | v_22340;
  assign v_22339 = mux_22339(v_1736);
  assign v_22340 = mux_22340(v_2595);
  assign v_22341 = mux_22341(v_22342);
  assign v_22342 = ~v_1731;
  assign v_22343 = ~v_845;
  assign v_22344 = v_22345 | v_22346;
  assign v_22345 = mux_22345(v_847);
  assign v_22346 = mux_22346(v_1725);
  assign v_22347 = mux_22347(v_22348);
  assign v_22348 = ~v_841;
  assign v_22349 = ~v_403;
  assign v_22350 = v_22351 | v_22352;
  assign v_22351 = mux_22351(v_405);
  assign v_22352 = mux_22352(v_835);
  assign v_22353 = mux_22353(v_22354);
  assign v_22354 = ~v_399;
  assign v_22355 = ~v_185;
  assign v_22356 = v_22357 | v_22358;
  assign v_22357 = mux_22357(v_187);
  assign v_22358 = mux_22358(v_393);
  assign v_22359 = mux_22359(v_22360);
  assign v_22360 = ~v_181;
  assign v_22361 = ~v_79;
  assign v_22362 = v_22363 | v_22364;
  assign v_22363 = mux_22363(v_81);
  assign v_22364 = mux_22364(v_175);
  assign v_22365 = mux_22365(v_22366);
  assign v_22366 = ~v_75;
  assign v_22367 = ~v_29;
  assign v_22368 = v_22369 | v_22370;
  assign v_22369 = mux_22369(v_31);
  assign v_22370 = mux_22370(v_69);
  assign v_22371 = mux_22371(v_22372);
  assign v_22372 = ~v_25;
  assign v_22373 = ~v_7;
  assign v_22374 = v_22375 | v_22376;
  assign v_22375 = mux_22375(v_9);
  assign v_22376 = mux_22376(v_19);
  assign v_22377 = mux_22377(v_22378);
  assign v_22378 = ~v_2;
  assign in0_consume_en = v_22380;
  assign v_22380 = mux_22380(v_22381);
  assign v_22381 = ~1'h0;
  assign out_canPeek = v_7971;
  assign out_peek = v_22384;
  assign v_22385 = v_22386 | v_22388;
  assign v_22386 = mux_22386(v_22387);
  assign v_22387 = ~act_7974;
  assign v_22388 = v_22389 | v_25967;
  assign v_22389 = mux_22389(v_7975);
  assign v_22391 = v_22392 | v_22394;
  assign v_22392 = mux_22392(v_22393);
  assign v_22393 = ~act_7981;
  assign v_22394 = v_22395 | v_24181;
  assign v_22395 = mux_22395(v_7982);
  assign v_22397 = v_22398 | v_22400;
  assign v_22398 = mux_22398(v_22399);
  assign v_22399 = ~act_15137;
  assign v_22400 = v_22401 | v_23291;
  assign v_22401 = mux_22401(v_15138);
  assign v_22403 = v_22404 | v_22406;
  assign v_22404 = mux_22404(v_22405);
  assign v_22405 = ~act_18709;
  assign v_22406 = v_22407 | v_22849;
  assign v_22407 = mux_22407(v_18710);
  assign v_22409 = v_22410 | v_22412;
  assign v_22410 = mux_22410(v_22411);
  assign v_22411 = ~act_20489;
  assign v_22412 = v_22413 | v_22631;
  assign v_22413 = mux_22413(v_20490);
  assign v_22415 = v_22416 | v_22418;
  assign v_22416 = mux_22416(v_22417);
  assign v_22417 = ~act_21373;
  assign v_22418 = v_22419 | v_22525;
  assign v_22419 = mux_22419(v_21374);
  assign v_22421 = v_22422 | v_22424;
  assign v_22422 = mux_22422(v_22423);
  assign v_22423 = ~act_21809;
  assign v_22424 = v_22425 | v_22475;
  assign v_22425 = mux_22425(v_21810);
  assign v_22427 = v_22428 | v_22430;
  assign v_22428 = mux_22428(v_22429);
  assign v_22429 = ~act_22021;
  assign v_22430 = v_22431 | v_22453;
  assign v_22431 = mux_22431(v_22022);
  assign v_22433 = v_22434 | v_22436;
  assign v_22434 = mux_22434(v_22435);
  assign v_22435 = ~act_22121;
  assign v_22436 = v_22437 | v_22445;
  assign v_22437 = mux_22437(v_22122);
  assign v_22439 = v_22440 | v_22442;
  assign v_22440 = mux_22440(v_22441);
  assign v_22441 = ~act_22165;
  assign v_22442 = v_22443 | v_22444;
  assign v_22443 = mux_22443(v_22166);
  assign v_22444 = mux_22444(v_22172);
  assign v_22445 = mux_22445(v_22152);
  assign v_22447 = v_22448 | v_22450;
  assign v_22448 = mux_22448(v_22449);
  assign v_22449 = ~act_22128;
  assign v_22450 = v_22451 | v_22452;
  assign v_22451 = mux_22451(v_22129);
  assign v_22452 = mux_22452(v_22135);
  assign v_22453 = mux_22453(v_22108);
  assign v_22455 = v_22456 | v_22458;
  assign v_22456 = mux_22456(v_22457);
  assign v_22457 = ~act_22028;
  assign v_22458 = v_22459 | v_22467;
  assign v_22459 = mux_22459(v_22029);
  assign v_22461 = v_22462 | v_22464;
  assign v_22462 = mux_22462(v_22463);
  assign v_22463 = ~act_22072;
  assign v_22464 = v_22465 | v_22466;
  assign v_22465 = mux_22465(v_22073);
  assign v_22466 = mux_22466(v_22079);
  assign v_22467 = mux_22467(v_22059);
  assign v_22469 = v_22470 | v_22472;
  assign v_22470 = mux_22470(v_22471);
  assign v_22471 = ~act_22035;
  assign v_22472 = v_22473 | v_22474;
  assign v_22473 = mux_22473(v_22036);
  assign v_22474 = mux_22474(v_22042);
  assign v_22475 = mux_22475(v_22008);
  assign v_22477 = v_22478 | v_22480;
  assign v_22478 = mux_22478(v_22479);
  assign v_22479 = ~act_21816;
  assign v_22480 = v_22481 | v_22503;
  assign v_22481 = mux_22481(v_21817);
  assign v_22483 = v_22484 | v_22486;
  assign v_22484 = mux_22484(v_22485);
  assign v_22485 = ~act_21916;
  assign v_22486 = v_22487 | v_22495;
  assign v_22487 = mux_22487(v_21917);
  assign v_22489 = v_22490 | v_22492;
  assign v_22490 = mux_22490(v_22491);
  assign v_22491 = ~act_21960;
  assign v_22492 = v_22493 | v_22494;
  assign v_22493 = mux_22493(v_21961);
  assign v_22494 = mux_22494(v_21967);
  assign v_22495 = mux_22495(v_21947);
  assign v_22497 = v_22498 | v_22500;
  assign v_22498 = mux_22498(v_22499);
  assign v_22499 = ~act_21923;
  assign v_22500 = v_22501 | v_22502;
  assign v_22501 = mux_22501(v_21924);
  assign v_22502 = mux_22502(v_21930);
  assign v_22503 = mux_22503(v_21903);
  assign v_22505 = v_22506 | v_22508;
  assign v_22506 = mux_22506(v_22507);
  assign v_22507 = ~act_21823;
  assign v_22508 = v_22509 | v_22517;
  assign v_22509 = mux_22509(v_21824);
  assign v_22511 = v_22512 | v_22514;
  assign v_22512 = mux_22512(v_22513);
  assign v_22513 = ~act_21867;
  assign v_22514 = v_22515 | v_22516;
  assign v_22515 = mux_22515(v_21868);
  assign v_22516 = mux_22516(v_21874);
  assign v_22517 = mux_22517(v_21854);
  assign v_22519 = v_22520 | v_22522;
  assign v_22520 = mux_22520(v_22521);
  assign v_22521 = ~act_21830;
  assign v_22522 = v_22523 | v_22524;
  assign v_22523 = mux_22523(v_21831);
  assign v_22524 = mux_22524(v_21837);
  assign v_22525 = mux_22525(v_21796);
  assign v_22527 = v_22528 | v_22530;
  assign v_22528 = mux_22528(v_22529);
  assign v_22529 = ~act_21380;
  assign v_22530 = v_22531 | v_22581;
  assign v_22531 = mux_22531(v_21381);
  assign v_22533 = v_22534 | v_22536;
  assign v_22534 = mux_22534(v_22535);
  assign v_22535 = ~act_21592;
  assign v_22536 = v_22537 | v_22559;
  assign v_22537 = mux_22537(v_21593);
  assign v_22539 = v_22540 | v_22542;
  assign v_22540 = mux_22540(v_22541);
  assign v_22541 = ~act_21692;
  assign v_22542 = v_22543 | v_22551;
  assign v_22543 = mux_22543(v_21693);
  assign v_22545 = v_22546 | v_22548;
  assign v_22546 = mux_22546(v_22547);
  assign v_22547 = ~act_21736;
  assign v_22548 = v_22549 | v_22550;
  assign v_22549 = mux_22549(v_21737);
  assign v_22550 = mux_22550(v_21743);
  assign v_22551 = mux_22551(v_21723);
  assign v_22553 = v_22554 | v_22556;
  assign v_22554 = mux_22554(v_22555);
  assign v_22555 = ~act_21699;
  assign v_22556 = v_22557 | v_22558;
  assign v_22557 = mux_22557(v_21700);
  assign v_22558 = mux_22558(v_21706);
  assign v_22559 = mux_22559(v_21679);
  assign v_22561 = v_22562 | v_22564;
  assign v_22562 = mux_22562(v_22563);
  assign v_22563 = ~act_21599;
  assign v_22564 = v_22565 | v_22573;
  assign v_22565 = mux_22565(v_21600);
  assign v_22567 = v_22568 | v_22570;
  assign v_22568 = mux_22568(v_22569);
  assign v_22569 = ~act_21643;
  assign v_22570 = v_22571 | v_22572;
  assign v_22571 = mux_22571(v_21644);
  assign v_22572 = mux_22572(v_21650);
  assign v_22573 = mux_22573(v_21630);
  assign v_22575 = v_22576 | v_22578;
  assign v_22576 = mux_22576(v_22577);
  assign v_22577 = ~act_21606;
  assign v_22578 = v_22579 | v_22580;
  assign v_22579 = mux_22579(v_21607);
  assign v_22580 = mux_22580(v_21613);
  assign v_22581 = mux_22581(v_21579);
  assign v_22583 = v_22584 | v_22586;
  assign v_22584 = mux_22584(v_22585);
  assign v_22585 = ~act_21387;
  assign v_22586 = v_22587 | v_22609;
  assign v_22587 = mux_22587(v_21388);
  assign v_22589 = v_22590 | v_22592;
  assign v_22590 = mux_22590(v_22591);
  assign v_22591 = ~act_21487;
  assign v_22592 = v_22593 | v_22601;
  assign v_22593 = mux_22593(v_21488);
  assign v_22595 = v_22596 | v_22598;
  assign v_22596 = mux_22596(v_22597);
  assign v_22597 = ~act_21531;
  assign v_22598 = v_22599 | v_22600;
  assign v_22599 = mux_22599(v_21532);
  assign v_22600 = mux_22600(v_21538);
  assign v_22601 = mux_22601(v_21518);
  assign v_22603 = v_22604 | v_22606;
  assign v_22604 = mux_22604(v_22605);
  assign v_22605 = ~act_21494;
  assign v_22606 = v_22607 | v_22608;
  assign v_22607 = mux_22607(v_21495);
  assign v_22608 = mux_22608(v_21501);
  assign v_22609 = mux_22609(v_21474);
  assign v_22611 = v_22612 | v_22614;
  assign v_22612 = mux_22612(v_22613);
  assign v_22613 = ~act_21394;
  assign v_22614 = v_22615 | v_22623;
  assign v_22615 = mux_22615(v_21395);
  assign v_22617 = v_22618 | v_22620;
  assign v_22618 = mux_22618(v_22619);
  assign v_22619 = ~act_21438;
  assign v_22620 = v_22621 | v_22622;
  assign v_22621 = mux_22621(v_21439);
  assign v_22622 = mux_22622(v_21445);
  assign v_22623 = mux_22623(v_21425);
  assign v_22625 = v_22626 | v_22628;
  assign v_22626 = mux_22626(v_22627);
  assign v_22627 = ~act_21401;
  assign v_22628 = v_22629 | v_22630;
  assign v_22629 = mux_22629(v_21402);
  assign v_22630 = mux_22630(v_21408);
  assign v_22631 = mux_22631(v_21360);
  assign v_22633 = v_22634 | v_22636;
  assign v_22634 = mux_22634(v_22635);
  assign v_22635 = ~act_20496;
  assign v_22636 = v_22637 | v_22743;
  assign v_22637 = mux_22637(v_20497);
  assign v_22639 = v_22640 | v_22642;
  assign v_22640 = mux_22640(v_22641);
  assign v_22641 = ~act_20932;
  assign v_22642 = v_22643 | v_22693;
  assign v_22643 = mux_22643(v_20933);
  assign v_22645 = v_22646 | v_22648;
  assign v_22646 = mux_22646(v_22647);
  assign v_22647 = ~act_21144;
  assign v_22648 = v_22649 | v_22671;
  assign v_22649 = mux_22649(v_21145);
  assign v_22651 = v_22652 | v_22654;
  assign v_22652 = mux_22652(v_22653);
  assign v_22653 = ~act_21244;
  assign v_22654 = v_22655 | v_22663;
  assign v_22655 = mux_22655(v_21245);
  assign v_22657 = v_22658 | v_22660;
  assign v_22658 = mux_22658(v_22659);
  assign v_22659 = ~act_21288;
  assign v_22660 = v_22661 | v_22662;
  assign v_22661 = mux_22661(v_21289);
  assign v_22662 = mux_22662(v_21295);
  assign v_22663 = mux_22663(v_21275);
  assign v_22665 = v_22666 | v_22668;
  assign v_22666 = mux_22666(v_22667);
  assign v_22667 = ~act_21251;
  assign v_22668 = v_22669 | v_22670;
  assign v_22669 = mux_22669(v_21252);
  assign v_22670 = mux_22670(v_21258);
  assign v_22671 = mux_22671(v_21231);
  assign v_22673 = v_22674 | v_22676;
  assign v_22674 = mux_22674(v_22675);
  assign v_22675 = ~act_21151;
  assign v_22676 = v_22677 | v_22685;
  assign v_22677 = mux_22677(v_21152);
  assign v_22679 = v_22680 | v_22682;
  assign v_22680 = mux_22680(v_22681);
  assign v_22681 = ~act_21195;
  assign v_22682 = v_22683 | v_22684;
  assign v_22683 = mux_22683(v_21196);
  assign v_22684 = mux_22684(v_21202);
  assign v_22685 = mux_22685(v_21182);
  assign v_22687 = v_22688 | v_22690;
  assign v_22688 = mux_22688(v_22689);
  assign v_22689 = ~act_21158;
  assign v_22690 = v_22691 | v_22692;
  assign v_22691 = mux_22691(v_21159);
  assign v_22692 = mux_22692(v_21165);
  assign v_22693 = mux_22693(v_21131);
  assign v_22695 = v_22696 | v_22698;
  assign v_22696 = mux_22696(v_22697);
  assign v_22697 = ~act_20939;
  assign v_22698 = v_22699 | v_22721;
  assign v_22699 = mux_22699(v_20940);
  assign v_22701 = v_22702 | v_22704;
  assign v_22702 = mux_22702(v_22703);
  assign v_22703 = ~act_21039;
  assign v_22704 = v_22705 | v_22713;
  assign v_22705 = mux_22705(v_21040);
  assign v_22707 = v_22708 | v_22710;
  assign v_22708 = mux_22708(v_22709);
  assign v_22709 = ~act_21083;
  assign v_22710 = v_22711 | v_22712;
  assign v_22711 = mux_22711(v_21084);
  assign v_22712 = mux_22712(v_21090);
  assign v_22713 = mux_22713(v_21070);
  assign v_22715 = v_22716 | v_22718;
  assign v_22716 = mux_22716(v_22717);
  assign v_22717 = ~act_21046;
  assign v_22718 = v_22719 | v_22720;
  assign v_22719 = mux_22719(v_21047);
  assign v_22720 = mux_22720(v_21053);
  assign v_22721 = mux_22721(v_21026);
  assign v_22723 = v_22724 | v_22726;
  assign v_22724 = mux_22724(v_22725);
  assign v_22725 = ~act_20946;
  assign v_22726 = v_22727 | v_22735;
  assign v_22727 = mux_22727(v_20947);
  assign v_22729 = v_22730 | v_22732;
  assign v_22730 = mux_22730(v_22731);
  assign v_22731 = ~act_20990;
  assign v_22732 = v_22733 | v_22734;
  assign v_22733 = mux_22733(v_20991);
  assign v_22734 = mux_22734(v_20997);
  assign v_22735 = mux_22735(v_20977);
  assign v_22737 = v_22738 | v_22740;
  assign v_22738 = mux_22738(v_22739);
  assign v_22739 = ~act_20953;
  assign v_22740 = v_22741 | v_22742;
  assign v_22741 = mux_22741(v_20954);
  assign v_22742 = mux_22742(v_20960);
  assign v_22743 = mux_22743(v_20919);
  assign v_22745 = v_22746 | v_22748;
  assign v_22746 = mux_22746(v_22747);
  assign v_22747 = ~act_20503;
  assign v_22748 = v_22749 | v_22799;
  assign v_22749 = mux_22749(v_20504);
  assign v_22751 = v_22752 | v_22754;
  assign v_22752 = mux_22752(v_22753);
  assign v_22753 = ~act_20715;
  assign v_22754 = v_22755 | v_22777;
  assign v_22755 = mux_22755(v_20716);
  assign v_22757 = v_22758 | v_22760;
  assign v_22758 = mux_22758(v_22759);
  assign v_22759 = ~act_20815;
  assign v_22760 = v_22761 | v_22769;
  assign v_22761 = mux_22761(v_20816);
  assign v_22763 = v_22764 | v_22766;
  assign v_22764 = mux_22764(v_22765);
  assign v_22765 = ~act_20859;
  assign v_22766 = v_22767 | v_22768;
  assign v_22767 = mux_22767(v_20860);
  assign v_22768 = mux_22768(v_20866);
  assign v_22769 = mux_22769(v_20846);
  assign v_22771 = v_22772 | v_22774;
  assign v_22772 = mux_22772(v_22773);
  assign v_22773 = ~act_20822;
  assign v_22774 = v_22775 | v_22776;
  assign v_22775 = mux_22775(v_20823);
  assign v_22776 = mux_22776(v_20829);
  assign v_22777 = mux_22777(v_20802);
  assign v_22779 = v_22780 | v_22782;
  assign v_22780 = mux_22780(v_22781);
  assign v_22781 = ~act_20722;
  assign v_22782 = v_22783 | v_22791;
  assign v_22783 = mux_22783(v_20723);
  assign v_22785 = v_22786 | v_22788;
  assign v_22786 = mux_22786(v_22787);
  assign v_22787 = ~act_20766;
  assign v_22788 = v_22789 | v_22790;
  assign v_22789 = mux_22789(v_20767);
  assign v_22790 = mux_22790(v_20773);
  assign v_22791 = mux_22791(v_20753);
  assign v_22793 = v_22794 | v_22796;
  assign v_22794 = mux_22794(v_22795);
  assign v_22795 = ~act_20729;
  assign v_22796 = v_22797 | v_22798;
  assign v_22797 = mux_22797(v_20730);
  assign v_22798 = mux_22798(v_20736);
  assign v_22799 = mux_22799(v_20702);
  assign v_22801 = v_22802 | v_22804;
  assign v_22802 = mux_22802(v_22803);
  assign v_22803 = ~act_20510;
  assign v_22804 = v_22805 | v_22827;
  assign v_22805 = mux_22805(v_20511);
  assign v_22807 = v_22808 | v_22810;
  assign v_22808 = mux_22808(v_22809);
  assign v_22809 = ~act_20610;
  assign v_22810 = v_22811 | v_22819;
  assign v_22811 = mux_22811(v_20611);
  assign v_22813 = v_22814 | v_22816;
  assign v_22814 = mux_22814(v_22815);
  assign v_22815 = ~act_20654;
  assign v_22816 = v_22817 | v_22818;
  assign v_22817 = mux_22817(v_20655);
  assign v_22818 = mux_22818(v_20661);
  assign v_22819 = mux_22819(v_20641);
  assign v_22821 = v_22822 | v_22824;
  assign v_22822 = mux_22822(v_22823);
  assign v_22823 = ~act_20617;
  assign v_22824 = v_22825 | v_22826;
  assign v_22825 = mux_22825(v_20618);
  assign v_22826 = mux_22826(v_20624);
  assign v_22827 = mux_22827(v_20597);
  assign v_22829 = v_22830 | v_22832;
  assign v_22830 = mux_22830(v_22831);
  assign v_22831 = ~act_20517;
  assign v_22832 = v_22833 | v_22841;
  assign v_22833 = mux_22833(v_20518);
  assign v_22835 = v_22836 | v_22838;
  assign v_22836 = mux_22836(v_22837);
  assign v_22837 = ~act_20561;
  assign v_22838 = v_22839 | v_22840;
  assign v_22839 = mux_22839(v_20562);
  assign v_22840 = mux_22840(v_20568);
  assign v_22841 = mux_22841(v_20548);
  assign v_22843 = v_22844 | v_22846;
  assign v_22844 = mux_22844(v_22845);
  assign v_22845 = ~act_20524;
  assign v_22846 = v_22847 | v_22848;
  assign v_22847 = mux_22847(v_20525);
  assign v_22848 = mux_22848(v_20531);
  assign v_22849 = mux_22849(v_20476);
  assign v_22851 = v_22852 | v_22854;
  assign v_22852 = mux_22852(v_22853);
  assign v_22853 = ~act_18716;
  assign v_22854 = v_22855 | v_23073;
  assign v_22855 = mux_22855(v_18717);
  assign v_22857 = v_22858 | v_22860;
  assign v_22858 = mux_22858(v_22859);
  assign v_22859 = ~act_19600;
  assign v_22860 = v_22861 | v_22967;
  assign v_22861 = mux_22861(v_19601);
  assign v_22863 = v_22864 | v_22866;
  assign v_22864 = mux_22864(v_22865);
  assign v_22865 = ~act_20036;
  assign v_22866 = v_22867 | v_22917;
  assign v_22867 = mux_22867(v_20037);
  assign v_22869 = v_22870 | v_22872;
  assign v_22870 = mux_22870(v_22871);
  assign v_22871 = ~act_20248;
  assign v_22872 = v_22873 | v_22895;
  assign v_22873 = mux_22873(v_20249);
  assign v_22875 = v_22876 | v_22878;
  assign v_22876 = mux_22876(v_22877);
  assign v_22877 = ~act_20348;
  assign v_22878 = v_22879 | v_22887;
  assign v_22879 = mux_22879(v_20349);
  assign v_22881 = v_22882 | v_22884;
  assign v_22882 = mux_22882(v_22883);
  assign v_22883 = ~act_20392;
  assign v_22884 = v_22885 | v_22886;
  assign v_22885 = mux_22885(v_20393);
  assign v_22886 = mux_22886(v_20399);
  assign v_22887 = mux_22887(v_20379);
  assign v_22889 = v_22890 | v_22892;
  assign v_22890 = mux_22890(v_22891);
  assign v_22891 = ~act_20355;
  assign v_22892 = v_22893 | v_22894;
  assign v_22893 = mux_22893(v_20356);
  assign v_22894 = mux_22894(v_20362);
  assign v_22895 = mux_22895(v_20335);
  assign v_22897 = v_22898 | v_22900;
  assign v_22898 = mux_22898(v_22899);
  assign v_22899 = ~act_20255;
  assign v_22900 = v_22901 | v_22909;
  assign v_22901 = mux_22901(v_20256);
  assign v_22903 = v_22904 | v_22906;
  assign v_22904 = mux_22904(v_22905);
  assign v_22905 = ~act_20299;
  assign v_22906 = v_22907 | v_22908;
  assign v_22907 = mux_22907(v_20300);
  assign v_22908 = mux_22908(v_20306);
  assign v_22909 = mux_22909(v_20286);
  assign v_22911 = v_22912 | v_22914;
  assign v_22912 = mux_22912(v_22913);
  assign v_22913 = ~act_20262;
  assign v_22914 = v_22915 | v_22916;
  assign v_22915 = mux_22915(v_20263);
  assign v_22916 = mux_22916(v_20269);
  assign v_22917 = mux_22917(v_20235);
  assign v_22919 = v_22920 | v_22922;
  assign v_22920 = mux_22920(v_22921);
  assign v_22921 = ~act_20043;
  assign v_22922 = v_22923 | v_22945;
  assign v_22923 = mux_22923(v_20044);
  assign v_22925 = v_22926 | v_22928;
  assign v_22926 = mux_22926(v_22927);
  assign v_22927 = ~act_20143;
  assign v_22928 = v_22929 | v_22937;
  assign v_22929 = mux_22929(v_20144);
  assign v_22931 = v_22932 | v_22934;
  assign v_22932 = mux_22932(v_22933);
  assign v_22933 = ~act_20187;
  assign v_22934 = v_22935 | v_22936;
  assign v_22935 = mux_22935(v_20188);
  assign v_22936 = mux_22936(v_20194);
  assign v_22937 = mux_22937(v_20174);
  assign v_22939 = v_22940 | v_22942;
  assign v_22940 = mux_22940(v_22941);
  assign v_22941 = ~act_20150;
  assign v_22942 = v_22943 | v_22944;
  assign v_22943 = mux_22943(v_20151);
  assign v_22944 = mux_22944(v_20157);
  assign v_22945 = mux_22945(v_20130);
  assign v_22947 = v_22948 | v_22950;
  assign v_22948 = mux_22948(v_22949);
  assign v_22949 = ~act_20050;
  assign v_22950 = v_22951 | v_22959;
  assign v_22951 = mux_22951(v_20051);
  assign v_22953 = v_22954 | v_22956;
  assign v_22954 = mux_22954(v_22955);
  assign v_22955 = ~act_20094;
  assign v_22956 = v_22957 | v_22958;
  assign v_22957 = mux_22957(v_20095);
  assign v_22958 = mux_22958(v_20101);
  assign v_22959 = mux_22959(v_20081);
  assign v_22961 = v_22962 | v_22964;
  assign v_22962 = mux_22962(v_22963);
  assign v_22963 = ~act_20057;
  assign v_22964 = v_22965 | v_22966;
  assign v_22965 = mux_22965(v_20058);
  assign v_22966 = mux_22966(v_20064);
  assign v_22967 = mux_22967(v_20023);
  assign v_22969 = v_22970 | v_22972;
  assign v_22970 = mux_22970(v_22971);
  assign v_22971 = ~act_19607;
  assign v_22972 = v_22973 | v_23023;
  assign v_22973 = mux_22973(v_19608);
  assign v_22975 = v_22976 | v_22978;
  assign v_22976 = mux_22976(v_22977);
  assign v_22977 = ~act_19819;
  assign v_22978 = v_22979 | v_23001;
  assign v_22979 = mux_22979(v_19820);
  assign v_22981 = v_22982 | v_22984;
  assign v_22982 = mux_22982(v_22983);
  assign v_22983 = ~act_19919;
  assign v_22984 = v_22985 | v_22993;
  assign v_22985 = mux_22985(v_19920);
  assign v_22987 = v_22988 | v_22990;
  assign v_22988 = mux_22988(v_22989);
  assign v_22989 = ~act_19963;
  assign v_22990 = v_22991 | v_22992;
  assign v_22991 = mux_22991(v_19964);
  assign v_22992 = mux_22992(v_19970);
  assign v_22993 = mux_22993(v_19950);
  assign v_22995 = v_22996 | v_22998;
  assign v_22996 = mux_22996(v_22997);
  assign v_22997 = ~act_19926;
  assign v_22998 = v_22999 | v_23000;
  assign v_22999 = mux_22999(v_19927);
  assign v_23000 = mux_23000(v_19933);
  assign v_23001 = mux_23001(v_19906);
  assign v_23003 = v_23004 | v_23006;
  assign v_23004 = mux_23004(v_23005);
  assign v_23005 = ~act_19826;
  assign v_23006 = v_23007 | v_23015;
  assign v_23007 = mux_23007(v_19827);
  assign v_23009 = v_23010 | v_23012;
  assign v_23010 = mux_23010(v_23011);
  assign v_23011 = ~act_19870;
  assign v_23012 = v_23013 | v_23014;
  assign v_23013 = mux_23013(v_19871);
  assign v_23014 = mux_23014(v_19877);
  assign v_23015 = mux_23015(v_19857);
  assign v_23017 = v_23018 | v_23020;
  assign v_23018 = mux_23018(v_23019);
  assign v_23019 = ~act_19833;
  assign v_23020 = v_23021 | v_23022;
  assign v_23021 = mux_23021(v_19834);
  assign v_23022 = mux_23022(v_19840);
  assign v_23023 = mux_23023(v_19806);
  assign v_23025 = v_23026 | v_23028;
  assign v_23026 = mux_23026(v_23027);
  assign v_23027 = ~act_19614;
  assign v_23028 = v_23029 | v_23051;
  assign v_23029 = mux_23029(v_19615);
  assign v_23031 = v_23032 | v_23034;
  assign v_23032 = mux_23032(v_23033);
  assign v_23033 = ~act_19714;
  assign v_23034 = v_23035 | v_23043;
  assign v_23035 = mux_23035(v_19715);
  assign v_23037 = v_23038 | v_23040;
  assign v_23038 = mux_23038(v_23039);
  assign v_23039 = ~act_19758;
  assign v_23040 = v_23041 | v_23042;
  assign v_23041 = mux_23041(v_19759);
  assign v_23042 = mux_23042(v_19765);
  assign v_23043 = mux_23043(v_19745);
  assign v_23045 = v_23046 | v_23048;
  assign v_23046 = mux_23046(v_23047);
  assign v_23047 = ~act_19721;
  assign v_23048 = v_23049 | v_23050;
  assign v_23049 = mux_23049(v_19722);
  assign v_23050 = mux_23050(v_19728);
  assign v_23051 = mux_23051(v_19701);
  assign v_23053 = v_23054 | v_23056;
  assign v_23054 = mux_23054(v_23055);
  assign v_23055 = ~act_19621;
  assign v_23056 = v_23057 | v_23065;
  assign v_23057 = mux_23057(v_19622);
  assign v_23059 = v_23060 | v_23062;
  assign v_23060 = mux_23060(v_23061);
  assign v_23061 = ~act_19665;
  assign v_23062 = v_23063 | v_23064;
  assign v_23063 = mux_23063(v_19666);
  assign v_23064 = mux_23064(v_19672);
  assign v_23065 = mux_23065(v_19652);
  assign v_23067 = v_23068 | v_23070;
  assign v_23068 = mux_23068(v_23069);
  assign v_23069 = ~act_19628;
  assign v_23070 = v_23071 | v_23072;
  assign v_23071 = mux_23071(v_19629);
  assign v_23072 = mux_23072(v_19635);
  assign v_23073 = mux_23073(v_19587);
  assign v_23075 = v_23076 | v_23078;
  assign v_23076 = mux_23076(v_23077);
  assign v_23077 = ~act_18723;
  assign v_23078 = v_23079 | v_23185;
  assign v_23079 = mux_23079(v_18724);
  assign v_23081 = v_23082 | v_23084;
  assign v_23082 = mux_23082(v_23083);
  assign v_23083 = ~act_19159;
  assign v_23084 = v_23085 | v_23135;
  assign v_23085 = mux_23085(v_19160);
  assign v_23087 = v_23088 | v_23090;
  assign v_23088 = mux_23088(v_23089);
  assign v_23089 = ~act_19371;
  assign v_23090 = v_23091 | v_23113;
  assign v_23091 = mux_23091(v_19372);
  assign v_23093 = v_23094 | v_23096;
  assign v_23094 = mux_23094(v_23095);
  assign v_23095 = ~act_19471;
  assign v_23096 = v_23097 | v_23105;
  assign v_23097 = mux_23097(v_19472);
  assign v_23099 = v_23100 | v_23102;
  assign v_23100 = mux_23100(v_23101);
  assign v_23101 = ~act_19515;
  assign v_23102 = v_23103 | v_23104;
  assign v_23103 = mux_23103(v_19516);
  assign v_23104 = mux_23104(v_19522);
  assign v_23105 = mux_23105(v_19502);
  assign v_23107 = v_23108 | v_23110;
  assign v_23108 = mux_23108(v_23109);
  assign v_23109 = ~act_19478;
  assign v_23110 = v_23111 | v_23112;
  assign v_23111 = mux_23111(v_19479);
  assign v_23112 = mux_23112(v_19485);
  assign v_23113 = mux_23113(v_19458);
  assign v_23115 = v_23116 | v_23118;
  assign v_23116 = mux_23116(v_23117);
  assign v_23117 = ~act_19378;
  assign v_23118 = v_23119 | v_23127;
  assign v_23119 = mux_23119(v_19379);
  assign v_23121 = v_23122 | v_23124;
  assign v_23122 = mux_23122(v_23123);
  assign v_23123 = ~act_19422;
  assign v_23124 = v_23125 | v_23126;
  assign v_23125 = mux_23125(v_19423);
  assign v_23126 = mux_23126(v_19429);
  assign v_23127 = mux_23127(v_19409);
  assign v_23129 = v_23130 | v_23132;
  assign v_23130 = mux_23130(v_23131);
  assign v_23131 = ~act_19385;
  assign v_23132 = v_23133 | v_23134;
  assign v_23133 = mux_23133(v_19386);
  assign v_23134 = mux_23134(v_19392);
  assign v_23135 = mux_23135(v_19358);
  assign v_23137 = v_23138 | v_23140;
  assign v_23138 = mux_23138(v_23139);
  assign v_23139 = ~act_19166;
  assign v_23140 = v_23141 | v_23163;
  assign v_23141 = mux_23141(v_19167);
  assign v_23143 = v_23144 | v_23146;
  assign v_23144 = mux_23144(v_23145);
  assign v_23145 = ~act_19266;
  assign v_23146 = v_23147 | v_23155;
  assign v_23147 = mux_23147(v_19267);
  assign v_23149 = v_23150 | v_23152;
  assign v_23150 = mux_23150(v_23151);
  assign v_23151 = ~act_19310;
  assign v_23152 = v_23153 | v_23154;
  assign v_23153 = mux_23153(v_19311);
  assign v_23154 = mux_23154(v_19317);
  assign v_23155 = mux_23155(v_19297);
  assign v_23157 = v_23158 | v_23160;
  assign v_23158 = mux_23158(v_23159);
  assign v_23159 = ~act_19273;
  assign v_23160 = v_23161 | v_23162;
  assign v_23161 = mux_23161(v_19274);
  assign v_23162 = mux_23162(v_19280);
  assign v_23163 = mux_23163(v_19253);
  assign v_23165 = v_23166 | v_23168;
  assign v_23166 = mux_23166(v_23167);
  assign v_23167 = ~act_19173;
  assign v_23168 = v_23169 | v_23177;
  assign v_23169 = mux_23169(v_19174);
  assign v_23171 = v_23172 | v_23174;
  assign v_23172 = mux_23172(v_23173);
  assign v_23173 = ~act_19217;
  assign v_23174 = v_23175 | v_23176;
  assign v_23175 = mux_23175(v_19218);
  assign v_23176 = mux_23176(v_19224);
  assign v_23177 = mux_23177(v_19204);
  assign v_23179 = v_23180 | v_23182;
  assign v_23180 = mux_23180(v_23181);
  assign v_23181 = ~act_19180;
  assign v_23182 = v_23183 | v_23184;
  assign v_23183 = mux_23183(v_19181);
  assign v_23184 = mux_23184(v_19187);
  assign v_23185 = mux_23185(v_19146);
  assign v_23187 = v_23188 | v_23190;
  assign v_23188 = mux_23188(v_23189);
  assign v_23189 = ~act_18730;
  assign v_23190 = v_23191 | v_23241;
  assign v_23191 = mux_23191(v_18731);
  assign v_23193 = v_23194 | v_23196;
  assign v_23194 = mux_23194(v_23195);
  assign v_23195 = ~act_18942;
  assign v_23196 = v_23197 | v_23219;
  assign v_23197 = mux_23197(v_18943);
  assign v_23199 = v_23200 | v_23202;
  assign v_23200 = mux_23200(v_23201);
  assign v_23201 = ~act_19042;
  assign v_23202 = v_23203 | v_23211;
  assign v_23203 = mux_23203(v_19043);
  assign v_23205 = v_23206 | v_23208;
  assign v_23206 = mux_23206(v_23207);
  assign v_23207 = ~act_19086;
  assign v_23208 = v_23209 | v_23210;
  assign v_23209 = mux_23209(v_19087);
  assign v_23210 = mux_23210(v_19093);
  assign v_23211 = mux_23211(v_19073);
  assign v_23213 = v_23214 | v_23216;
  assign v_23214 = mux_23214(v_23215);
  assign v_23215 = ~act_19049;
  assign v_23216 = v_23217 | v_23218;
  assign v_23217 = mux_23217(v_19050);
  assign v_23218 = mux_23218(v_19056);
  assign v_23219 = mux_23219(v_19029);
  assign v_23221 = v_23222 | v_23224;
  assign v_23222 = mux_23222(v_23223);
  assign v_23223 = ~act_18949;
  assign v_23224 = v_23225 | v_23233;
  assign v_23225 = mux_23225(v_18950);
  assign v_23227 = v_23228 | v_23230;
  assign v_23228 = mux_23228(v_23229);
  assign v_23229 = ~act_18993;
  assign v_23230 = v_23231 | v_23232;
  assign v_23231 = mux_23231(v_18994);
  assign v_23232 = mux_23232(v_19000);
  assign v_23233 = mux_23233(v_18980);
  assign v_23235 = v_23236 | v_23238;
  assign v_23236 = mux_23236(v_23237);
  assign v_23237 = ~act_18956;
  assign v_23238 = v_23239 | v_23240;
  assign v_23239 = mux_23239(v_18957);
  assign v_23240 = mux_23240(v_18963);
  assign v_23241 = mux_23241(v_18929);
  assign v_23243 = v_23244 | v_23246;
  assign v_23244 = mux_23244(v_23245);
  assign v_23245 = ~act_18737;
  assign v_23246 = v_23247 | v_23269;
  assign v_23247 = mux_23247(v_18738);
  assign v_23249 = v_23250 | v_23252;
  assign v_23250 = mux_23250(v_23251);
  assign v_23251 = ~act_18837;
  assign v_23252 = v_23253 | v_23261;
  assign v_23253 = mux_23253(v_18838);
  assign v_23255 = v_23256 | v_23258;
  assign v_23256 = mux_23256(v_23257);
  assign v_23257 = ~act_18881;
  assign v_23258 = v_23259 | v_23260;
  assign v_23259 = mux_23259(v_18882);
  assign v_23260 = mux_23260(v_18888);
  assign v_23261 = mux_23261(v_18868);
  assign v_23263 = v_23264 | v_23266;
  assign v_23264 = mux_23264(v_23265);
  assign v_23265 = ~act_18844;
  assign v_23266 = v_23267 | v_23268;
  assign v_23267 = mux_23267(v_18845);
  assign v_23268 = mux_23268(v_18851);
  assign v_23269 = mux_23269(v_18824);
  assign v_23271 = v_23272 | v_23274;
  assign v_23272 = mux_23272(v_23273);
  assign v_23273 = ~act_18744;
  assign v_23274 = v_23275 | v_23283;
  assign v_23275 = mux_23275(v_18745);
  assign v_23277 = v_23278 | v_23280;
  assign v_23278 = mux_23278(v_23279);
  assign v_23279 = ~act_18788;
  assign v_23280 = v_23281 | v_23282;
  assign v_23281 = mux_23281(v_18789);
  assign v_23282 = mux_23282(v_18795);
  assign v_23283 = mux_23283(v_18775);
  assign v_23285 = v_23286 | v_23288;
  assign v_23286 = mux_23286(v_23287);
  assign v_23287 = ~act_18751;
  assign v_23288 = v_23289 | v_23290;
  assign v_23289 = mux_23289(v_18752);
  assign v_23290 = mux_23290(v_18758);
  assign v_23291 = mux_23291(v_18696);
  assign v_23293 = v_23294 | v_23296;
  assign v_23294 = mux_23294(v_23295);
  assign v_23295 = ~act_15144;
  assign v_23296 = v_23297 | v_23739;
  assign v_23297 = mux_23297(v_15145);
  assign v_23299 = v_23300 | v_23302;
  assign v_23300 = mux_23300(v_23301);
  assign v_23301 = ~act_16924;
  assign v_23302 = v_23303 | v_23521;
  assign v_23303 = mux_23303(v_16925);
  assign v_23305 = v_23306 | v_23308;
  assign v_23306 = mux_23306(v_23307);
  assign v_23307 = ~act_17808;
  assign v_23308 = v_23309 | v_23415;
  assign v_23309 = mux_23309(v_17809);
  assign v_23311 = v_23312 | v_23314;
  assign v_23312 = mux_23312(v_23313);
  assign v_23313 = ~act_18244;
  assign v_23314 = v_23315 | v_23365;
  assign v_23315 = mux_23315(v_18245);
  assign v_23317 = v_23318 | v_23320;
  assign v_23318 = mux_23318(v_23319);
  assign v_23319 = ~act_18456;
  assign v_23320 = v_23321 | v_23343;
  assign v_23321 = mux_23321(v_18457);
  assign v_23323 = v_23324 | v_23326;
  assign v_23324 = mux_23324(v_23325);
  assign v_23325 = ~act_18556;
  assign v_23326 = v_23327 | v_23335;
  assign v_23327 = mux_23327(v_18557);
  assign v_23329 = v_23330 | v_23332;
  assign v_23330 = mux_23330(v_23331);
  assign v_23331 = ~act_18600;
  assign v_23332 = v_23333 | v_23334;
  assign v_23333 = mux_23333(v_18601);
  assign v_23334 = mux_23334(v_18607);
  assign v_23335 = mux_23335(v_18587);
  assign v_23337 = v_23338 | v_23340;
  assign v_23338 = mux_23338(v_23339);
  assign v_23339 = ~act_18563;
  assign v_23340 = v_23341 | v_23342;
  assign v_23341 = mux_23341(v_18564);
  assign v_23342 = mux_23342(v_18570);
  assign v_23343 = mux_23343(v_18543);
  assign v_23345 = v_23346 | v_23348;
  assign v_23346 = mux_23346(v_23347);
  assign v_23347 = ~act_18463;
  assign v_23348 = v_23349 | v_23357;
  assign v_23349 = mux_23349(v_18464);
  assign v_23351 = v_23352 | v_23354;
  assign v_23352 = mux_23352(v_23353);
  assign v_23353 = ~act_18507;
  assign v_23354 = v_23355 | v_23356;
  assign v_23355 = mux_23355(v_18508);
  assign v_23356 = mux_23356(v_18514);
  assign v_23357 = mux_23357(v_18494);
  assign v_23359 = v_23360 | v_23362;
  assign v_23360 = mux_23360(v_23361);
  assign v_23361 = ~act_18470;
  assign v_23362 = v_23363 | v_23364;
  assign v_23363 = mux_23363(v_18471);
  assign v_23364 = mux_23364(v_18477);
  assign v_23365 = mux_23365(v_18443);
  assign v_23367 = v_23368 | v_23370;
  assign v_23368 = mux_23368(v_23369);
  assign v_23369 = ~act_18251;
  assign v_23370 = v_23371 | v_23393;
  assign v_23371 = mux_23371(v_18252);
  assign v_23373 = v_23374 | v_23376;
  assign v_23374 = mux_23374(v_23375);
  assign v_23375 = ~act_18351;
  assign v_23376 = v_23377 | v_23385;
  assign v_23377 = mux_23377(v_18352);
  assign v_23379 = v_23380 | v_23382;
  assign v_23380 = mux_23380(v_23381);
  assign v_23381 = ~act_18395;
  assign v_23382 = v_23383 | v_23384;
  assign v_23383 = mux_23383(v_18396);
  assign v_23384 = mux_23384(v_18402);
  assign v_23385 = mux_23385(v_18382);
  assign v_23387 = v_23388 | v_23390;
  assign v_23388 = mux_23388(v_23389);
  assign v_23389 = ~act_18358;
  assign v_23390 = v_23391 | v_23392;
  assign v_23391 = mux_23391(v_18359);
  assign v_23392 = mux_23392(v_18365);
  assign v_23393 = mux_23393(v_18338);
  assign v_23395 = v_23396 | v_23398;
  assign v_23396 = mux_23396(v_23397);
  assign v_23397 = ~act_18258;
  assign v_23398 = v_23399 | v_23407;
  assign v_23399 = mux_23399(v_18259);
  assign v_23401 = v_23402 | v_23404;
  assign v_23402 = mux_23402(v_23403);
  assign v_23403 = ~act_18302;
  assign v_23404 = v_23405 | v_23406;
  assign v_23405 = mux_23405(v_18303);
  assign v_23406 = mux_23406(v_18309);
  assign v_23407 = mux_23407(v_18289);
  assign v_23409 = v_23410 | v_23412;
  assign v_23410 = mux_23410(v_23411);
  assign v_23411 = ~act_18265;
  assign v_23412 = v_23413 | v_23414;
  assign v_23413 = mux_23413(v_18266);
  assign v_23414 = mux_23414(v_18272);
  assign v_23415 = mux_23415(v_18231);
  assign v_23417 = v_23418 | v_23420;
  assign v_23418 = mux_23418(v_23419);
  assign v_23419 = ~act_17815;
  assign v_23420 = v_23421 | v_23471;
  assign v_23421 = mux_23421(v_17816);
  assign v_23423 = v_23424 | v_23426;
  assign v_23424 = mux_23424(v_23425);
  assign v_23425 = ~act_18027;
  assign v_23426 = v_23427 | v_23449;
  assign v_23427 = mux_23427(v_18028);
  assign v_23429 = v_23430 | v_23432;
  assign v_23430 = mux_23430(v_23431);
  assign v_23431 = ~act_18127;
  assign v_23432 = v_23433 | v_23441;
  assign v_23433 = mux_23433(v_18128);
  assign v_23435 = v_23436 | v_23438;
  assign v_23436 = mux_23436(v_23437);
  assign v_23437 = ~act_18171;
  assign v_23438 = v_23439 | v_23440;
  assign v_23439 = mux_23439(v_18172);
  assign v_23440 = mux_23440(v_18178);
  assign v_23441 = mux_23441(v_18158);
  assign v_23443 = v_23444 | v_23446;
  assign v_23444 = mux_23444(v_23445);
  assign v_23445 = ~act_18134;
  assign v_23446 = v_23447 | v_23448;
  assign v_23447 = mux_23447(v_18135);
  assign v_23448 = mux_23448(v_18141);
  assign v_23449 = mux_23449(v_18114);
  assign v_23451 = v_23452 | v_23454;
  assign v_23452 = mux_23452(v_23453);
  assign v_23453 = ~act_18034;
  assign v_23454 = v_23455 | v_23463;
  assign v_23455 = mux_23455(v_18035);
  assign v_23457 = v_23458 | v_23460;
  assign v_23458 = mux_23458(v_23459);
  assign v_23459 = ~act_18078;
  assign v_23460 = v_23461 | v_23462;
  assign v_23461 = mux_23461(v_18079);
  assign v_23462 = mux_23462(v_18085);
  assign v_23463 = mux_23463(v_18065);
  assign v_23465 = v_23466 | v_23468;
  assign v_23466 = mux_23466(v_23467);
  assign v_23467 = ~act_18041;
  assign v_23468 = v_23469 | v_23470;
  assign v_23469 = mux_23469(v_18042);
  assign v_23470 = mux_23470(v_18048);
  assign v_23471 = mux_23471(v_18014);
  assign v_23473 = v_23474 | v_23476;
  assign v_23474 = mux_23474(v_23475);
  assign v_23475 = ~act_17822;
  assign v_23476 = v_23477 | v_23499;
  assign v_23477 = mux_23477(v_17823);
  assign v_23479 = v_23480 | v_23482;
  assign v_23480 = mux_23480(v_23481);
  assign v_23481 = ~act_17922;
  assign v_23482 = v_23483 | v_23491;
  assign v_23483 = mux_23483(v_17923);
  assign v_23485 = v_23486 | v_23488;
  assign v_23486 = mux_23486(v_23487);
  assign v_23487 = ~act_17966;
  assign v_23488 = v_23489 | v_23490;
  assign v_23489 = mux_23489(v_17967);
  assign v_23490 = mux_23490(v_17973);
  assign v_23491 = mux_23491(v_17953);
  assign v_23493 = v_23494 | v_23496;
  assign v_23494 = mux_23494(v_23495);
  assign v_23495 = ~act_17929;
  assign v_23496 = v_23497 | v_23498;
  assign v_23497 = mux_23497(v_17930);
  assign v_23498 = mux_23498(v_17936);
  assign v_23499 = mux_23499(v_17909);
  assign v_23501 = v_23502 | v_23504;
  assign v_23502 = mux_23502(v_23503);
  assign v_23503 = ~act_17829;
  assign v_23504 = v_23505 | v_23513;
  assign v_23505 = mux_23505(v_17830);
  assign v_23507 = v_23508 | v_23510;
  assign v_23508 = mux_23508(v_23509);
  assign v_23509 = ~act_17873;
  assign v_23510 = v_23511 | v_23512;
  assign v_23511 = mux_23511(v_17874);
  assign v_23512 = mux_23512(v_17880);
  assign v_23513 = mux_23513(v_17860);
  assign v_23515 = v_23516 | v_23518;
  assign v_23516 = mux_23516(v_23517);
  assign v_23517 = ~act_17836;
  assign v_23518 = v_23519 | v_23520;
  assign v_23519 = mux_23519(v_17837);
  assign v_23520 = mux_23520(v_17843);
  assign v_23521 = mux_23521(v_17795);
  assign v_23523 = v_23524 | v_23526;
  assign v_23524 = mux_23524(v_23525);
  assign v_23525 = ~act_16931;
  assign v_23526 = v_23527 | v_23633;
  assign v_23527 = mux_23527(v_16932);
  assign v_23529 = v_23530 | v_23532;
  assign v_23530 = mux_23530(v_23531);
  assign v_23531 = ~act_17367;
  assign v_23532 = v_23533 | v_23583;
  assign v_23533 = mux_23533(v_17368);
  assign v_23535 = v_23536 | v_23538;
  assign v_23536 = mux_23536(v_23537);
  assign v_23537 = ~act_17579;
  assign v_23538 = v_23539 | v_23561;
  assign v_23539 = mux_23539(v_17580);
  assign v_23541 = v_23542 | v_23544;
  assign v_23542 = mux_23542(v_23543);
  assign v_23543 = ~act_17679;
  assign v_23544 = v_23545 | v_23553;
  assign v_23545 = mux_23545(v_17680);
  assign v_23547 = v_23548 | v_23550;
  assign v_23548 = mux_23548(v_23549);
  assign v_23549 = ~act_17723;
  assign v_23550 = v_23551 | v_23552;
  assign v_23551 = mux_23551(v_17724);
  assign v_23552 = mux_23552(v_17730);
  assign v_23553 = mux_23553(v_17710);
  assign v_23555 = v_23556 | v_23558;
  assign v_23556 = mux_23556(v_23557);
  assign v_23557 = ~act_17686;
  assign v_23558 = v_23559 | v_23560;
  assign v_23559 = mux_23559(v_17687);
  assign v_23560 = mux_23560(v_17693);
  assign v_23561 = mux_23561(v_17666);
  assign v_23563 = v_23564 | v_23566;
  assign v_23564 = mux_23564(v_23565);
  assign v_23565 = ~act_17586;
  assign v_23566 = v_23567 | v_23575;
  assign v_23567 = mux_23567(v_17587);
  assign v_23569 = v_23570 | v_23572;
  assign v_23570 = mux_23570(v_23571);
  assign v_23571 = ~act_17630;
  assign v_23572 = v_23573 | v_23574;
  assign v_23573 = mux_23573(v_17631);
  assign v_23574 = mux_23574(v_17637);
  assign v_23575 = mux_23575(v_17617);
  assign v_23577 = v_23578 | v_23580;
  assign v_23578 = mux_23578(v_23579);
  assign v_23579 = ~act_17593;
  assign v_23580 = v_23581 | v_23582;
  assign v_23581 = mux_23581(v_17594);
  assign v_23582 = mux_23582(v_17600);
  assign v_23583 = mux_23583(v_17566);
  assign v_23585 = v_23586 | v_23588;
  assign v_23586 = mux_23586(v_23587);
  assign v_23587 = ~act_17374;
  assign v_23588 = v_23589 | v_23611;
  assign v_23589 = mux_23589(v_17375);
  assign v_23591 = v_23592 | v_23594;
  assign v_23592 = mux_23592(v_23593);
  assign v_23593 = ~act_17474;
  assign v_23594 = v_23595 | v_23603;
  assign v_23595 = mux_23595(v_17475);
  assign v_23597 = v_23598 | v_23600;
  assign v_23598 = mux_23598(v_23599);
  assign v_23599 = ~act_17518;
  assign v_23600 = v_23601 | v_23602;
  assign v_23601 = mux_23601(v_17519);
  assign v_23602 = mux_23602(v_17525);
  assign v_23603 = mux_23603(v_17505);
  assign v_23605 = v_23606 | v_23608;
  assign v_23606 = mux_23606(v_23607);
  assign v_23607 = ~act_17481;
  assign v_23608 = v_23609 | v_23610;
  assign v_23609 = mux_23609(v_17482);
  assign v_23610 = mux_23610(v_17488);
  assign v_23611 = mux_23611(v_17461);
  assign v_23613 = v_23614 | v_23616;
  assign v_23614 = mux_23614(v_23615);
  assign v_23615 = ~act_17381;
  assign v_23616 = v_23617 | v_23625;
  assign v_23617 = mux_23617(v_17382);
  assign v_23619 = v_23620 | v_23622;
  assign v_23620 = mux_23620(v_23621);
  assign v_23621 = ~act_17425;
  assign v_23622 = v_23623 | v_23624;
  assign v_23623 = mux_23623(v_17426);
  assign v_23624 = mux_23624(v_17432);
  assign v_23625 = mux_23625(v_17412);
  assign v_23627 = v_23628 | v_23630;
  assign v_23628 = mux_23628(v_23629);
  assign v_23629 = ~act_17388;
  assign v_23630 = v_23631 | v_23632;
  assign v_23631 = mux_23631(v_17389);
  assign v_23632 = mux_23632(v_17395);
  assign v_23633 = mux_23633(v_17354);
  assign v_23635 = v_23636 | v_23638;
  assign v_23636 = mux_23636(v_23637);
  assign v_23637 = ~act_16938;
  assign v_23638 = v_23639 | v_23689;
  assign v_23639 = mux_23639(v_16939);
  assign v_23641 = v_23642 | v_23644;
  assign v_23642 = mux_23642(v_23643);
  assign v_23643 = ~act_17150;
  assign v_23644 = v_23645 | v_23667;
  assign v_23645 = mux_23645(v_17151);
  assign v_23647 = v_23648 | v_23650;
  assign v_23648 = mux_23648(v_23649);
  assign v_23649 = ~act_17250;
  assign v_23650 = v_23651 | v_23659;
  assign v_23651 = mux_23651(v_17251);
  assign v_23653 = v_23654 | v_23656;
  assign v_23654 = mux_23654(v_23655);
  assign v_23655 = ~act_17294;
  assign v_23656 = v_23657 | v_23658;
  assign v_23657 = mux_23657(v_17295);
  assign v_23658 = mux_23658(v_17301);
  assign v_23659 = mux_23659(v_17281);
  assign v_23661 = v_23662 | v_23664;
  assign v_23662 = mux_23662(v_23663);
  assign v_23663 = ~act_17257;
  assign v_23664 = v_23665 | v_23666;
  assign v_23665 = mux_23665(v_17258);
  assign v_23666 = mux_23666(v_17264);
  assign v_23667 = mux_23667(v_17237);
  assign v_23669 = v_23670 | v_23672;
  assign v_23670 = mux_23670(v_23671);
  assign v_23671 = ~act_17157;
  assign v_23672 = v_23673 | v_23681;
  assign v_23673 = mux_23673(v_17158);
  assign v_23675 = v_23676 | v_23678;
  assign v_23676 = mux_23676(v_23677);
  assign v_23677 = ~act_17201;
  assign v_23678 = v_23679 | v_23680;
  assign v_23679 = mux_23679(v_17202);
  assign v_23680 = mux_23680(v_17208);
  assign v_23681 = mux_23681(v_17188);
  assign v_23683 = v_23684 | v_23686;
  assign v_23684 = mux_23684(v_23685);
  assign v_23685 = ~act_17164;
  assign v_23686 = v_23687 | v_23688;
  assign v_23687 = mux_23687(v_17165);
  assign v_23688 = mux_23688(v_17171);
  assign v_23689 = mux_23689(v_17137);
  assign v_23691 = v_23692 | v_23694;
  assign v_23692 = mux_23692(v_23693);
  assign v_23693 = ~act_16945;
  assign v_23694 = v_23695 | v_23717;
  assign v_23695 = mux_23695(v_16946);
  assign v_23697 = v_23698 | v_23700;
  assign v_23698 = mux_23698(v_23699);
  assign v_23699 = ~act_17045;
  assign v_23700 = v_23701 | v_23709;
  assign v_23701 = mux_23701(v_17046);
  assign v_23703 = v_23704 | v_23706;
  assign v_23704 = mux_23704(v_23705);
  assign v_23705 = ~act_17089;
  assign v_23706 = v_23707 | v_23708;
  assign v_23707 = mux_23707(v_17090);
  assign v_23708 = mux_23708(v_17096);
  assign v_23709 = mux_23709(v_17076);
  assign v_23711 = v_23712 | v_23714;
  assign v_23712 = mux_23712(v_23713);
  assign v_23713 = ~act_17052;
  assign v_23714 = v_23715 | v_23716;
  assign v_23715 = mux_23715(v_17053);
  assign v_23716 = mux_23716(v_17059);
  assign v_23717 = mux_23717(v_17032);
  assign v_23719 = v_23720 | v_23722;
  assign v_23720 = mux_23720(v_23721);
  assign v_23721 = ~act_16952;
  assign v_23722 = v_23723 | v_23731;
  assign v_23723 = mux_23723(v_16953);
  assign v_23725 = v_23726 | v_23728;
  assign v_23726 = mux_23726(v_23727);
  assign v_23727 = ~act_16996;
  assign v_23728 = v_23729 | v_23730;
  assign v_23729 = mux_23729(v_16997);
  assign v_23730 = mux_23730(v_17003);
  assign v_23731 = mux_23731(v_16983);
  assign v_23733 = v_23734 | v_23736;
  assign v_23734 = mux_23734(v_23735);
  assign v_23735 = ~act_16959;
  assign v_23736 = v_23737 | v_23738;
  assign v_23737 = mux_23737(v_16960);
  assign v_23738 = mux_23738(v_16966);
  assign v_23739 = mux_23739(v_16911);
  assign v_23741 = v_23742 | v_23744;
  assign v_23742 = mux_23742(v_23743);
  assign v_23743 = ~act_15151;
  assign v_23744 = v_23745 | v_23963;
  assign v_23745 = mux_23745(v_15152);
  assign v_23747 = v_23748 | v_23750;
  assign v_23748 = mux_23748(v_23749);
  assign v_23749 = ~act_16035;
  assign v_23750 = v_23751 | v_23857;
  assign v_23751 = mux_23751(v_16036);
  assign v_23753 = v_23754 | v_23756;
  assign v_23754 = mux_23754(v_23755);
  assign v_23755 = ~act_16471;
  assign v_23756 = v_23757 | v_23807;
  assign v_23757 = mux_23757(v_16472);
  assign v_23759 = v_23760 | v_23762;
  assign v_23760 = mux_23760(v_23761);
  assign v_23761 = ~act_16683;
  assign v_23762 = v_23763 | v_23785;
  assign v_23763 = mux_23763(v_16684);
  assign v_23765 = v_23766 | v_23768;
  assign v_23766 = mux_23766(v_23767);
  assign v_23767 = ~act_16783;
  assign v_23768 = v_23769 | v_23777;
  assign v_23769 = mux_23769(v_16784);
  assign v_23771 = v_23772 | v_23774;
  assign v_23772 = mux_23772(v_23773);
  assign v_23773 = ~act_16827;
  assign v_23774 = v_23775 | v_23776;
  assign v_23775 = mux_23775(v_16828);
  assign v_23776 = mux_23776(v_16834);
  assign v_23777 = mux_23777(v_16814);
  assign v_23779 = v_23780 | v_23782;
  assign v_23780 = mux_23780(v_23781);
  assign v_23781 = ~act_16790;
  assign v_23782 = v_23783 | v_23784;
  assign v_23783 = mux_23783(v_16791);
  assign v_23784 = mux_23784(v_16797);
  assign v_23785 = mux_23785(v_16770);
  assign v_23787 = v_23788 | v_23790;
  assign v_23788 = mux_23788(v_23789);
  assign v_23789 = ~act_16690;
  assign v_23790 = v_23791 | v_23799;
  assign v_23791 = mux_23791(v_16691);
  assign v_23793 = v_23794 | v_23796;
  assign v_23794 = mux_23794(v_23795);
  assign v_23795 = ~act_16734;
  assign v_23796 = v_23797 | v_23798;
  assign v_23797 = mux_23797(v_16735);
  assign v_23798 = mux_23798(v_16741);
  assign v_23799 = mux_23799(v_16721);
  assign v_23801 = v_23802 | v_23804;
  assign v_23802 = mux_23802(v_23803);
  assign v_23803 = ~act_16697;
  assign v_23804 = v_23805 | v_23806;
  assign v_23805 = mux_23805(v_16698);
  assign v_23806 = mux_23806(v_16704);
  assign v_23807 = mux_23807(v_16670);
  assign v_23809 = v_23810 | v_23812;
  assign v_23810 = mux_23810(v_23811);
  assign v_23811 = ~act_16478;
  assign v_23812 = v_23813 | v_23835;
  assign v_23813 = mux_23813(v_16479);
  assign v_23815 = v_23816 | v_23818;
  assign v_23816 = mux_23816(v_23817);
  assign v_23817 = ~act_16578;
  assign v_23818 = v_23819 | v_23827;
  assign v_23819 = mux_23819(v_16579);
  assign v_23821 = v_23822 | v_23824;
  assign v_23822 = mux_23822(v_23823);
  assign v_23823 = ~act_16622;
  assign v_23824 = v_23825 | v_23826;
  assign v_23825 = mux_23825(v_16623);
  assign v_23826 = mux_23826(v_16629);
  assign v_23827 = mux_23827(v_16609);
  assign v_23829 = v_23830 | v_23832;
  assign v_23830 = mux_23830(v_23831);
  assign v_23831 = ~act_16585;
  assign v_23832 = v_23833 | v_23834;
  assign v_23833 = mux_23833(v_16586);
  assign v_23834 = mux_23834(v_16592);
  assign v_23835 = mux_23835(v_16565);
  assign v_23837 = v_23838 | v_23840;
  assign v_23838 = mux_23838(v_23839);
  assign v_23839 = ~act_16485;
  assign v_23840 = v_23841 | v_23849;
  assign v_23841 = mux_23841(v_16486);
  assign v_23843 = v_23844 | v_23846;
  assign v_23844 = mux_23844(v_23845);
  assign v_23845 = ~act_16529;
  assign v_23846 = v_23847 | v_23848;
  assign v_23847 = mux_23847(v_16530);
  assign v_23848 = mux_23848(v_16536);
  assign v_23849 = mux_23849(v_16516);
  assign v_23851 = v_23852 | v_23854;
  assign v_23852 = mux_23852(v_23853);
  assign v_23853 = ~act_16492;
  assign v_23854 = v_23855 | v_23856;
  assign v_23855 = mux_23855(v_16493);
  assign v_23856 = mux_23856(v_16499);
  assign v_23857 = mux_23857(v_16458);
  assign v_23859 = v_23860 | v_23862;
  assign v_23860 = mux_23860(v_23861);
  assign v_23861 = ~act_16042;
  assign v_23862 = v_23863 | v_23913;
  assign v_23863 = mux_23863(v_16043);
  assign v_23865 = v_23866 | v_23868;
  assign v_23866 = mux_23866(v_23867);
  assign v_23867 = ~act_16254;
  assign v_23868 = v_23869 | v_23891;
  assign v_23869 = mux_23869(v_16255);
  assign v_23871 = v_23872 | v_23874;
  assign v_23872 = mux_23872(v_23873);
  assign v_23873 = ~act_16354;
  assign v_23874 = v_23875 | v_23883;
  assign v_23875 = mux_23875(v_16355);
  assign v_23877 = v_23878 | v_23880;
  assign v_23878 = mux_23878(v_23879);
  assign v_23879 = ~act_16398;
  assign v_23880 = v_23881 | v_23882;
  assign v_23881 = mux_23881(v_16399);
  assign v_23882 = mux_23882(v_16405);
  assign v_23883 = mux_23883(v_16385);
  assign v_23885 = v_23886 | v_23888;
  assign v_23886 = mux_23886(v_23887);
  assign v_23887 = ~act_16361;
  assign v_23888 = v_23889 | v_23890;
  assign v_23889 = mux_23889(v_16362);
  assign v_23890 = mux_23890(v_16368);
  assign v_23891 = mux_23891(v_16341);
  assign v_23893 = v_23894 | v_23896;
  assign v_23894 = mux_23894(v_23895);
  assign v_23895 = ~act_16261;
  assign v_23896 = v_23897 | v_23905;
  assign v_23897 = mux_23897(v_16262);
  assign v_23899 = v_23900 | v_23902;
  assign v_23900 = mux_23900(v_23901);
  assign v_23901 = ~act_16305;
  assign v_23902 = v_23903 | v_23904;
  assign v_23903 = mux_23903(v_16306);
  assign v_23904 = mux_23904(v_16312);
  assign v_23905 = mux_23905(v_16292);
  assign v_23907 = v_23908 | v_23910;
  assign v_23908 = mux_23908(v_23909);
  assign v_23909 = ~act_16268;
  assign v_23910 = v_23911 | v_23912;
  assign v_23911 = mux_23911(v_16269);
  assign v_23912 = mux_23912(v_16275);
  assign v_23913 = mux_23913(v_16241);
  assign v_23915 = v_23916 | v_23918;
  assign v_23916 = mux_23916(v_23917);
  assign v_23917 = ~act_16049;
  assign v_23918 = v_23919 | v_23941;
  assign v_23919 = mux_23919(v_16050);
  assign v_23921 = v_23922 | v_23924;
  assign v_23922 = mux_23922(v_23923);
  assign v_23923 = ~act_16149;
  assign v_23924 = v_23925 | v_23933;
  assign v_23925 = mux_23925(v_16150);
  assign v_23927 = v_23928 | v_23930;
  assign v_23928 = mux_23928(v_23929);
  assign v_23929 = ~act_16193;
  assign v_23930 = v_23931 | v_23932;
  assign v_23931 = mux_23931(v_16194);
  assign v_23932 = mux_23932(v_16200);
  assign v_23933 = mux_23933(v_16180);
  assign v_23935 = v_23936 | v_23938;
  assign v_23936 = mux_23936(v_23937);
  assign v_23937 = ~act_16156;
  assign v_23938 = v_23939 | v_23940;
  assign v_23939 = mux_23939(v_16157);
  assign v_23940 = mux_23940(v_16163);
  assign v_23941 = mux_23941(v_16136);
  assign v_23943 = v_23944 | v_23946;
  assign v_23944 = mux_23944(v_23945);
  assign v_23945 = ~act_16056;
  assign v_23946 = v_23947 | v_23955;
  assign v_23947 = mux_23947(v_16057);
  assign v_23949 = v_23950 | v_23952;
  assign v_23950 = mux_23950(v_23951);
  assign v_23951 = ~act_16100;
  assign v_23952 = v_23953 | v_23954;
  assign v_23953 = mux_23953(v_16101);
  assign v_23954 = mux_23954(v_16107);
  assign v_23955 = mux_23955(v_16087);
  assign v_23957 = v_23958 | v_23960;
  assign v_23958 = mux_23958(v_23959);
  assign v_23959 = ~act_16063;
  assign v_23960 = v_23961 | v_23962;
  assign v_23961 = mux_23961(v_16064);
  assign v_23962 = mux_23962(v_16070);
  assign v_23963 = mux_23963(v_16022);
  assign v_23965 = v_23966 | v_23968;
  assign v_23966 = mux_23966(v_23967);
  assign v_23967 = ~act_15158;
  assign v_23968 = v_23969 | v_24075;
  assign v_23969 = mux_23969(v_15159);
  assign v_23971 = v_23972 | v_23974;
  assign v_23972 = mux_23972(v_23973);
  assign v_23973 = ~act_15594;
  assign v_23974 = v_23975 | v_24025;
  assign v_23975 = mux_23975(v_15595);
  assign v_23977 = v_23978 | v_23980;
  assign v_23978 = mux_23978(v_23979);
  assign v_23979 = ~act_15806;
  assign v_23980 = v_23981 | v_24003;
  assign v_23981 = mux_23981(v_15807);
  assign v_23983 = v_23984 | v_23986;
  assign v_23984 = mux_23984(v_23985);
  assign v_23985 = ~act_15906;
  assign v_23986 = v_23987 | v_23995;
  assign v_23987 = mux_23987(v_15907);
  assign v_23989 = v_23990 | v_23992;
  assign v_23990 = mux_23990(v_23991);
  assign v_23991 = ~act_15950;
  assign v_23992 = v_23993 | v_23994;
  assign v_23993 = mux_23993(v_15951);
  assign v_23994 = mux_23994(v_15957);
  assign v_23995 = mux_23995(v_15937);
  assign v_23997 = v_23998 | v_24000;
  assign v_23998 = mux_23998(v_23999);
  assign v_23999 = ~act_15913;
  assign v_24000 = v_24001 | v_24002;
  assign v_24001 = mux_24001(v_15914);
  assign v_24002 = mux_24002(v_15920);
  assign v_24003 = mux_24003(v_15893);
  assign v_24005 = v_24006 | v_24008;
  assign v_24006 = mux_24006(v_24007);
  assign v_24007 = ~act_15813;
  assign v_24008 = v_24009 | v_24017;
  assign v_24009 = mux_24009(v_15814);
  assign v_24011 = v_24012 | v_24014;
  assign v_24012 = mux_24012(v_24013);
  assign v_24013 = ~act_15857;
  assign v_24014 = v_24015 | v_24016;
  assign v_24015 = mux_24015(v_15858);
  assign v_24016 = mux_24016(v_15864);
  assign v_24017 = mux_24017(v_15844);
  assign v_24019 = v_24020 | v_24022;
  assign v_24020 = mux_24020(v_24021);
  assign v_24021 = ~act_15820;
  assign v_24022 = v_24023 | v_24024;
  assign v_24023 = mux_24023(v_15821);
  assign v_24024 = mux_24024(v_15827);
  assign v_24025 = mux_24025(v_15793);
  assign v_24027 = v_24028 | v_24030;
  assign v_24028 = mux_24028(v_24029);
  assign v_24029 = ~act_15601;
  assign v_24030 = v_24031 | v_24053;
  assign v_24031 = mux_24031(v_15602);
  assign v_24033 = v_24034 | v_24036;
  assign v_24034 = mux_24034(v_24035);
  assign v_24035 = ~act_15701;
  assign v_24036 = v_24037 | v_24045;
  assign v_24037 = mux_24037(v_15702);
  assign v_24039 = v_24040 | v_24042;
  assign v_24040 = mux_24040(v_24041);
  assign v_24041 = ~act_15745;
  assign v_24042 = v_24043 | v_24044;
  assign v_24043 = mux_24043(v_15746);
  assign v_24044 = mux_24044(v_15752);
  assign v_24045 = mux_24045(v_15732);
  assign v_24047 = v_24048 | v_24050;
  assign v_24048 = mux_24048(v_24049);
  assign v_24049 = ~act_15708;
  assign v_24050 = v_24051 | v_24052;
  assign v_24051 = mux_24051(v_15709);
  assign v_24052 = mux_24052(v_15715);
  assign v_24053 = mux_24053(v_15688);
  assign v_24055 = v_24056 | v_24058;
  assign v_24056 = mux_24056(v_24057);
  assign v_24057 = ~act_15608;
  assign v_24058 = v_24059 | v_24067;
  assign v_24059 = mux_24059(v_15609);
  assign v_24061 = v_24062 | v_24064;
  assign v_24062 = mux_24062(v_24063);
  assign v_24063 = ~act_15652;
  assign v_24064 = v_24065 | v_24066;
  assign v_24065 = mux_24065(v_15653);
  assign v_24066 = mux_24066(v_15659);
  assign v_24067 = mux_24067(v_15639);
  assign v_24069 = v_24070 | v_24072;
  assign v_24070 = mux_24070(v_24071);
  assign v_24071 = ~act_15615;
  assign v_24072 = v_24073 | v_24074;
  assign v_24073 = mux_24073(v_15616);
  assign v_24074 = mux_24074(v_15622);
  assign v_24075 = mux_24075(v_15581);
  assign v_24077 = v_24078 | v_24080;
  assign v_24078 = mux_24078(v_24079);
  assign v_24079 = ~act_15165;
  assign v_24080 = v_24081 | v_24131;
  assign v_24081 = mux_24081(v_15166);
  assign v_24083 = v_24084 | v_24086;
  assign v_24084 = mux_24084(v_24085);
  assign v_24085 = ~act_15377;
  assign v_24086 = v_24087 | v_24109;
  assign v_24087 = mux_24087(v_15378);
  assign v_24089 = v_24090 | v_24092;
  assign v_24090 = mux_24090(v_24091);
  assign v_24091 = ~act_15477;
  assign v_24092 = v_24093 | v_24101;
  assign v_24093 = mux_24093(v_15478);
  assign v_24095 = v_24096 | v_24098;
  assign v_24096 = mux_24096(v_24097);
  assign v_24097 = ~act_15521;
  assign v_24098 = v_24099 | v_24100;
  assign v_24099 = mux_24099(v_15522);
  assign v_24100 = mux_24100(v_15528);
  assign v_24101 = mux_24101(v_15508);
  assign v_24103 = v_24104 | v_24106;
  assign v_24104 = mux_24104(v_24105);
  assign v_24105 = ~act_15484;
  assign v_24106 = v_24107 | v_24108;
  assign v_24107 = mux_24107(v_15485);
  assign v_24108 = mux_24108(v_15491);
  assign v_24109 = mux_24109(v_15464);
  assign v_24111 = v_24112 | v_24114;
  assign v_24112 = mux_24112(v_24113);
  assign v_24113 = ~act_15384;
  assign v_24114 = v_24115 | v_24123;
  assign v_24115 = mux_24115(v_15385);
  assign v_24117 = v_24118 | v_24120;
  assign v_24118 = mux_24118(v_24119);
  assign v_24119 = ~act_15428;
  assign v_24120 = v_24121 | v_24122;
  assign v_24121 = mux_24121(v_15429);
  assign v_24122 = mux_24122(v_15435);
  assign v_24123 = mux_24123(v_15415);
  assign v_24125 = v_24126 | v_24128;
  assign v_24126 = mux_24126(v_24127);
  assign v_24127 = ~act_15391;
  assign v_24128 = v_24129 | v_24130;
  assign v_24129 = mux_24129(v_15392);
  assign v_24130 = mux_24130(v_15398);
  assign v_24131 = mux_24131(v_15364);
  assign v_24133 = v_24134 | v_24136;
  assign v_24134 = mux_24134(v_24135);
  assign v_24135 = ~act_15172;
  assign v_24136 = v_24137 | v_24159;
  assign v_24137 = mux_24137(v_15173);
  assign v_24139 = v_24140 | v_24142;
  assign v_24140 = mux_24140(v_24141);
  assign v_24141 = ~act_15272;
  assign v_24142 = v_24143 | v_24151;
  assign v_24143 = mux_24143(v_15273);
  assign v_24145 = v_24146 | v_24148;
  assign v_24146 = mux_24146(v_24147);
  assign v_24147 = ~act_15316;
  assign v_24148 = v_24149 | v_24150;
  assign v_24149 = mux_24149(v_15317);
  assign v_24150 = mux_24150(v_15323);
  assign v_24151 = mux_24151(v_15303);
  assign v_24153 = v_24154 | v_24156;
  assign v_24154 = mux_24154(v_24155);
  assign v_24155 = ~act_15279;
  assign v_24156 = v_24157 | v_24158;
  assign v_24157 = mux_24157(v_15280);
  assign v_24158 = mux_24158(v_15286);
  assign v_24159 = mux_24159(v_15259);
  assign v_24161 = v_24162 | v_24164;
  assign v_24162 = mux_24162(v_24163);
  assign v_24163 = ~act_15179;
  assign v_24164 = v_24165 | v_24173;
  assign v_24165 = mux_24165(v_15180);
  assign v_24167 = v_24168 | v_24170;
  assign v_24168 = mux_24168(v_24169);
  assign v_24169 = ~act_15223;
  assign v_24170 = v_24171 | v_24172;
  assign v_24171 = mux_24171(v_15224);
  assign v_24172 = mux_24172(v_15230);
  assign v_24173 = mux_24173(v_15210);
  assign v_24175 = v_24176 | v_24178;
  assign v_24176 = mux_24176(v_24177);
  assign v_24177 = ~act_15186;
  assign v_24178 = v_24179 | v_24180;
  assign v_24179 = mux_24179(v_15187);
  assign v_24180 = mux_24180(v_15193);
  assign v_24181 = mux_24181(v_15124);
  assign v_24183 = v_24184 | v_24186;
  assign v_24184 = mux_24184(v_24185);
  assign v_24185 = ~act_7988;
  assign v_24186 = v_24187 | v_25077;
  assign v_24187 = mux_24187(v_7989);
  assign v_24189 = v_24190 | v_24192;
  assign v_24190 = mux_24190(v_24191);
  assign v_24191 = ~act_11560;
  assign v_24192 = v_24193 | v_24635;
  assign v_24193 = mux_24193(v_11561);
  assign v_24195 = v_24196 | v_24198;
  assign v_24196 = mux_24196(v_24197);
  assign v_24197 = ~act_13340;
  assign v_24198 = v_24199 | v_24417;
  assign v_24199 = mux_24199(v_13341);
  assign v_24201 = v_24202 | v_24204;
  assign v_24202 = mux_24202(v_24203);
  assign v_24203 = ~act_14224;
  assign v_24204 = v_24205 | v_24311;
  assign v_24205 = mux_24205(v_14225);
  assign v_24207 = v_24208 | v_24210;
  assign v_24208 = mux_24208(v_24209);
  assign v_24209 = ~act_14660;
  assign v_24210 = v_24211 | v_24261;
  assign v_24211 = mux_24211(v_14661);
  assign v_24213 = v_24214 | v_24216;
  assign v_24214 = mux_24214(v_24215);
  assign v_24215 = ~act_14872;
  assign v_24216 = v_24217 | v_24239;
  assign v_24217 = mux_24217(v_14873);
  assign v_24219 = v_24220 | v_24222;
  assign v_24220 = mux_24220(v_24221);
  assign v_24221 = ~act_14972;
  assign v_24222 = v_24223 | v_24231;
  assign v_24223 = mux_24223(v_14973);
  assign v_24225 = v_24226 | v_24228;
  assign v_24226 = mux_24226(v_24227);
  assign v_24227 = ~act_15016;
  assign v_24228 = v_24229 | v_24230;
  assign v_24229 = mux_24229(v_15017);
  assign v_24230 = mux_24230(v_15023);
  assign v_24231 = mux_24231(v_15003);
  assign v_24233 = v_24234 | v_24236;
  assign v_24234 = mux_24234(v_24235);
  assign v_24235 = ~act_14979;
  assign v_24236 = v_24237 | v_24238;
  assign v_24237 = mux_24237(v_14980);
  assign v_24238 = mux_24238(v_14986);
  assign v_24239 = mux_24239(v_14959);
  assign v_24241 = v_24242 | v_24244;
  assign v_24242 = mux_24242(v_24243);
  assign v_24243 = ~act_14879;
  assign v_24244 = v_24245 | v_24253;
  assign v_24245 = mux_24245(v_14880);
  assign v_24247 = v_24248 | v_24250;
  assign v_24248 = mux_24248(v_24249);
  assign v_24249 = ~act_14923;
  assign v_24250 = v_24251 | v_24252;
  assign v_24251 = mux_24251(v_14924);
  assign v_24252 = mux_24252(v_14930);
  assign v_24253 = mux_24253(v_14910);
  assign v_24255 = v_24256 | v_24258;
  assign v_24256 = mux_24256(v_24257);
  assign v_24257 = ~act_14886;
  assign v_24258 = v_24259 | v_24260;
  assign v_24259 = mux_24259(v_14887);
  assign v_24260 = mux_24260(v_14893);
  assign v_24261 = mux_24261(v_14859);
  assign v_24263 = v_24264 | v_24266;
  assign v_24264 = mux_24264(v_24265);
  assign v_24265 = ~act_14667;
  assign v_24266 = v_24267 | v_24289;
  assign v_24267 = mux_24267(v_14668);
  assign v_24269 = v_24270 | v_24272;
  assign v_24270 = mux_24270(v_24271);
  assign v_24271 = ~act_14767;
  assign v_24272 = v_24273 | v_24281;
  assign v_24273 = mux_24273(v_14768);
  assign v_24275 = v_24276 | v_24278;
  assign v_24276 = mux_24276(v_24277);
  assign v_24277 = ~act_14811;
  assign v_24278 = v_24279 | v_24280;
  assign v_24279 = mux_24279(v_14812);
  assign v_24280 = mux_24280(v_14818);
  assign v_24281 = mux_24281(v_14798);
  assign v_24283 = v_24284 | v_24286;
  assign v_24284 = mux_24284(v_24285);
  assign v_24285 = ~act_14774;
  assign v_24286 = v_24287 | v_24288;
  assign v_24287 = mux_24287(v_14775);
  assign v_24288 = mux_24288(v_14781);
  assign v_24289 = mux_24289(v_14754);
  assign v_24291 = v_24292 | v_24294;
  assign v_24292 = mux_24292(v_24293);
  assign v_24293 = ~act_14674;
  assign v_24294 = v_24295 | v_24303;
  assign v_24295 = mux_24295(v_14675);
  assign v_24297 = v_24298 | v_24300;
  assign v_24298 = mux_24298(v_24299);
  assign v_24299 = ~act_14718;
  assign v_24300 = v_24301 | v_24302;
  assign v_24301 = mux_24301(v_14719);
  assign v_24302 = mux_24302(v_14725);
  assign v_24303 = mux_24303(v_14705);
  assign v_24305 = v_24306 | v_24308;
  assign v_24306 = mux_24306(v_24307);
  assign v_24307 = ~act_14681;
  assign v_24308 = v_24309 | v_24310;
  assign v_24309 = mux_24309(v_14682);
  assign v_24310 = mux_24310(v_14688);
  assign v_24311 = mux_24311(v_14647);
  assign v_24313 = v_24314 | v_24316;
  assign v_24314 = mux_24314(v_24315);
  assign v_24315 = ~act_14231;
  assign v_24316 = v_24317 | v_24367;
  assign v_24317 = mux_24317(v_14232);
  assign v_24319 = v_24320 | v_24322;
  assign v_24320 = mux_24320(v_24321);
  assign v_24321 = ~act_14443;
  assign v_24322 = v_24323 | v_24345;
  assign v_24323 = mux_24323(v_14444);
  assign v_24325 = v_24326 | v_24328;
  assign v_24326 = mux_24326(v_24327);
  assign v_24327 = ~act_14543;
  assign v_24328 = v_24329 | v_24337;
  assign v_24329 = mux_24329(v_14544);
  assign v_24331 = v_24332 | v_24334;
  assign v_24332 = mux_24332(v_24333);
  assign v_24333 = ~act_14587;
  assign v_24334 = v_24335 | v_24336;
  assign v_24335 = mux_24335(v_14588);
  assign v_24336 = mux_24336(v_14594);
  assign v_24337 = mux_24337(v_14574);
  assign v_24339 = v_24340 | v_24342;
  assign v_24340 = mux_24340(v_24341);
  assign v_24341 = ~act_14550;
  assign v_24342 = v_24343 | v_24344;
  assign v_24343 = mux_24343(v_14551);
  assign v_24344 = mux_24344(v_14557);
  assign v_24345 = mux_24345(v_14530);
  assign v_24347 = v_24348 | v_24350;
  assign v_24348 = mux_24348(v_24349);
  assign v_24349 = ~act_14450;
  assign v_24350 = v_24351 | v_24359;
  assign v_24351 = mux_24351(v_14451);
  assign v_24353 = v_24354 | v_24356;
  assign v_24354 = mux_24354(v_24355);
  assign v_24355 = ~act_14494;
  assign v_24356 = v_24357 | v_24358;
  assign v_24357 = mux_24357(v_14495);
  assign v_24358 = mux_24358(v_14501);
  assign v_24359 = mux_24359(v_14481);
  assign v_24361 = v_24362 | v_24364;
  assign v_24362 = mux_24362(v_24363);
  assign v_24363 = ~act_14457;
  assign v_24364 = v_24365 | v_24366;
  assign v_24365 = mux_24365(v_14458);
  assign v_24366 = mux_24366(v_14464);
  assign v_24367 = mux_24367(v_14430);
  assign v_24369 = v_24370 | v_24372;
  assign v_24370 = mux_24370(v_24371);
  assign v_24371 = ~act_14238;
  assign v_24372 = v_24373 | v_24395;
  assign v_24373 = mux_24373(v_14239);
  assign v_24375 = v_24376 | v_24378;
  assign v_24376 = mux_24376(v_24377);
  assign v_24377 = ~act_14338;
  assign v_24378 = v_24379 | v_24387;
  assign v_24379 = mux_24379(v_14339);
  assign v_24381 = v_24382 | v_24384;
  assign v_24382 = mux_24382(v_24383);
  assign v_24383 = ~act_14382;
  assign v_24384 = v_24385 | v_24386;
  assign v_24385 = mux_24385(v_14383);
  assign v_24386 = mux_24386(v_14389);
  assign v_24387 = mux_24387(v_14369);
  assign v_24389 = v_24390 | v_24392;
  assign v_24390 = mux_24390(v_24391);
  assign v_24391 = ~act_14345;
  assign v_24392 = v_24393 | v_24394;
  assign v_24393 = mux_24393(v_14346);
  assign v_24394 = mux_24394(v_14352);
  assign v_24395 = mux_24395(v_14325);
  assign v_24397 = v_24398 | v_24400;
  assign v_24398 = mux_24398(v_24399);
  assign v_24399 = ~act_14245;
  assign v_24400 = v_24401 | v_24409;
  assign v_24401 = mux_24401(v_14246);
  assign v_24403 = v_24404 | v_24406;
  assign v_24404 = mux_24404(v_24405);
  assign v_24405 = ~act_14289;
  assign v_24406 = v_24407 | v_24408;
  assign v_24407 = mux_24407(v_14290);
  assign v_24408 = mux_24408(v_14296);
  assign v_24409 = mux_24409(v_14276);
  assign v_24411 = v_24412 | v_24414;
  assign v_24412 = mux_24412(v_24413);
  assign v_24413 = ~act_14252;
  assign v_24414 = v_24415 | v_24416;
  assign v_24415 = mux_24415(v_14253);
  assign v_24416 = mux_24416(v_14259);
  assign v_24417 = mux_24417(v_14211);
  assign v_24419 = v_24420 | v_24422;
  assign v_24420 = mux_24420(v_24421);
  assign v_24421 = ~act_13347;
  assign v_24422 = v_24423 | v_24529;
  assign v_24423 = mux_24423(v_13348);
  assign v_24425 = v_24426 | v_24428;
  assign v_24426 = mux_24426(v_24427);
  assign v_24427 = ~act_13783;
  assign v_24428 = v_24429 | v_24479;
  assign v_24429 = mux_24429(v_13784);
  assign v_24431 = v_24432 | v_24434;
  assign v_24432 = mux_24432(v_24433);
  assign v_24433 = ~act_13995;
  assign v_24434 = v_24435 | v_24457;
  assign v_24435 = mux_24435(v_13996);
  assign v_24437 = v_24438 | v_24440;
  assign v_24438 = mux_24438(v_24439);
  assign v_24439 = ~act_14095;
  assign v_24440 = v_24441 | v_24449;
  assign v_24441 = mux_24441(v_14096);
  assign v_24443 = v_24444 | v_24446;
  assign v_24444 = mux_24444(v_24445);
  assign v_24445 = ~act_14139;
  assign v_24446 = v_24447 | v_24448;
  assign v_24447 = mux_24447(v_14140);
  assign v_24448 = mux_24448(v_14146);
  assign v_24449 = mux_24449(v_14126);
  assign v_24451 = v_24452 | v_24454;
  assign v_24452 = mux_24452(v_24453);
  assign v_24453 = ~act_14102;
  assign v_24454 = v_24455 | v_24456;
  assign v_24455 = mux_24455(v_14103);
  assign v_24456 = mux_24456(v_14109);
  assign v_24457 = mux_24457(v_14082);
  assign v_24459 = v_24460 | v_24462;
  assign v_24460 = mux_24460(v_24461);
  assign v_24461 = ~act_14002;
  assign v_24462 = v_24463 | v_24471;
  assign v_24463 = mux_24463(v_14003);
  assign v_24465 = v_24466 | v_24468;
  assign v_24466 = mux_24466(v_24467);
  assign v_24467 = ~act_14046;
  assign v_24468 = v_24469 | v_24470;
  assign v_24469 = mux_24469(v_14047);
  assign v_24470 = mux_24470(v_14053);
  assign v_24471 = mux_24471(v_14033);
  assign v_24473 = v_24474 | v_24476;
  assign v_24474 = mux_24474(v_24475);
  assign v_24475 = ~act_14009;
  assign v_24476 = v_24477 | v_24478;
  assign v_24477 = mux_24477(v_14010);
  assign v_24478 = mux_24478(v_14016);
  assign v_24479 = mux_24479(v_13982);
  assign v_24481 = v_24482 | v_24484;
  assign v_24482 = mux_24482(v_24483);
  assign v_24483 = ~act_13790;
  assign v_24484 = v_24485 | v_24507;
  assign v_24485 = mux_24485(v_13791);
  assign v_24487 = v_24488 | v_24490;
  assign v_24488 = mux_24488(v_24489);
  assign v_24489 = ~act_13890;
  assign v_24490 = v_24491 | v_24499;
  assign v_24491 = mux_24491(v_13891);
  assign v_24493 = v_24494 | v_24496;
  assign v_24494 = mux_24494(v_24495);
  assign v_24495 = ~act_13934;
  assign v_24496 = v_24497 | v_24498;
  assign v_24497 = mux_24497(v_13935);
  assign v_24498 = mux_24498(v_13941);
  assign v_24499 = mux_24499(v_13921);
  assign v_24501 = v_24502 | v_24504;
  assign v_24502 = mux_24502(v_24503);
  assign v_24503 = ~act_13897;
  assign v_24504 = v_24505 | v_24506;
  assign v_24505 = mux_24505(v_13898);
  assign v_24506 = mux_24506(v_13904);
  assign v_24507 = mux_24507(v_13877);
  assign v_24509 = v_24510 | v_24512;
  assign v_24510 = mux_24510(v_24511);
  assign v_24511 = ~act_13797;
  assign v_24512 = v_24513 | v_24521;
  assign v_24513 = mux_24513(v_13798);
  assign v_24515 = v_24516 | v_24518;
  assign v_24516 = mux_24516(v_24517);
  assign v_24517 = ~act_13841;
  assign v_24518 = v_24519 | v_24520;
  assign v_24519 = mux_24519(v_13842);
  assign v_24520 = mux_24520(v_13848);
  assign v_24521 = mux_24521(v_13828);
  assign v_24523 = v_24524 | v_24526;
  assign v_24524 = mux_24524(v_24525);
  assign v_24525 = ~act_13804;
  assign v_24526 = v_24527 | v_24528;
  assign v_24527 = mux_24527(v_13805);
  assign v_24528 = mux_24528(v_13811);
  assign v_24529 = mux_24529(v_13770);
  assign v_24531 = v_24532 | v_24534;
  assign v_24532 = mux_24532(v_24533);
  assign v_24533 = ~act_13354;
  assign v_24534 = v_24535 | v_24585;
  assign v_24535 = mux_24535(v_13355);
  assign v_24537 = v_24538 | v_24540;
  assign v_24538 = mux_24538(v_24539);
  assign v_24539 = ~act_13566;
  assign v_24540 = v_24541 | v_24563;
  assign v_24541 = mux_24541(v_13567);
  assign v_24543 = v_24544 | v_24546;
  assign v_24544 = mux_24544(v_24545);
  assign v_24545 = ~act_13666;
  assign v_24546 = v_24547 | v_24555;
  assign v_24547 = mux_24547(v_13667);
  assign v_24549 = v_24550 | v_24552;
  assign v_24550 = mux_24550(v_24551);
  assign v_24551 = ~act_13710;
  assign v_24552 = v_24553 | v_24554;
  assign v_24553 = mux_24553(v_13711);
  assign v_24554 = mux_24554(v_13717);
  assign v_24555 = mux_24555(v_13697);
  assign v_24557 = v_24558 | v_24560;
  assign v_24558 = mux_24558(v_24559);
  assign v_24559 = ~act_13673;
  assign v_24560 = v_24561 | v_24562;
  assign v_24561 = mux_24561(v_13674);
  assign v_24562 = mux_24562(v_13680);
  assign v_24563 = mux_24563(v_13653);
  assign v_24565 = v_24566 | v_24568;
  assign v_24566 = mux_24566(v_24567);
  assign v_24567 = ~act_13573;
  assign v_24568 = v_24569 | v_24577;
  assign v_24569 = mux_24569(v_13574);
  assign v_24571 = v_24572 | v_24574;
  assign v_24572 = mux_24572(v_24573);
  assign v_24573 = ~act_13617;
  assign v_24574 = v_24575 | v_24576;
  assign v_24575 = mux_24575(v_13618);
  assign v_24576 = mux_24576(v_13624);
  assign v_24577 = mux_24577(v_13604);
  assign v_24579 = v_24580 | v_24582;
  assign v_24580 = mux_24580(v_24581);
  assign v_24581 = ~act_13580;
  assign v_24582 = v_24583 | v_24584;
  assign v_24583 = mux_24583(v_13581);
  assign v_24584 = mux_24584(v_13587);
  assign v_24585 = mux_24585(v_13553);
  assign v_24587 = v_24588 | v_24590;
  assign v_24588 = mux_24588(v_24589);
  assign v_24589 = ~act_13361;
  assign v_24590 = v_24591 | v_24613;
  assign v_24591 = mux_24591(v_13362);
  assign v_24593 = v_24594 | v_24596;
  assign v_24594 = mux_24594(v_24595);
  assign v_24595 = ~act_13461;
  assign v_24596 = v_24597 | v_24605;
  assign v_24597 = mux_24597(v_13462);
  assign v_24599 = v_24600 | v_24602;
  assign v_24600 = mux_24600(v_24601);
  assign v_24601 = ~act_13505;
  assign v_24602 = v_24603 | v_24604;
  assign v_24603 = mux_24603(v_13506);
  assign v_24604 = mux_24604(v_13512);
  assign v_24605 = mux_24605(v_13492);
  assign v_24607 = v_24608 | v_24610;
  assign v_24608 = mux_24608(v_24609);
  assign v_24609 = ~act_13468;
  assign v_24610 = v_24611 | v_24612;
  assign v_24611 = mux_24611(v_13469);
  assign v_24612 = mux_24612(v_13475);
  assign v_24613 = mux_24613(v_13448);
  assign v_24615 = v_24616 | v_24618;
  assign v_24616 = mux_24616(v_24617);
  assign v_24617 = ~act_13368;
  assign v_24618 = v_24619 | v_24627;
  assign v_24619 = mux_24619(v_13369);
  assign v_24621 = v_24622 | v_24624;
  assign v_24622 = mux_24622(v_24623);
  assign v_24623 = ~act_13412;
  assign v_24624 = v_24625 | v_24626;
  assign v_24625 = mux_24625(v_13413);
  assign v_24626 = mux_24626(v_13419);
  assign v_24627 = mux_24627(v_13399);
  assign v_24629 = v_24630 | v_24632;
  assign v_24630 = mux_24630(v_24631);
  assign v_24631 = ~act_13375;
  assign v_24632 = v_24633 | v_24634;
  assign v_24633 = mux_24633(v_13376);
  assign v_24634 = mux_24634(v_13382);
  assign v_24635 = mux_24635(v_13327);
  assign v_24637 = v_24638 | v_24640;
  assign v_24638 = mux_24638(v_24639);
  assign v_24639 = ~act_11567;
  assign v_24640 = v_24641 | v_24859;
  assign v_24641 = mux_24641(v_11568);
  assign v_24643 = v_24644 | v_24646;
  assign v_24644 = mux_24644(v_24645);
  assign v_24645 = ~act_12451;
  assign v_24646 = v_24647 | v_24753;
  assign v_24647 = mux_24647(v_12452);
  assign v_24649 = v_24650 | v_24652;
  assign v_24650 = mux_24650(v_24651);
  assign v_24651 = ~act_12887;
  assign v_24652 = v_24653 | v_24703;
  assign v_24653 = mux_24653(v_12888);
  assign v_24655 = v_24656 | v_24658;
  assign v_24656 = mux_24656(v_24657);
  assign v_24657 = ~act_13099;
  assign v_24658 = v_24659 | v_24681;
  assign v_24659 = mux_24659(v_13100);
  assign v_24661 = v_24662 | v_24664;
  assign v_24662 = mux_24662(v_24663);
  assign v_24663 = ~act_13199;
  assign v_24664 = v_24665 | v_24673;
  assign v_24665 = mux_24665(v_13200);
  assign v_24667 = v_24668 | v_24670;
  assign v_24668 = mux_24668(v_24669);
  assign v_24669 = ~act_13243;
  assign v_24670 = v_24671 | v_24672;
  assign v_24671 = mux_24671(v_13244);
  assign v_24672 = mux_24672(v_13250);
  assign v_24673 = mux_24673(v_13230);
  assign v_24675 = v_24676 | v_24678;
  assign v_24676 = mux_24676(v_24677);
  assign v_24677 = ~act_13206;
  assign v_24678 = v_24679 | v_24680;
  assign v_24679 = mux_24679(v_13207);
  assign v_24680 = mux_24680(v_13213);
  assign v_24681 = mux_24681(v_13186);
  assign v_24683 = v_24684 | v_24686;
  assign v_24684 = mux_24684(v_24685);
  assign v_24685 = ~act_13106;
  assign v_24686 = v_24687 | v_24695;
  assign v_24687 = mux_24687(v_13107);
  assign v_24689 = v_24690 | v_24692;
  assign v_24690 = mux_24690(v_24691);
  assign v_24691 = ~act_13150;
  assign v_24692 = v_24693 | v_24694;
  assign v_24693 = mux_24693(v_13151);
  assign v_24694 = mux_24694(v_13157);
  assign v_24695 = mux_24695(v_13137);
  assign v_24697 = v_24698 | v_24700;
  assign v_24698 = mux_24698(v_24699);
  assign v_24699 = ~act_13113;
  assign v_24700 = v_24701 | v_24702;
  assign v_24701 = mux_24701(v_13114);
  assign v_24702 = mux_24702(v_13120);
  assign v_24703 = mux_24703(v_13086);
  assign v_24705 = v_24706 | v_24708;
  assign v_24706 = mux_24706(v_24707);
  assign v_24707 = ~act_12894;
  assign v_24708 = v_24709 | v_24731;
  assign v_24709 = mux_24709(v_12895);
  assign v_24711 = v_24712 | v_24714;
  assign v_24712 = mux_24712(v_24713);
  assign v_24713 = ~act_12994;
  assign v_24714 = v_24715 | v_24723;
  assign v_24715 = mux_24715(v_12995);
  assign v_24717 = v_24718 | v_24720;
  assign v_24718 = mux_24718(v_24719);
  assign v_24719 = ~act_13038;
  assign v_24720 = v_24721 | v_24722;
  assign v_24721 = mux_24721(v_13039);
  assign v_24722 = mux_24722(v_13045);
  assign v_24723 = mux_24723(v_13025);
  assign v_24725 = v_24726 | v_24728;
  assign v_24726 = mux_24726(v_24727);
  assign v_24727 = ~act_13001;
  assign v_24728 = v_24729 | v_24730;
  assign v_24729 = mux_24729(v_13002);
  assign v_24730 = mux_24730(v_13008);
  assign v_24731 = mux_24731(v_12981);
  assign v_24733 = v_24734 | v_24736;
  assign v_24734 = mux_24734(v_24735);
  assign v_24735 = ~act_12901;
  assign v_24736 = v_24737 | v_24745;
  assign v_24737 = mux_24737(v_12902);
  assign v_24739 = v_24740 | v_24742;
  assign v_24740 = mux_24740(v_24741);
  assign v_24741 = ~act_12945;
  assign v_24742 = v_24743 | v_24744;
  assign v_24743 = mux_24743(v_12946);
  assign v_24744 = mux_24744(v_12952);
  assign v_24745 = mux_24745(v_12932);
  assign v_24747 = v_24748 | v_24750;
  assign v_24748 = mux_24748(v_24749);
  assign v_24749 = ~act_12908;
  assign v_24750 = v_24751 | v_24752;
  assign v_24751 = mux_24751(v_12909);
  assign v_24752 = mux_24752(v_12915);
  assign v_24753 = mux_24753(v_12874);
  assign v_24755 = v_24756 | v_24758;
  assign v_24756 = mux_24756(v_24757);
  assign v_24757 = ~act_12458;
  assign v_24758 = v_24759 | v_24809;
  assign v_24759 = mux_24759(v_12459);
  assign v_24761 = v_24762 | v_24764;
  assign v_24762 = mux_24762(v_24763);
  assign v_24763 = ~act_12670;
  assign v_24764 = v_24765 | v_24787;
  assign v_24765 = mux_24765(v_12671);
  assign v_24767 = v_24768 | v_24770;
  assign v_24768 = mux_24768(v_24769);
  assign v_24769 = ~act_12770;
  assign v_24770 = v_24771 | v_24779;
  assign v_24771 = mux_24771(v_12771);
  assign v_24773 = v_24774 | v_24776;
  assign v_24774 = mux_24774(v_24775);
  assign v_24775 = ~act_12814;
  assign v_24776 = v_24777 | v_24778;
  assign v_24777 = mux_24777(v_12815);
  assign v_24778 = mux_24778(v_12821);
  assign v_24779 = mux_24779(v_12801);
  assign v_24781 = v_24782 | v_24784;
  assign v_24782 = mux_24782(v_24783);
  assign v_24783 = ~act_12777;
  assign v_24784 = v_24785 | v_24786;
  assign v_24785 = mux_24785(v_12778);
  assign v_24786 = mux_24786(v_12784);
  assign v_24787 = mux_24787(v_12757);
  assign v_24789 = v_24790 | v_24792;
  assign v_24790 = mux_24790(v_24791);
  assign v_24791 = ~act_12677;
  assign v_24792 = v_24793 | v_24801;
  assign v_24793 = mux_24793(v_12678);
  assign v_24795 = v_24796 | v_24798;
  assign v_24796 = mux_24796(v_24797);
  assign v_24797 = ~act_12721;
  assign v_24798 = v_24799 | v_24800;
  assign v_24799 = mux_24799(v_12722);
  assign v_24800 = mux_24800(v_12728);
  assign v_24801 = mux_24801(v_12708);
  assign v_24803 = v_24804 | v_24806;
  assign v_24804 = mux_24804(v_24805);
  assign v_24805 = ~act_12684;
  assign v_24806 = v_24807 | v_24808;
  assign v_24807 = mux_24807(v_12685);
  assign v_24808 = mux_24808(v_12691);
  assign v_24809 = mux_24809(v_12657);
  assign v_24811 = v_24812 | v_24814;
  assign v_24812 = mux_24812(v_24813);
  assign v_24813 = ~act_12465;
  assign v_24814 = v_24815 | v_24837;
  assign v_24815 = mux_24815(v_12466);
  assign v_24817 = v_24818 | v_24820;
  assign v_24818 = mux_24818(v_24819);
  assign v_24819 = ~act_12565;
  assign v_24820 = v_24821 | v_24829;
  assign v_24821 = mux_24821(v_12566);
  assign v_24823 = v_24824 | v_24826;
  assign v_24824 = mux_24824(v_24825);
  assign v_24825 = ~act_12609;
  assign v_24826 = v_24827 | v_24828;
  assign v_24827 = mux_24827(v_12610);
  assign v_24828 = mux_24828(v_12616);
  assign v_24829 = mux_24829(v_12596);
  assign v_24831 = v_24832 | v_24834;
  assign v_24832 = mux_24832(v_24833);
  assign v_24833 = ~act_12572;
  assign v_24834 = v_24835 | v_24836;
  assign v_24835 = mux_24835(v_12573);
  assign v_24836 = mux_24836(v_12579);
  assign v_24837 = mux_24837(v_12552);
  assign v_24839 = v_24840 | v_24842;
  assign v_24840 = mux_24840(v_24841);
  assign v_24841 = ~act_12472;
  assign v_24842 = v_24843 | v_24851;
  assign v_24843 = mux_24843(v_12473);
  assign v_24845 = v_24846 | v_24848;
  assign v_24846 = mux_24846(v_24847);
  assign v_24847 = ~act_12516;
  assign v_24848 = v_24849 | v_24850;
  assign v_24849 = mux_24849(v_12517);
  assign v_24850 = mux_24850(v_12523);
  assign v_24851 = mux_24851(v_12503);
  assign v_24853 = v_24854 | v_24856;
  assign v_24854 = mux_24854(v_24855);
  assign v_24855 = ~act_12479;
  assign v_24856 = v_24857 | v_24858;
  assign v_24857 = mux_24857(v_12480);
  assign v_24858 = mux_24858(v_12486);
  assign v_24859 = mux_24859(v_12438);
  assign v_24861 = v_24862 | v_24864;
  assign v_24862 = mux_24862(v_24863);
  assign v_24863 = ~act_11574;
  assign v_24864 = v_24865 | v_24971;
  assign v_24865 = mux_24865(v_11575);
  assign v_24867 = v_24868 | v_24870;
  assign v_24868 = mux_24868(v_24869);
  assign v_24869 = ~act_12010;
  assign v_24870 = v_24871 | v_24921;
  assign v_24871 = mux_24871(v_12011);
  assign v_24873 = v_24874 | v_24876;
  assign v_24874 = mux_24874(v_24875);
  assign v_24875 = ~act_12222;
  assign v_24876 = v_24877 | v_24899;
  assign v_24877 = mux_24877(v_12223);
  assign v_24879 = v_24880 | v_24882;
  assign v_24880 = mux_24880(v_24881);
  assign v_24881 = ~act_12322;
  assign v_24882 = v_24883 | v_24891;
  assign v_24883 = mux_24883(v_12323);
  assign v_24885 = v_24886 | v_24888;
  assign v_24886 = mux_24886(v_24887);
  assign v_24887 = ~act_12366;
  assign v_24888 = v_24889 | v_24890;
  assign v_24889 = mux_24889(v_12367);
  assign v_24890 = mux_24890(v_12373);
  assign v_24891 = mux_24891(v_12353);
  assign v_24893 = v_24894 | v_24896;
  assign v_24894 = mux_24894(v_24895);
  assign v_24895 = ~act_12329;
  assign v_24896 = v_24897 | v_24898;
  assign v_24897 = mux_24897(v_12330);
  assign v_24898 = mux_24898(v_12336);
  assign v_24899 = mux_24899(v_12309);
  assign v_24901 = v_24902 | v_24904;
  assign v_24902 = mux_24902(v_24903);
  assign v_24903 = ~act_12229;
  assign v_24904 = v_24905 | v_24913;
  assign v_24905 = mux_24905(v_12230);
  assign v_24907 = v_24908 | v_24910;
  assign v_24908 = mux_24908(v_24909);
  assign v_24909 = ~act_12273;
  assign v_24910 = v_24911 | v_24912;
  assign v_24911 = mux_24911(v_12274);
  assign v_24912 = mux_24912(v_12280);
  assign v_24913 = mux_24913(v_12260);
  assign v_24915 = v_24916 | v_24918;
  assign v_24916 = mux_24916(v_24917);
  assign v_24917 = ~act_12236;
  assign v_24918 = v_24919 | v_24920;
  assign v_24919 = mux_24919(v_12237);
  assign v_24920 = mux_24920(v_12243);
  assign v_24921 = mux_24921(v_12209);
  assign v_24923 = v_24924 | v_24926;
  assign v_24924 = mux_24924(v_24925);
  assign v_24925 = ~act_12017;
  assign v_24926 = v_24927 | v_24949;
  assign v_24927 = mux_24927(v_12018);
  assign v_24929 = v_24930 | v_24932;
  assign v_24930 = mux_24930(v_24931);
  assign v_24931 = ~act_12117;
  assign v_24932 = v_24933 | v_24941;
  assign v_24933 = mux_24933(v_12118);
  assign v_24935 = v_24936 | v_24938;
  assign v_24936 = mux_24936(v_24937);
  assign v_24937 = ~act_12161;
  assign v_24938 = v_24939 | v_24940;
  assign v_24939 = mux_24939(v_12162);
  assign v_24940 = mux_24940(v_12168);
  assign v_24941 = mux_24941(v_12148);
  assign v_24943 = v_24944 | v_24946;
  assign v_24944 = mux_24944(v_24945);
  assign v_24945 = ~act_12124;
  assign v_24946 = v_24947 | v_24948;
  assign v_24947 = mux_24947(v_12125);
  assign v_24948 = mux_24948(v_12131);
  assign v_24949 = mux_24949(v_12104);
  assign v_24951 = v_24952 | v_24954;
  assign v_24952 = mux_24952(v_24953);
  assign v_24953 = ~act_12024;
  assign v_24954 = v_24955 | v_24963;
  assign v_24955 = mux_24955(v_12025);
  assign v_24957 = v_24958 | v_24960;
  assign v_24958 = mux_24958(v_24959);
  assign v_24959 = ~act_12068;
  assign v_24960 = v_24961 | v_24962;
  assign v_24961 = mux_24961(v_12069);
  assign v_24962 = mux_24962(v_12075);
  assign v_24963 = mux_24963(v_12055);
  assign v_24965 = v_24966 | v_24968;
  assign v_24966 = mux_24966(v_24967);
  assign v_24967 = ~act_12031;
  assign v_24968 = v_24969 | v_24970;
  assign v_24969 = mux_24969(v_12032);
  assign v_24970 = mux_24970(v_12038);
  assign v_24971 = mux_24971(v_11997);
  assign v_24973 = v_24974 | v_24976;
  assign v_24974 = mux_24974(v_24975);
  assign v_24975 = ~act_11581;
  assign v_24976 = v_24977 | v_25027;
  assign v_24977 = mux_24977(v_11582);
  assign v_24979 = v_24980 | v_24982;
  assign v_24980 = mux_24980(v_24981);
  assign v_24981 = ~act_11793;
  assign v_24982 = v_24983 | v_25005;
  assign v_24983 = mux_24983(v_11794);
  assign v_24985 = v_24986 | v_24988;
  assign v_24986 = mux_24986(v_24987);
  assign v_24987 = ~act_11893;
  assign v_24988 = v_24989 | v_24997;
  assign v_24989 = mux_24989(v_11894);
  assign v_24991 = v_24992 | v_24994;
  assign v_24992 = mux_24992(v_24993);
  assign v_24993 = ~act_11937;
  assign v_24994 = v_24995 | v_24996;
  assign v_24995 = mux_24995(v_11938);
  assign v_24996 = mux_24996(v_11944);
  assign v_24997 = mux_24997(v_11924);
  assign v_24999 = v_25000 | v_25002;
  assign v_25000 = mux_25000(v_25001);
  assign v_25001 = ~act_11900;
  assign v_25002 = v_25003 | v_25004;
  assign v_25003 = mux_25003(v_11901);
  assign v_25004 = mux_25004(v_11907);
  assign v_25005 = mux_25005(v_11880);
  assign v_25007 = v_25008 | v_25010;
  assign v_25008 = mux_25008(v_25009);
  assign v_25009 = ~act_11800;
  assign v_25010 = v_25011 | v_25019;
  assign v_25011 = mux_25011(v_11801);
  assign v_25013 = v_25014 | v_25016;
  assign v_25014 = mux_25014(v_25015);
  assign v_25015 = ~act_11844;
  assign v_25016 = v_25017 | v_25018;
  assign v_25017 = mux_25017(v_11845);
  assign v_25018 = mux_25018(v_11851);
  assign v_25019 = mux_25019(v_11831);
  assign v_25021 = v_25022 | v_25024;
  assign v_25022 = mux_25022(v_25023);
  assign v_25023 = ~act_11807;
  assign v_25024 = v_25025 | v_25026;
  assign v_25025 = mux_25025(v_11808);
  assign v_25026 = mux_25026(v_11814);
  assign v_25027 = mux_25027(v_11780);
  assign v_25029 = v_25030 | v_25032;
  assign v_25030 = mux_25030(v_25031);
  assign v_25031 = ~act_11588;
  assign v_25032 = v_25033 | v_25055;
  assign v_25033 = mux_25033(v_11589);
  assign v_25035 = v_25036 | v_25038;
  assign v_25036 = mux_25036(v_25037);
  assign v_25037 = ~act_11688;
  assign v_25038 = v_25039 | v_25047;
  assign v_25039 = mux_25039(v_11689);
  assign v_25041 = v_25042 | v_25044;
  assign v_25042 = mux_25042(v_25043);
  assign v_25043 = ~act_11732;
  assign v_25044 = v_25045 | v_25046;
  assign v_25045 = mux_25045(v_11733);
  assign v_25046 = mux_25046(v_11739);
  assign v_25047 = mux_25047(v_11719);
  assign v_25049 = v_25050 | v_25052;
  assign v_25050 = mux_25050(v_25051);
  assign v_25051 = ~act_11695;
  assign v_25052 = v_25053 | v_25054;
  assign v_25053 = mux_25053(v_11696);
  assign v_25054 = mux_25054(v_11702);
  assign v_25055 = mux_25055(v_11675);
  assign v_25057 = v_25058 | v_25060;
  assign v_25058 = mux_25058(v_25059);
  assign v_25059 = ~act_11595;
  assign v_25060 = v_25061 | v_25069;
  assign v_25061 = mux_25061(v_11596);
  assign v_25063 = v_25064 | v_25066;
  assign v_25064 = mux_25064(v_25065);
  assign v_25065 = ~act_11639;
  assign v_25066 = v_25067 | v_25068;
  assign v_25067 = mux_25067(v_11640);
  assign v_25068 = mux_25068(v_11646);
  assign v_25069 = mux_25069(v_11626);
  assign v_25071 = v_25072 | v_25074;
  assign v_25072 = mux_25072(v_25073);
  assign v_25073 = ~act_11602;
  assign v_25074 = v_25075 | v_25076;
  assign v_25075 = mux_25075(v_11603);
  assign v_25076 = mux_25076(v_11609);
  assign v_25077 = mux_25077(v_11547);
  assign v_25079 = v_25080 | v_25082;
  assign v_25080 = mux_25080(v_25081);
  assign v_25081 = ~act_7995;
  assign v_25082 = v_25083 | v_25525;
  assign v_25083 = mux_25083(v_7996);
  assign v_25085 = v_25086 | v_25088;
  assign v_25086 = mux_25086(v_25087);
  assign v_25087 = ~act_9775;
  assign v_25088 = v_25089 | v_25307;
  assign v_25089 = mux_25089(v_9776);
  assign v_25091 = v_25092 | v_25094;
  assign v_25092 = mux_25092(v_25093);
  assign v_25093 = ~act_10659;
  assign v_25094 = v_25095 | v_25201;
  assign v_25095 = mux_25095(v_10660);
  assign v_25097 = v_25098 | v_25100;
  assign v_25098 = mux_25098(v_25099);
  assign v_25099 = ~act_11095;
  assign v_25100 = v_25101 | v_25151;
  assign v_25101 = mux_25101(v_11096);
  assign v_25103 = v_25104 | v_25106;
  assign v_25104 = mux_25104(v_25105);
  assign v_25105 = ~act_11307;
  assign v_25106 = v_25107 | v_25129;
  assign v_25107 = mux_25107(v_11308);
  assign v_25109 = v_25110 | v_25112;
  assign v_25110 = mux_25110(v_25111);
  assign v_25111 = ~act_11407;
  assign v_25112 = v_25113 | v_25121;
  assign v_25113 = mux_25113(v_11408);
  assign v_25115 = v_25116 | v_25118;
  assign v_25116 = mux_25116(v_25117);
  assign v_25117 = ~act_11451;
  assign v_25118 = v_25119 | v_25120;
  assign v_25119 = mux_25119(v_11452);
  assign v_25120 = mux_25120(v_11458);
  assign v_25121 = mux_25121(v_11438);
  assign v_25123 = v_25124 | v_25126;
  assign v_25124 = mux_25124(v_25125);
  assign v_25125 = ~act_11414;
  assign v_25126 = v_25127 | v_25128;
  assign v_25127 = mux_25127(v_11415);
  assign v_25128 = mux_25128(v_11421);
  assign v_25129 = mux_25129(v_11394);
  assign v_25131 = v_25132 | v_25134;
  assign v_25132 = mux_25132(v_25133);
  assign v_25133 = ~act_11314;
  assign v_25134 = v_25135 | v_25143;
  assign v_25135 = mux_25135(v_11315);
  assign v_25137 = v_25138 | v_25140;
  assign v_25138 = mux_25138(v_25139);
  assign v_25139 = ~act_11358;
  assign v_25140 = v_25141 | v_25142;
  assign v_25141 = mux_25141(v_11359);
  assign v_25142 = mux_25142(v_11365);
  assign v_25143 = mux_25143(v_11345);
  assign v_25145 = v_25146 | v_25148;
  assign v_25146 = mux_25146(v_25147);
  assign v_25147 = ~act_11321;
  assign v_25148 = v_25149 | v_25150;
  assign v_25149 = mux_25149(v_11322);
  assign v_25150 = mux_25150(v_11328);
  assign v_25151 = mux_25151(v_11294);
  assign v_25153 = v_25154 | v_25156;
  assign v_25154 = mux_25154(v_25155);
  assign v_25155 = ~act_11102;
  assign v_25156 = v_25157 | v_25179;
  assign v_25157 = mux_25157(v_11103);
  assign v_25159 = v_25160 | v_25162;
  assign v_25160 = mux_25160(v_25161);
  assign v_25161 = ~act_11202;
  assign v_25162 = v_25163 | v_25171;
  assign v_25163 = mux_25163(v_11203);
  assign v_25165 = v_25166 | v_25168;
  assign v_25166 = mux_25166(v_25167);
  assign v_25167 = ~act_11246;
  assign v_25168 = v_25169 | v_25170;
  assign v_25169 = mux_25169(v_11247);
  assign v_25170 = mux_25170(v_11253);
  assign v_25171 = mux_25171(v_11233);
  assign v_25173 = v_25174 | v_25176;
  assign v_25174 = mux_25174(v_25175);
  assign v_25175 = ~act_11209;
  assign v_25176 = v_25177 | v_25178;
  assign v_25177 = mux_25177(v_11210);
  assign v_25178 = mux_25178(v_11216);
  assign v_25179 = mux_25179(v_11189);
  assign v_25181 = v_25182 | v_25184;
  assign v_25182 = mux_25182(v_25183);
  assign v_25183 = ~act_11109;
  assign v_25184 = v_25185 | v_25193;
  assign v_25185 = mux_25185(v_11110);
  assign v_25187 = v_25188 | v_25190;
  assign v_25188 = mux_25188(v_25189);
  assign v_25189 = ~act_11153;
  assign v_25190 = v_25191 | v_25192;
  assign v_25191 = mux_25191(v_11154);
  assign v_25192 = mux_25192(v_11160);
  assign v_25193 = mux_25193(v_11140);
  assign v_25195 = v_25196 | v_25198;
  assign v_25196 = mux_25196(v_25197);
  assign v_25197 = ~act_11116;
  assign v_25198 = v_25199 | v_25200;
  assign v_25199 = mux_25199(v_11117);
  assign v_25200 = mux_25200(v_11123);
  assign v_25201 = mux_25201(v_11082);
  assign v_25203 = v_25204 | v_25206;
  assign v_25204 = mux_25204(v_25205);
  assign v_25205 = ~act_10666;
  assign v_25206 = v_25207 | v_25257;
  assign v_25207 = mux_25207(v_10667);
  assign v_25209 = v_25210 | v_25212;
  assign v_25210 = mux_25210(v_25211);
  assign v_25211 = ~act_10878;
  assign v_25212 = v_25213 | v_25235;
  assign v_25213 = mux_25213(v_10879);
  assign v_25215 = v_25216 | v_25218;
  assign v_25216 = mux_25216(v_25217);
  assign v_25217 = ~act_10978;
  assign v_25218 = v_25219 | v_25227;
  assign v_25219 = mux_25219(v_10979);
  assign v_25221 = v_25222 | v_25224;
  assign v_25222 = mux_25222(v_25223);
  assign v_25223 = ~act_11022;
  assign v_25224 = v_25225 | v_25226;
  assign v_25225 = mux_25225(v_11023);
  assign v_25226 = mux_25226(v_11029);
  assign v_25227 = mux_25227(v_11009);
  assign v_25229 = v_25230 | v_25232;
  assign v_25230 = mux_25230(v_25231);
  assign v_25231 = ~act_10985;
  assign v_25232 = v_25233 | v_25234;
  assign v_25233 = mux_25233(v_10986);
  assign v_25234 = mux_25234(v_10992);
  assign v_25235 = mux_25235(v_10965);
  assign v_25237 = v_25238 | v_25240;
  assign v_25238 = mux_25238(v_25239);
  assign v_25239 = ~act_10885;
  assign v_25240 = v_25241 | v_25249;
  assign v_25241 = mux_25241(v_10886);
  assign v_25243 = v_25244 | v_25246;
  assign v_25244 = mux_25244(v_25245);
  assign v_25245 = ~act_10929;
  assign v_25246 = v_25247 | v_25248;
  assign v_25247 = mux_25247(v_10930);
  assign v_25248 = mux_25248(v_10936);
  assign v_25249 = mux_25249(v_10916);
  assign v_25251 = v_25252 | v_25254;
  assign v_25252 = mux_25252(v_25253);
  assign v_25253 = ~act_10892;
  assign v_25254 = v_25255 | v_25256;
  assign v_25255 = mux_25255(v_10893);
  assign v_25256 = mux_25256(v_10899);
  assign v_25257 = mux_25257(v_10865);
  assign v_25259 = v_25260 | v_25262;
  assign v_25260 = mux_25260(v_25261);
  assign v_25261 = ~act_10673;
  assign v_25262 = v_25263 | v_25285;
  assign v_25263 = mux_25263(v_10674);
  assign v_25265 = v_25266 | v_25268;
  assign v_25266 = mux_25266(v_25267);
  assign v_25267 = ~act_10773;
  assign v_25268 = v_25269 | v_25277;
  assign v_25269 = mux_25269(v_10774);
  assign v_25271 = v_25272 | v_25274;
  assign v_25272 = mux_25272(v_25273);
  assign v_25273 = ~act_10817;
  assign v_25274 = v_25275 | v_25276;
  assign v_25275 = mux_25275(v_10818);
  assign v_25276 = mux_25276(v_10824);
  assign v_25277 = mux_25277(v_10804);
  assign v_25279 = v_25280 | v_25282;
  assign v_25280 = mux_25280(v_25281);
  assign v_25281 = ~act_10780;
  assign v_25282 = v_25283 | v_25284;
  assign v_25283 = mux_25283(v_10781);
  assign v_25284 = mux_25284(v_10787);
  assign v_25285 = mux_25285(v_10760);
  assign v_25287 = v_25288 | v_25290;
  assign v_25288 = mux_25288(v_25289);
  assign v_25289 = ~act_10680;
  assign v_25290 = v_25291 | v_25299;
  assign v_25291 = mux_25291(v_10681);
  assign v_25293 = v_25294 | v_25296;
  assign v_25294 = mux_25294(v_25295);
  assign v_25295 = ~act_10724;
  assign v_25296 = v_25297 | v_25298;
  assign v_25297 = mux_25297(v_10725);
  assign v_25298 = mux_25298(v_10731);
  assign v_25299 = mux_25299(v_10711);
  assign v_25301 = v_25302 | v_25304;
  assign v_25302 = mux_25302(v_25303);
  assign v_25303 = ~act_10687;
  assign v_25304 = v_25305 | v_25306;
  assign v_25305 = mux_25305(v_10688);
  assign v_25306 = mux_25306(v_10694);
  assign v_25307 = mux_25307(v_10646);
  assign v_25309 = v_25310 | v_25312;
  assign v_25310 = mux_25310(v_25311);
  assign v_25311 = ~act_9782;
  assign v_25312 = v_25313 | v_25419;
  assign v_25313 = mux_25313(v_9783);
  assign v_25315 = v_25316 | v_25318;
  assign v_25316 = mux_25316(v_25317);
  assign v_25317 = ~act_10218;
  assign v_25318 = v_25319 | v_25369;
  assign v_25319 = mux_25319(v_10219);
  assign v_25321 = v_25322 | v_25324;
  assign v_25322 = mux_25322(v_25323);
  assign v_25323 = ~act_10430;
  assign v_25324 = v_25325 | v_25347;
  assign v_25325 = mux_25325(v_10431);
  assign v_25327 = v_25328 | v_25330;
  assign v_25328 = mux_25328(v_25329);
  assign v_25329 = ~act_10530;
  assign v_25330 = v_25331 | v_25339;
  assign v_25331 = mux_25331(v_10531);
  assign v_25333 = v_25334 | v_25336;
  assign v_25334 = mux_25334(v_25335);
  assign v_25335 = ~act_10574;
  assign v_25336 = v_25337 | v_25338;
  assign v_25337 = mux_25337(v_10575);
  assign v_25338 = mux_25338(v_10581);
  assign v_25339 = mux_25339(v_10561);
  assign v_25341 = v_25342 | v_25344;
  assign v_25342 = mux_25342(v_25343);
  assign v_25343 = ~act_10537;
  assign v_25344 = v_25345 | v_25346;
  assign v_25345 = mux_25345(v_10538);
  assign v_25346 = mux_25346(v_10544);
  assign v_25347 = mux_25347(v_10517);
  assign v_25349 = v_25350 | v_25352;
  assign v_25350 = mux_25350(v_25351);
  assign v_25351 = ~act_10437;
  assign v_25352 = v_25353 | v_25361;
  assign v_25353 = mux_25353(v_10438);
  assign v_25355 = v_25356 | v_25358;
  assign v_25356 = mux_25356(v_25357);
  assign v_25357 = ~act_10481;
  assign v_25358 = v_25359 | v_25360;
  assign v_25359 = mux_25359(v_10482);
  assign v_25360 = mux_25360(v_10488);
  assign v_25361 = mux_25361(v_10468);
  assign v_25363 = v_25364 | v_25366;
  assign v_25364 = mux_25364(v_25365);
  assign v_25365 = ~act_10444;
  assign v_25366 = v_25367 | v_25368;
  assign v_25367 = mux_25367(v_10445);
  assign v_25368 = mux_25368(v_10451);
  assign v_25369 = mux_25369(v_10417);
  assign v_25371 = v_25372 | v_25374;
  assign v_25372 = mux_25372(v_25373);
  assign v_25373 = ~act_10225;
  assign v_25374 = v_25375 | v_25397;
  assign v_25375 = mux_25375(v_10226);
  assign v_25377 = v_25378 | v_25380;
  assign v_25378 = mux_25378(v_25379);
  assign v_25379 = ~act_10325;
  assign v_25380 = v_25381 | v_25389;
  assign v_25381 = mux_25381(v_10326);
  assign v_25383 = v_25384 | v_25386;
  assign v_25384 = mux_25384(v_25385);
  assign v_25385 = ~act_10369;
  assign v_25386 = v_25387 | v_25388;
  assign v_25387 = mux_25387(v_10370);
  assign v_25388 = mux_25388(v_10376);
  assign v_25389 = mux_25389(v_10356);
  assign v_25391 = v_25392 | v_25394;
  assign v_25392 = mux_25392(v_25393);
  assign v_25393 = ~act_10332;
  assign v_25394 = v_25395 | v_25396;
  assign v_25395 = mux_25395(v_10333);
  assign v_25396 = mux_25396(v_10339);
  assign v_25397 = mux_25397(v_10312);
  assign v_25399 = v_25400 | v_25402;
  assign v_25400 = mux_25400(v_25401);
  assign v_25401 = ~act_10232;
  assign v_25402 = v_25403 | v_25411;
  assign v_25403 = mux_25403(v_10233);
  assign v_25405 = v_25406 | v_25408;
  assign v_25406 = mux_25406(v_25407);
  assign v_25407 = ~act_10276;
  assign v_25408 = v_25409 | v_25410;
  assign v_25409 = mux_25409(v_10277);
  assign v_25410 = mux_25410(v_10283);
  assign v_25411 = mux_25411(v_10263);
  assign v_25413 = v_25414 | v_25416;
  assign v_25414 = mux_25414(v_25415);
  assign v_25415 = ~act_10239;
  assign v_25416 = v_25417 | v_25418;
  assign v_25417 = mux_25417(v_10240);
  assign v_25418 = mux_25418(v_10246);
  assign v_25419 = mux_25419(v_10205);
  assign v_25421 = v_25422 | v_25424;
  assign v_25422 = mux_25422(v_25423);
  assign v_25423 = ~act_9789;
  assign v_25424 = v_25425 | v_25475;
  assign v_25425 = mux_25425(v_9790);
  assign v_25427 = v_25428 | v_25430;
  assign v_25428 = mux_25428(v_25429);
  assign v_25429 = ~act_10001;
  assign v_25430 = v_25431 | v_25453;
  assign v_25431 = mux_25431(v_10002);
  assign v_25433 = v_25434 | v_25436;
  assign v_25434 = mux_25434(v_25435);
  assign v_25435 = ~act_10101;
  assign v_25436 = v_25437 | v_25445;
  assign v_25437 = mux_25437(v_10102);
  assign v_25439 = v_25440 | v_25442;
  assign v_25440 = mux_25440(v_25441);
  assign v_25441 = ~act_10145;
  assign v_25442 = v_25443 | v_25444;
  assign v_25443 = mux_25443(v_10146);
  assign v_25444 = mux_25444(v_10152);
  assign v_25445 = mux_25445(v_10132);
  assign v_25447 = v_25448 | v_25450;
  assign v_25448 = mux_25448(v_25449);
  assign v_25449 = ~act_10108;
  assign v_25450 = v_25451 | v_25452;
  assign v_25451 = mux_25451(v_10109);
  assign v_25452 = mux_25452(v_10115);
  assign v_25453 = mux_25453(v_10088);
  assign v_25455 = v_25456 | v_25458;
  assign v_25456 = mux_25456(v_25457);
  assign v_25457 = ~act_10008;
  assign v_25458 = v_25459 | v_25467;
  assign v_25459 = mux_25459(v_10009);
  assign v_25461 = v_25462 | v_25464;
  assign v_25462 = mux_25462(v_25463);
  assign v_25463 = ~act_10052;
  assign v_25464 = v_25465 | v_25466;
  assign v_25465 = mux_25465(v_10053);
  assign v_25466 = mux_25466(v_10059);
  assign v_25467 = mux_25467(v_10039);
  assign v_25469 = v_25470 | v_25472;
  assign v_25470 = mux_25470(v_25471);
  assign v_25471 = ~act_10015;
  assign v_25472 = v_25473 | v_25474;
  assign v_25473 = mux_25473(v_10016);
  assign v_25474 = mux_25474(v_10022);
  assign v_25475 = mux_25475(v_9988);
  assign v_25477 = v_25478 | v_25480;
  assign v_25478 = mux_25478(v_25479);
  assign v_25479 = ~act_9796;
  assign v_25480 = v_25481 | v_25503;
  assign v_25481 = mux_25481(v_9797);
  assign v_25483 = v_25484 | v_25486;
  assign v_25484 = mux_25484(v_25485);
  assign v_25485 = ~act_9896;
  assign v_25486 = v_25487 | v_25495;
  assign v_25487 = mux_25487(v_9897);
  assign v_25489 = v_25490 | v_25492;
  assign v_25490 = mux_25490(v_25491);
  assign v_25491 = ~act_9940;
  assign v_25492 = v_25493 | v_25494;
  assign v_25493 = mux_25493(v_9941);
  assign v_25494 = mux_25494(v_9947);
  assign v_25495 = mux_25495(v_9927);
  assign v_25497 = v_25498 | v_25500;
  assign v_25498 = mux_25498(v_25499);
  assign v_25499 = ~act_9903;
  assign v_25500 = v_25501 | v_25502;
  assign v_25501 = mux_25501(v_9904);
  assign v_25502 = mux_25502(v_9910);
  assign v_25503 = mux_25503(v_9883);
  assign v_25505 = v_25506 | v_25508;
  assign v_25506 = mux_25506(v_25507);
  assign v_25507 = ~act_9803;
  assign v_25508 = v_25509 | v_25517;
  assign v_25509 = mux_25509(v_9804);
  assign v_25511 = v_25512 | v_25514;
  assign v_25512 = mux_25512(v_25513);
  assign v_25513 = ~act_9847;
  assign v_25514 = v_25515 | v_25516;
  assign v_25515 = mux_25515(v_9848);
  assign v_25516 = mux_25516(v_9854);
  assign v_25517 = mux_25517(v_9834);
  assign v_25519 = v_25520 | v_25522;
  assign v_25520 = mux_25520(v_25521);
  assign v_25521 = ~act_9810;
  assign v_25522 = v_25523 | v_25524;
  assign v_25523 = mux_25523(v_9811);
  assign v_25524 = mux_25524(v_9817);
  assign v_25525 = mux_25525(v_9762);
  assign v_25527 = v_25528 | v_25530;
  assign v_25528 = mux_25528(v_25529);
  assign v_25529 = ~act_8002;
  assign v_25530 = v_25531 | v_25749;
  assign v_25531 = mux_25531(v_8003);
  assign v_25533 = v_25534 | v_25536;
  assign v_25534 = mux_25534(v_25535);
  assign v_25535 = ~act_8886;
  assign v_25536 = v_25537 | v_25643;
  assign v_25537 = mux_25537(v_8887);
  assign v_25539 = v_25540 | v_25542;
  assign v_25540 = mux_25540(v_25541);
  assign v_25541 = ~act_9322;
  assign v_25542 = v_25543 | v_25593;
  assign v_25543 = mux_25543(v_9323);
  assign v_25545 = v_25546 | v_25548;
  assign v_25546 = mux_25546(v_25547);
  assign v_25547 = ~act_9534;
  assign v_25548 = v_25549 | v_25571;
  assign v_25549 = mux_25549(v_9535);
  assign v_25551 = v_25552 | v_25554;
  assign v_25552 = mux_25552(v_25553);
  assign v_25553 = ~act_9634;
  assign v_25554 = v_25555 | v_25563;
  assign v_25555 = mux_25555(v_9635);
  assign v_25557 = v_25558 | v_25560;
  assign v_25558 = mux_25558(v_25559);
  assign v_25559 = ~act_9678;
  assign v_25560 = v_25561 | v_25562;
  assign v_25561 = mux_25561(v_9679);
  assign v_25562 = mux_25562(v_9685);
  assign v_25563 = mux_25563(v_9665);
  assign v_25565 = v_25566 | v_25568;
  assign v_25566 = mux_25566(v_25567);
  assign v_25567 = ~act_9641;
  assign v_25568 = v_25569 | v_25570;
  assign v_25569 = mux_25569(v_9642);
  assign v_25570 = mux_25570(v_9648);
  assign v_25571 = mux_25571(v_9621);
  assign v_25573 = v_25574 | v_25576;
  assign v_25574 = mux_25574(v_25575);
  assign v_25575 = ~act_9541;
  assign v_25576 = v_25577 | v_25585;
  assign v_25577 = mux_25577(v_9542);
  assign v_25579 = v_25580 | v_25582;
  assign v_25580 = mux_25580(v_25581);
  assign v_25581 = ~act_9585;
  assign v_25582 = v_25583 | v_25584;
  assign v_25583 = mux_25583(v_9586);
  assign v_25584 = mux_25584(v_9592);
  assign v_25585 = mux_25585(v_9572);
  assign v_25587 = v_25588 | v_25590;
  assign v_25588 = mux_25588(v_25589);
  assign v_25589 = ~act_9548;
  assign v_25590 = v_25591 | v_25592;
  assign v_25591 = mux_25591(v_9549);
  assign v_25592 = mux_25592(v_9555);
  assign v_25593 = mux_25593(v_9521);
  assign v_25595 = v_25596 | v_25598;
  assign v_25596 = mux_25596(v_25597);
  assign v_25597 = ~act_9329;
  assign v_25598 = v_25599 | v_25621;
  assign v_25599 = mux_25599(v_9330);
  assign v_25601 = v_25602 | v_25604;
  assign v_25602 = mux_25602(v_25603);
  assign v_25603 = ~act_9429;
  assign v_25604 = v_25605 | v_25613;
  assign v_25605 = mux_25605(v_9430);
  assign v_25607 = v_25608 | v_25610;
  assign v_25608 = mux_25608(v_25609);
  assign v_25609 = ~act_9473;
  assign v_25610 = v_25611 | v_25612;
  assign v_25611 = mux_25611(v_9474);
  assign v_25612 = mux_25612(v_9480);
  assign v_25613 = mux_25613(v_9460);
  assign v_25615 = v_25616 | v_25618;
  assign v_25616 = mux_25616(v_25617);
  assign v_25617 = ~act_9436;
  assign v_25618 = v_25619 | v_25620;
  assign v_25619 = mux_25619(v_9437);
  assign v_25620 = mux_25620(v_9443);
  assign v_25621 = mux_25621(v_9416);
  assign v_25623 = v_25624 | v_25626;
  assign v_25624 = mux_25624(v_25625);
  assign v_25625 = ~act_9336;
  assign v_25626 = v_25627 | v_25635;
  assign v_25627 = mux_25627(v_9337);
  assign v_25629 = v_25630 | v_25632;
  assign v_25630 = mux_25630(v_25631);
  assign v_25631 = ~act_9380;
  assign v_25632 = v_25633 | v_25634;
  assign v_25633 = mux_25633(v_9381);
  assign v_25634 = mux_25634(v_9387);
  assign v_25635 = mux_25635(v_9367);
  assign v_25637 = v_25638 | v_25640;
  assign v_25638 = mux_25638(v_25639);
  assign v_25639 = ~act_9343;
  assign v_25640 = v_25641 | v_25642;
  assign v_25641 = mux_25641(v_9344);
  assign v_25642 = mux_25642(v_9350);
  assign v_25643 = mux_25643(v_9309);
  assign v_25645 = v_25646 | v_25648;
  assign v_25646 = mux_25646(v_25647);
  assign v_25647 = ~act_8893;
  assign v_25648 = v_25649 | v_25699;
  assign v_25649 = mux_25649(v_8894);
  assign v_25651 = v_25652 | v_25654;
  assign v_25652 = mux_25652(v_25653);
  assign v_25653 = ~act_9105;
  assign v_25654 = v_25655 | v_25677;
  assign v_25655 = mux_25655(v_9106);
  assign v_25657 = v_25658 | v_25660;
  assign v_25658 = mux_25658(v_25659);
  assign v_25659 = ~act_9205;
  assign v_25660 = v_25661 | v_25669;
  assign v_25661 = mux_25661(v_9206);
  assign v_25663 = v_25664 | v_25666;
  assign v_25664 = mux_25664(v_25665);
  assign v_25665 = ~act_9249;
  assign v_25666 = v_25667 | v_25668;
  assign v_25667 = mux_25667(v_9250);
  assign v_25668 = mux_25668(v_9256);
  assign v_25669 = mux_25669(v_9236);
  assign v_25671 = v_25672 | v_25674;
  assign v_25672 = mux_25672(v_25673);
  assign v_25673 = ~act_9212;
  assign v_25674 = v_25675 | v_25676;
  assign v_25675 = mux_25675(v_9213);
  assign v_25676 = mux_25676(v_9219);
  assign v_25677 = mux_25677(v_9192);
  assign v_25679 = v_25680 | v_25682;
  assign v_25680 = mux_25680(v_25681);
  assign v_25681 = ~act_9112;
  assign v_25682 = v_25683 | v_25691;
  assign v_25683 = mux_25683(v_9113);
  assign v_25685 = v_25686 | v_25688;
  assign v_25686 = mux_25686(v_25687);
  assign v_25687 = ~act_9156;
  assign v_25688 = v_25689 | v_25690;
  assign v_25689 = mux_25689(v_9157);
  assign v_25690 = mux_25690(v_9163);
  assign v_25691 = mux_25691(v_9143);
  assign v_25693 = v_25694 | v_25696;
  assign v_25694 = mux_25694(v_25695);
  assign v_25695 = ~act_9119;
  assign v_25696 = v_25697 | v_25698;
  assign v_25697 = mux_25697(v_9120);
  assign v_25698 = mux_25698(v_9126);
  assign v_25699 = mux_25699(v_9092);
  assign v_25701 = v_25702 | v_25704;
  assign v_25702 = mux_25702(v_25703);
  assign v_25703 = ~act_8900;
  assign v_25704 = v_25705 | v_25727;
  assign v_25705 = mux_25705(v_8901);
  assign v_25707 = v_25708 | v_25710;
  assign v_25708 = mux_25708(v_25709);
  assign v_25709 = ~act_9000;
  assign v_25710 = v_25711 | v_25719;
  assign v_25711 = mux_25711(v_9001);
  assign v_25713 = v_25714 | v_25716;
  assign v_25714 = mux_25714(v_25715);
  assign v_25715 = ~act_9044;
  assign v_25716 = v_25717 | v_25718;
  assign v_25717 = mux_25717(v_9045);
  assign v_25718 = mux_25718(v_9051);
  assign v_25719 = mux_25719(v_9031);
  assign v_25721 = v_25722 | v_25724;
  assign v_25722 = mux_25722(v_25723);
  assign v_25723 = ~act_9007;
  assign v_25724 = v_25725 | v_25726;
  assign v_25725 = mux_25725(v_9008);
  assign v_25726 = mux_25726(v_9014);
  assign v_25727 = mux_25727(v_8987);
  assign v_25729 = v_25730 | v_25732;
  assign v_25730 = mux_25730(v_25731);
  assign v_25731 = ~act_8907;
  assign v_25732 = v_25733 | v_25741;
  assign v_25733 = mux_25733(v_8908);
  assign v_25735 = v_25736 | v_25738;
  assign v_25736 = mux_25736(v_25737);
  assign v_25737 = ~act_8951;
  assign v_25738 = v_25739 | v_25740;
  assign v_25739 = mux_25739(v_8952);
  assign v_25740 = mux_25740(v_8958);
  assign v_25741 = mux_25741(v_8938);
  assign v_25743 = v_25744 | v_25746;
  assign v_25744 = mux_25744(v_25745);
  assign v_25745 = ~act_8914;
  assign v_25746 = v_25747 | v_25748;
  assign v_25747 = mux_25747(v_8915);
  assign v_25748 = mux_25748(v_8921);
  assign v_25749 = mux_25749(v_8873);
  assign v_25751 = v_25752 | v_25754;
  assign v_25752 = mux_25752(v_25753);
  assign v_25753 = ~act_8009;
  assign v_25754 = v_25755 | v_25861;
  assign v_25755 = mux_25755(v_8010);
  assign v_25757 = v_25758 | v_25760;
  assign v_25758 = mux_25758(v_25759);
  assign v_25759 = ~act_8445;
  assign v_25760 = v_25761 | v_25811;
  assign v_25761 = mux_25761(v_8446);
  assign v_25763 = v_25764 | v_25766;
  assign v_25764 = mux_25764(v_25765);
  assign v_25765 = ~act_8657;
  assign v_25766 = v_25767 | v_25789;
  assign v_25767 = mux_25767(v_8658);
  assign v_25769 = v_25770 | v_25772;
  assign v_25770 = mux_25770(v_25771);
  assign v_25771 = ~act_8757;
  assign v_25772 = v_25773 | v_25781;
  assign v_25773 = mux_25773(v_8758);
  assign v_25775 = v_25776 | v_25778;
  assign v_25776 = mux_25776(v_25777);
  assign v_25777 = ~act_8801;
  assign v_25778 = v_25779 | v_25780;
  assign v_25779 = mux_25779(v_8802);
  assign v_25780 = mux_25780(v_8808);
  assign v_25781 = mux_25781(v_8788);
  assign v_25783 = v_25784 | v_25786;
  assign v_25784 = mux_25784(v_25785);
  assign v_25785 = ~act_8764;
  assign v_25786 = v_25787 | v_25788;
  assign v_25787 = mux_25787(v_8765);
  assign v_25788 = mux_25788(v_8771);
  assign v_25789 = mux_25789(v_8744);
  assign v_25791 = v_25792 | v_25794;
  assign v_25792 = mux_25792(v_25793);
  assign v_25793 = ~act_8664;
  assign v_25794 = v_25795 | v_25803;
  assign v_25795 = mux_25795(v_8665);
  assign v_25797 = v_25798 | v_25800;
  assign v_25798 = mux_25798(v_25799);
  assign v_25799 = ~act_8708;
  assign v_25800 = v_25801 | v_25802;
  assign v_25801 = mux_25801(v_8709);
  assign v_25802 = mux_25802(v_8715);
  assign v_25803 = mux_25803(v_8695);
  assign v_25805 = v_25806 | v_25808;
  assign v_25806 = mux_25806(v_25807);
  assign v_25807 = ~act_8671;
  assign v_25808 = v_25809 | v_25810;
  assign v_25809 = mux_25809(v_8672);
  assign v_25810 = mux_25810(v_8678);
  assign v_25811 = mux_25811(v_8644);
  assign v_25813 = v_25814 | v_25816;
  assign v_25814 = mux_25814(v_25815);
  assign v_25815 = ~act_8452;
  assign v_25816 = v_25817 | v_25839;
  assign v_25817 = mux_25817(v_8453);
  assign v_25819 = v_25820 | v_25822;
  assign v_25820 = mux_25820(v_25821);
  assign v_25821 = ~act_8552;
  assign v_25822 = v_25823 | v_25831;
  assign v_25823 = mux_25823(v_8553);
  assign v_25825 = v_25826 | v_25828;
  assign v_25826 = mux_25826(v_25827);
  assign v_25827 = ~act_8596;
  assign v_25828 = v_25829 | v_25830;
  assign v_25829 = mux_25829(v_8597);
  assign v_25830 = mux_25830(v_8603);
  assign v_25831 = mux_25831(v_8583);
  assign v_25833 = v_25834 | v_25836;
  assign v_25834 = mux_25834(v_25835);
  assign v_25835 = ~act_8559;
  assign v_25836 = v_25837 | v_25838;
  assign v_25837 = mux_25837(v_8560);
  assign v_25838 = mux_25838(v_8566);
  assign v_25839 = mux_25839(v_8539);
  assign v_25841 = v_25842 | v_25844;
  assign v_25842 = mux_25842(v_25843);
  assign v_25843 = ~act_8459;
  assign v_25844 = v_25845 | v_25853;
  assign v_25845 = mux_25845(v_8460);
  assign v_25847 = v_25848 | v_25850;
  assign v_25848 = mux_25848(v_25849);
  assign v_25849 = ~act_8503;
  assign v_25850 = v_25851 | v_25852;
  assign v_25851 = mux_25851(v_8504);
  assign v_25852 = mux_25852(v_8510);
  assign v_25853 = mux_25853(v_8490);
  assign v_25855 = v_25856 | v_25858;
  assign v_25856 = mux_25856(v_25857);
  assign v_25857 = ~act_8466;
  assign v_25858 = v_25859 | v_25860;
  assign v_25859 = mux_25859(v_8467);
  assign v_25860 = mux_25860(v_8473);
  assign v_25861 = mux_25861(v_8432);
  assign v_25863 = v_25864 | v_25866;
  assign v_25864 = mux_25864(v_25865);
  assign v_25865 = ~act_8016;
  assign v_25866 = v_25867 | v_25917;
  assign v_25867 = mux_25867(v_8017);
  assign v_25869 = v_25870 | v_25872;
  assign v_25870 = mux_25870(v_25871);
  assign v_25871 = ~act_8228;
  assign v_25872 = v_25873 | v_25895;
  assign v_25873 = mux_25873(v_8229);
  assign v_25875 = v_25876 | v_25878;
  assign v_25876 = mux_25876(v_25877);
  assign v_25877 = ~act_8328;
  assign v_25878 = v_25879 | v_25887;
  assign v_25879 = mux_25879(v_8329);
  assign v_25881 = v_25882 | v_25884;
  assign v_25882 = mux_25882(v_25883);
  assign v_25883 = ~act_8372;
  assign v_25884 = v_25885 | v_25886;
  assign v_25885 = mux_25885(v_8373);
  assign v_25886 = mux_25886(v_8379);
  assign v_25887 = mux_25887(v_8359);
  assign v_25889 = v_25890 | v_25892;
  assign v_25890 = mux_25890(v_25891);
  assign v_25891 = ~act_8335;
  assign v_25892 = v_25893 | v_25894;
  assign v_25893 = mux_25893(v_8336);
  assign v_25894 = mux_25894(v_8342);
  assign v_25895 = mux_25895(v_8315);
  assign v_25897 = v_25898 | v_25900;
  assign v_25898 = mux_25898(v_25899);
  assign v_25899 = ~act_8235;
  assign v_25900 = v_25901 | v_25909;
  assign v_25901 = mux_25901(v_8236);
  assign v_25903 = v_25904 | v_25906;
  assign v_25904 = mux_25904(v_25905);
  assign v_25905 = ~act_8279;
  assign v_25906 = v_25907 | v_25908;
  assign v_25907 = mux_25907(v_8280);
  assign v_25908 = mux_25908(v_8286);
  assign v_25909 = mux_25909(v_8266);
  assign v_25911 = v_25912 | v_25914;
  assign v_25912 = mux_25912(v_25913);
  assign v_25913 = ~act_8242;
  assign v_25914 = v_25915 | v_25916;
  assign v_25915 = mux_25915(v_8243);
  assign v_25916 = mux_25916(v_8249);
  assign v_25917 = mux_25917(v_8215);
  assign v_25919 = v_25920 | v_25922;
  assign v_25920 = mux_25920(v_25921);
  assign v_25921 = ~act_8023;
  assign v_25922 = v_25923 | v_25945;
  assign v_25923 = mux_25923(v_8024);
  assign v_25925 = v_25926 | v_25928;
  assign v_25926 = mux_25926(v_25927);
  assign v_25927 = ~act_8123;
  assign v_25928 = v_25929 | v_25937;
  assign v_25929 = mux_25929(v_8124);
  assign v_25931 = v_25932 | v_25934;
  assign v_25932 = mux_25932(v_25933);
  assign v_25933 = ~act_8167;
  assign v_25934 = v_25935 | v_25936;
  assign v_25935 = mux_25935(v_8168);
  assign v_25936 = mux_25936(v_8174);
  assign v_25937 = mux_25937(v_8154);
  assign v_25939 = v_25940 | v_25942;
  assign v_25940 = mux_25940(v_25941);
  assign v_25941 = ~act_8130;
  assign v_25942 = v_25943 | v_25944;
  assign v_25943 = mux_25943(v_8131);
  assign v_25944 = mux_25944(v_8137);
  assign v_25945 = mux_25945(v_8110);
  assign v_25947 = v_25948 | v_25950;
  assign v_25948 = mux_25948(v_25949);
  assign v_25949 = ~act_8030;
  assign v_25950 = v_25951 | v_25959;
  assign v_25951 = mux_25951(v_8031);
  assign v_25953 = v_25954 | v_25956;
  assign v_25954 = mux_25954(v_25955);
  assign v_25955 = ~act_8074;
  assign v_25956 = v_25957 | v_25958;
  assign v_25957 = mux_25957(v_8075);
  assign v_25958 = mux_25958(v_8081);
  assign v_25959 = mux_25959(v_8061);
  assign v_25961 = v_25962 | v_25964;
  assign v_25962 = mux_25962(v_25963);
  assign v_25963 = ~act_8037;
  assign v_25964 = v_25965 | v_25966;
  assign v_25965 = mux_25965(v_8038);
  assign v_25966 = mux_25966(v_8044);
  assign v_25967 = mux_25967(v_7967);
  assign v_25969 = v_25970 | v_25972;
  assign v_25970 = mux_25970(v_25971);
  assign v_25971 = ~act_7960;
  assign v_25972 = v_25973 | v_27087;
  assign v_25973 = mux_25973(v_4395);
  assign v_25975 = v_25976 | v_25978;
  assign v_25976 = mux_25976(v_25977);
  assign v_25977 = ~act_4388;
  assign v_25978 = v_25979 | v_26645;
  assign v_25979 = mux_25979(v_2615);
  assign v_25981 = v_25982 | v_25984;
  assign v_25982 = mux_25982(v_25983);
  assign v_25983 = ~act_2608;
  assign v_25984 = v_25985 | v_26427;
  assign v_25985 = mux_25985(v_1731);
  assign v_25987 = v_25988 | v_25990;
  assign v_25988 = mux_25988(v_25989);
  assign v_25989 = ~act_848;
  assign v_25990 = v_25991 | v_26209;
  assign v_25991 = mux_25991(v_849);
  assign v_25993 = v_25994 | v_25996;
  assign v_25994 = mux_25994(v_25995);
  assign v_25995 = ~act_855;
  assign v_25996 = v_25997 | v_26103;
  assign v_25997 = mux_25997(v_856);
  assign v_25999 = v_26000 | v_26002;
  assign v_26000 = mux_26000(v_26001);
  assign v_26001 = ~act_1291;
  assign v_26002 = v_26003 | v_26053;
  assign v_26003 = mux_26003(v_1292);
  assign v_26005 = v_26006 | v_26008;
  assign v_26006 = mux_26006(v_26007);
  assign v_26007 = ~act_1503;
  assign v_26008 = v_26009 | v_26031;
  assign v_26009 = mux_26009(v_1504);
  assign v_26011 = v_26012 | v_26014;
  assign v_26012 = mux_26012(v_26013);
  assign v_26013 = ~act_1603;
  assign v_26014 = v_26015 | v_26023;
  assign v_26015 = mux_26015(v_1604);
  assign v_26017 = v_26018 | v_26020;
  assign v_26018 = mux_26018(v_26019);
  assign v_26019 = ~act_1647;
  assign v_26020 = v_26021 | v_26022;
  assign v_26021 = mux_26021(v_1648);
  assign v_26022 = mux_26022(v_1654);
  assign v_26023 = mux_26023(v_1634);
  assign v_26025 = v_26026 | v_26028;
  assign v_26026 = mux_26026(v_26027);
  assign v_26027 = ~act_1610;
  assign v_26028 = v_26029 | v_26030;
  assign v_26029 = mux_26029(v_1611);
  assign v_26030 = mux_26030(v_1617);
  assign v_26031 = mux_26031(v_1590);
  assign v_26033 = v_26034 | v_26036;
  assign v_26034 = mux_26034(v_26035);
  assign v_26035 = ~act_1510;
  assign v_26036 = v_26037 | v_26045;
  assign v_26037 = mux_26037(v_1511);
  assign v_26039 = v_26040 | v_26042;
  assign v_26040 = mux_26040(v_26041);
  assign v_26041 = ~act_1554;
  assign v_26042 = v_26043 | v_26044;
  assign v_26043 = mux_26043(v_1555);
  assign v_26044 = mux_26044(v_1561);
  assign v_26045 = mux_26045(v_1541);
  assign v_26047 = v_26048 | v_26050;
  assign v_26048 = mux_26048(v_26049);
  assign v_26049 = ~act_1517;
  assign v_26050 = v_26051 | v_26052;
  assign v_26051 = mux_26051(v_1518);
  assign v_26052 = mux_26052(v_1524);
  assign v_26053 = mux_26053(v_1490);
  assign v_26055 = v_26056 | v_26058;
  assign v_26056 = mux_26056(v_26057);
  assign v_26057 = ~act_1298;
  assign v_26058 = v_26059 | v_26081;
  assign v_26059 = mux_26059(v_1299);
  assign v_26061 = v_26062 | v_26064;
  assign v_26062 = mux_26062(v_26063);
  assign v_26063 = ~act_1398;
  assign v_26064 = v_26065 | v_26073;
  assign v_26065 = mux_26065(v_1399);
  assign v_26067 = v_26068 | v_26070;
  assign v_26068 = mux_26068(v_26069);
  assign v_26069 = ~act_1442;
  assign v_26070 = v_26071 | v_26072;
  assign v_26071 = mux_26071(v_1443);
  assign v_26072 = mux_26072(v_1449);
  assign v_26073 = mux_26073(v_1429);
  assign v_26075 = v_26076 | v_26078;
  assign v_26076 = mux_26076(v_26077);
  assign v_26077 = ~act_1405;
  assign v_26078 = v_26079 | v_26080;
  assign v_26079 = mux_26079(v_1406);
  assign v_26080 = mux_26080(v_1412);
  assign v_26081 = mux_26081(v_1385);
  assign v_26083 = v_26084 | v_26086;
  assign v_26084 = mux_26084(v_26085);
  assign v_26085 = ~act_1305;
  assign v_26086 = v_26087 | v_26095;
  assign v_26087 = mux_26087(v_1306);
  assign v_26089 = v_26090 | v_26092;
  assign v_26090 = mux_26090(v_26091);
  assign v_26091 = ~act_1349;
  assign v_26092 = v_26093 | v_26094;
  assign v_26093 = mux_26093(v_1350);
  assign v_26094 = mux_26094(v_1356);
  assign v_26095 = mux_26095(v_1336);
  assign v_26097 = v_26098 | v_26100;
  assign v_26098 = mux_26098(v_26099);
  assign v_26099 = ~act_1312;
  assign v_26100 = v_26101 | v_26102;
  assign v_26101 = mux_26101(v_1313);
  assign v_26102 = mux_26102(v_1319);
  assign v_26103 = mux_26103(v_1278);
  assign v_26105 = v_26106 | v_26108;
  assign v_26106 = mux_26106(v_26107);
  assign v_26107 = ~act_862;
  assign v_26108 = v_26109 | v_26159;
  assign v_26109 = mux_26109(v_863);
  assign v_26111 = v_26112 | v_26114;
  assign v_26112 = mux_26112(v_26113);
  assign v_26113 = ~act_1074;
  assign v_26114 = v_26115 | v_26137;
  assign v_26115 = mux_26115(v_1075);
  assign v_26117 = v_26118 | v_26120;
  assign v_26118 = mux_26118(v_26119);
  assign v_26119 = ~act_1174;
  assign v_26120 = v_26121 | v_26129;
  assign v_26121 = mux_26121(v_1175);
  assign v_26123 = v_26124 | v_26126;
  assign v_26124 = mux_26124(v_26125);
  assign v_26125 = ~act_1218;
  assign v_26126 = v_26127 | v_26128;
  assign v_26127 = mux_26127(v_1219);
  assign v_26128 = mux_26128(v_1225);
  assign v_26129 = mux_26129(v_1205);
  assign v_26131 = v_26132 | v_26134;
  assign v_26132 = mux_26132(v_26133);
  assign v_26133 = ~act_1181;
  assign v_26134 = v_26135 | v_26136;
  assign v_26135 = mux_26135(v_1182);
  assign v_26136 = mux_26136(v_1188);
  assign v_26137 = mux_26137(v_1161);
  assign v_26139 = v_26140 | v_26142;
  assign v_26140 = mux_26140(v_26141);
  assign v_26141 = ~act_1081;
  assign v_26142 = v_26143 | v_26151;
  assign v_26143 = mux_26143(v_1082);
  assign v_26145 = v_26146 | v_26148;
  assign v_26146 = mux_26146(v_26147);
  assign v_26147 = ~act_1125;
  assign v_26148 = v_26149 | v_26150;
  assign v_26149 = mux_26149(v_1126);
  assign v_26150 = mux_26150(v_1132);
  assign v_26151 = mux_26151(v_1112);
  assign v_26153 = v_26154 | v_26156;
  assign v_26154 = mux_26154(v_26155);
  assign v_26155 = ~act_1088;
  assign v_26156 = v_26157 | v_26158;
  assign v_26157 = mux_26157(v_1089);
  assign v_26158 = mux_26158(v_1095);
  assign v_26159 = mux_26159(v_1061);
  assign v_26161 = v_26162 | v_26164;
  assign v_26162 = mux_26162(v_26163);
  assign v_26163 = ~act_869;
  assign v_26164 = v_26165 | v_26187;
  assign v_26165 = mux_26165(v_870);
  assign v_26167 = v_26168 | v_26170;
  assign v_26168 = mux_26168(v_26169);
  assign v_26169 = ~act_969;
  assign v_26170 = v_26171 | v_26179;
  assign v_26171 = mux_26171(v_970);
  assign v_26173 = v_26174 | v_26176;
  assign v_26174 = mux_26174(v_26175);
  assign v_26175 = ~act_1013;
  assign v_26176 = v_26177 | v_26178;
  assign v_26177 = mux_26177(v_1014);
  assign v_26178 = mux_26178(v_1020);
  assign v_26179 = mux_26179(v_1000);
  assign v_26181 = v_26182 | v_26184;
  assign v_26182 = mux_26182(v_26183);
  assign v_26183 = ~act_976;
  assign v_26184 = v_26185 | v_26186;
  assign v_26185 = mux_26185(v_977);
  assign v_26186 = mux_26186(v_983);
  assign v_26187 = mux_26187(v_956);
  assign v_26189 = v_26190 | v_26192;
  assign v_26190 = mux_26190(v_26191);
  assign v_26191 = ~act_876;
  assign v_26192 = v_26193 | v_26201;
  assign v_26193 = mux_26193(v_877);
  assign v_26195 = v_26196 | v_26198;
  assign v_26196 = mux_26196(v_26197);
  assign v_26197 = ~act_920;
  assign v_26198 = v_26199 | v_26200;
  assign v_26199 = mux_26199(v_921);
  assign v_26200 = mux_26200(v_927);
  assign v_26201 = mux_26201(v_907);
  assign v_26203 = v_26204 | v_26206;
  assign v_26204 = mux_26204(v_26205);
  assign v_26205 = ~act_883;
  assign v_26206 = v_26207 | v_26208;
  assign v_26207 = mux_26207(v_884);
  assign v_26208 = mux_26208(v_890);
  assign v_26209 = mux_26209(v_841);
  assign v_26211 = v_26212 | v_26214;
  assign v_26212 = mux_26212(v_26213);
  assign v_26213 = ~act_406;
  assign v_26214 = v_26215 | v_26321;
  assign v_26215 = mux_26215(v_407);
  assign v_26217 = v_26218 | v_26220;
  assign v_26218 = mux_26218(v_26219);
  assign v_26219 = ~act_413;
  assign v_26220 = v_26221 | v_26271;
  assign v_26221 = mux_26221(v_414);
  assign v_26223 = v_26224 | v_26226;
  assign v_26224 = mux_26224(v_26225);
  assign v_26225 = ~act_625;
  assign v_26226 = v_26227 | v_26249;
  assign v_26227 = mux_26227(v_626);
  assign v_26229 = v_26230 | v_26232;
  assign v_26230 = mux_26230(v_26231);
  assign v_26231 = ~act_725;
  assign v_26232 = v_26233 | v_26241;
  assign v_26233 = mux_26233(v_726);
  assign v_26235 = v_26236 | v_26238;
  assign v_26236 = mux_26236(v_26237);
  assign v_26237 = ~act_769;
  assign v_26238 = v_26239 | v_26240;
  assign v_26239 = mux_26239(v_770);
  assign v_26240 = mux_26240(v_776);
  assign v_26241 = mux_26241(v_756);
  assign v_26243 = v_26244 | v_26246;
  assign v_26244 = mux_26244(v_26245);
  assign v_26245 = ~act_732;
  assign v_26246 = v_26247 | v_26248;
  assign v_26247 = mux_26247(v_733);
  assign v_26248 = mux_26248(v_739);
  assign v_26249 = mux_26249(v_712);
  assign v_26251 = v_26252 | v_26254;
  assign v_26252 = mux_26252(v_26253);
  assign v_26253 = ~act_632;
  assign v_26254 = v_26255 | v_26263;
  assign v_26255 = mux_26255(v_633);
  assign v_26257 = v_26258 | v_26260;
  assign v_26258 = mux_26258(v_26259);
  assign v_26259 = ~act_676;
  assign v_26260 = v_26261 | v_26262;
  assign v_26261 = mux_26261(v_677);
  assign v_26262 = mux_26262(v_683);
  assign v_26263 = mux_26263(v_663);
  assign v_26265 = v_26266 | v_26268;
  assign v_26266 = mux_26266(v_26267);
  assign v_26267 = ~act_639;
  assign v_26268 = v_26269 | v_26270;
  assign v_26269 = mux_26269(v_640);
  assign v_26270 = mux_26270(v_646);
  assign v_26271 = mux_26271(v_612);
  assign v_26273 = v_26274 | v_26276;
  assign v_26274 = mux_26274(v_26275);
  assign v_26275 = ~act_420;
  assign v_26276 = v_26277 | v_26299;
  assign v_26277 = mux_26277(v_421);
  assign v_26279 = v_26280 | v_26282;
  assign v_26280 = mux_26280(v_26281);
  assign v_26281 = ~act_520;
  assign v_26282 = v_26283 | v_26291;
  assign v_26283 = mux_26283(v_521);
  assign v_26285 = v_26286 | v_26288;
  assign v_26286 = mux_26286(v_26287);
  assign v_26287 = ~act_564;
  assign v_26288 = v_26289 | v_26290;
  assign v_26289 = mux_26289(v_565);
  assign v_26290 = mux_26290(v_571);
  assign v_26291 = mux_26291(v_551);
  assign v_26293 = v_26294 | v_26296;
  assign v_26294 = mux_26294(v_26295);
  assign v_26295 = ~act_527;
  assign v_26296 = v_26297 | v_26298;
  assign v_26297 = mux_26297(v_528);
  assign v_26298 = mux_26298(v_534);
  assign v_26299 = mux_26299(v_507);
  assign v_26301 = v_26302 | v_26304;
  assign v_26302 = mux_26302(v_26303);
  assign v_26303 = ~act_427;
  assign v_26304 = v_26305 | v_26313;
  assign v_26305 = mux_26305(v_428);
  assign v_26307 = v_26308 | v_26310;
  assign v_26308 = mux_26308(v_26309);
  assign v_26309 = ~act_471;
  assign v_26310 = v_26311 | v_26312;
  assign v_26311 = mux_26311(v_472);
  assign v_26312 = mux_26312(v_478);
  assign v_26313 = mux_26313(v_458);
  assign v_26315 = v_26316 | v_26318;
  assign v_26316 = mux_26316(v_26317);
  assign v_26317 = ~act_434;
  assign v_26318 = v_26319 | v_26320;
  assign v_26319 = mux_26319(v_435);
  assign v_26320 = mux_26320(v_441);
  assign v_26321 = mux_26321(v_399);
  assign v_26323 = v_26324 | v_26326;
  assign v_26324 = mux_26324(v_26325);
  assign v_26325 = ~act_188;
  assign v_26326 = v_26327 | v_26377;
  assign v_26327 = mux_26327(v_189);
  assign v_26329 = v_26330 | v_26332;
  assign v_26330 = mux_26330(v_26331);
  assign v_26331 = ~act_195;
  assign v_26332 = v_26333 | v_26355;
  assign v_26333 = mux_26333(v_196);
  assign v_26335 = v_26336 | v_26338;
  assign v_26336 = mux_26336(v_26337);
  assign v_26337 = ~act_295;
  assign v_26338 = v_26339 | v_26347;
  assign v_26339 = mux_26339(v_296);
  assign v_26341 = v_26342 | v_26344;
  assign v_26342 = mux_26342(v_26343);
  assign v_26343 = ~act_339;
  assign v_26344 = v_26345 | v_26346;
  assign v_26345 = mux_26345(v_340);
  assign v_26346 = mux_26346(v_346);
  assign v_26347 = mux_26347(v_326);
  assign v_26349 = v_26350 | v_26352;
  assign v_26350 = mux_26350(v_26351);
  assign v_26351 = ~act_302;
  assign v_26352 = v_26353 | v_26354;
  assign v_26353 = mux_26353(v_303);
  assign v_26354 = mux_26354(v_309);
  assign v_26355 = mux_26355(v_282);
  assign v_26357 = v_26358 | v_26360;
  assign v_26358 = mux_26358(v_26359);
  assign v_26359 = ~act_202;
  assign v_26360 = v_26361 | v_26369;
  assign v_26361 = mux_26361(v_203);
  assign v_26363 = v_26364 | v_26366;
  assign v_26364 = mux_26364(v_26365);
  assign v_26365 = ~act_246;
  assign v_26366 = v_26367 | v_26368;
  assign v_26367 = mux_26367(v_247);
  assign v_26368 = mux_26368(v_253);
  assign v_26369 = mux_26369(v_233);
  assign v_26371 = v_26372 | v_26374;
  assign v_26372 = mux_26372(v_26373);
  assign v_26373 = ~act_209;
  assign v_26374 = v_26375 | v_26376;
  assign v_26375 = mux_26375(v_210);
  assign v_26376 = mux_26376(v_216);
  assign v_26377 = mux_26377(v_181);
  assign v_26379 = v_26380 | v_26382;
  assign v_26380 = mux_26380(v_26381);
  assign v_26381 = ~act_82;
  assign v_26382 = v_26383 | v_26405;
  assign v_26383 = mux_26383(v_83);
  assign v_26385 = v_26386 | v_26388;
  assign v_26386 = mux_26386(v_26387);
  assign v_26387 = ~act_89;
  assign v_26388 = v_26389 | v_26397;
  assign v_26389 = mux_26389(v_90);
  assign v_26391 = v_26392 | v_26394;
  assign v_26392 = mux_26392(v_26393);
  assign v_26393 = ~act_133;
  assign v_26394 = v_26395 | v_26396;
  assign v_26395 = mux_26395(v_134);
  assign v_26396 = mux_26396(v_140);
  assign v_26397 = mux_26397(v_120);
  assign v_26399 = v_26400 | v_26402;
  assign v_26400 = mux_26400(v_26401);
  assign v_26401 = ~act_96;
  assign v_26402 = v_26403 | v_26404;
  assign v_26403 = mux_26403(v_97);
  assign v_26404 = mux_26404(v_103);
  assign v_26405 = mux_26405(v_75);
  assign v_26407 = v_26408 | v_26410;
  assign v_26408 = mux_26408(v_26409);
  assign v_26409 = ~act_32;
  assign v_26410 = v_26411 | v_26419;
  assign v_26411 = mux_26411(v_33);
  assign v_26413 = v_26414 | v_26416;
  assign v_26414 = mux_26414(v_26415);
  assign v_26415 = ~act_39;
  assign v_26416 = v_26417 | v_26418;
  assign v_26417 = mux_26417(v_40);
  assign v_26418 = mux_26418(v_46);
  assign v_26419 = mux_26419(v_25);
  assign v_26421 = v_26422 | v_26424;
  assign v_26422 = mux_26422(v_26423);
  assign v_26423 = ~act_10;
  assign v_26424 = v_26425 | v_26426;
  assign v_26425 = mux_26425(v_11);
  assign v_26426 = mux_26426(v_2);
  assign v_26427 = mux_26427(v_2601);
  assign v_26429 = v_26430 | v_26432;
  assign v_26430 = mux_26430(v_26431);
  assign v_26431 = ~act_1737;
  assign v_26432 = v_26433 | v_26539;
  assign v_26433 = mux_26433(v_1738);
  assign v_26435 = v_26436 | v_26438;
  assign v_26436 = mux_26436(v_26437);
  assign v_26437 = ~act_2173;
  assign v_26438 = v_26439 | v_26489;
  assign v_26439 = mux_26439(v_2174);
  assign v_26441 = v_26442 | v_26444;
  assign v_26442 = mux_26442(v_26443);
  assign v_26443 = ~act_2385;
  assign v_26444 = v_26445 | v_26467;
  assign v_26445 = mux_26445(v_2386);
  assign v_26447 = v_26448 | v_26450;
  assign v_26448 = mux_26448(v_26449);
  assign v_26449 = ~act_2485;
  assign v_26450 = v_26451 | v_26459;
  assign v_26451 = mux_26451(v_2486);
  assign v_26453 = v_26454 | v_26456;
  assign v_26454 = mux_26454(v_26455);
  assign v_26455 = ~act_2529;
  assign v_26456 = v_26457 | v_26458;
  assign v_26457 = mux_26457(v_2530);
  assign v_26458 = mux_26458(v_2536);
  assign v_26459 = mux_26459(v_2516);
  assign v_26461 = v_26462 | v_26464;
  assign v_26462 = mux_26462(v_26463);
  assign v_26463 = ~act_2492;
  assign v_26464 = v_26465 | v_26466;
  assign v_26465 = mux_26465(v_2493);
  assign v_26466 = mux_26466(v_2499);
  assign v_26467 = mux_26467(v_2472);
  assign v_26469 = v_26470 | v_26472;
  assign v_26470 = mux_26470(v_26471);
  assign v_26471 = ~act_2392;
  assign v_26472 = v_26473 | v_26481;
  assign v_26473 = mux_26473(v_2393);
  assign v_26475 = v_26476 | v_26478;
  assign v_26476 = mux_26476(v_26477);
  assign v_26477 = ~act_2436;
  assign v_26478 = v_26479 | v_26480;
  assign v_26479 = mux_26479(v_2437);
  assign v_26480 = mux_26480(v_2443);
  assign v_26481 = mux_26481(v_2423);
  assign v_26483 = v_26484 | v_26486;
  assign v_26484 = mux_26484(v_26485);
  assign v_26485 = ~act_2399;
  assign v_26486 = v_26487 | v_26488;
  assign v_26487 = mux_26487(v_2400);
  assign v_26488 = mux_26488(v_2406);
  assign v_26489 = mux_26489(v_2372);
  assign v_26491 = v_26492 | v_26494;
  assign v_26492 = mux_26492(v_26493);
  assign v_26493 = ~act_2180;
  assign v_26494 = v_26495 | v_26517;
  assign v_26495 = mux_26495(v_2181);
  assign v_26497 = v_26498 | v_26500;
  assign v_26498 = mux_26498(v_26499);
  assign v_26499 = ~act_2280;
  assign v_26500 = v_26501 | v_26509;
  assign v_26501 = mux_26501(v_2281);
  assign v_26503 = v_26504 | v_26506;
  assign v_26504 = mux_26504(v_26505);
  assign v_26505 = ~act_2324;
  assign v_26506 = v_26507 | v_26508;
  assign v_26507 = mux_26507(v_2325);
  assign v_26508 = mux_26508(v_2331);
  assign v_26509 = mux_26509(v_2311);
  assign v_26511 = v_26512 | v_26514;
  assign v_26512 = mux_26512(v_26513);
  assign v_26513 = ~act_2287;
  assign v_26514 = v_26515 | v_26516;
  assign v_26515 = mux_26515(v_2288);
  assign v_26516 = mux_26516(v_2294);
  assign v_26517 = mux_26517(v_2267);
  assign v_26519 = v_26520 | v_26522;
  assign v_26520 = mux_26520(v_26521);
  assign v_26521 = ~act_2187;
  assign v_26522 = v_26523 | v_26531;
  assign v_26523 = mux_26523(v_2188);
  assign v_26525 = v_26526 | v_26528;
  assign v_26526 = mux_26526(v_26527);
  assign v_26527 = ~act_2231;
  assign v_26528 = v_26529 | v_26530;
  assign v_26529 = mux_26529(v_2232);
  assign v_26530 = mux_26530(v_2238);
  assign v_26531 = mux_26531(v_2218);
  assign v_26533 = v_26534 | v_26536;
  assign v_26534 = mux_26534(v_26535);
  assign v_26535 = ~act_2194;
  assign v_26536 = v_26537 | v_26538;
  assign v_26537 = mux_26537(v_2195);
  assign v_26538 = mux_26538(v_2201);
  assign v_26539 = mux_26539(v_2160);
  assign v_26541 = v_26542 | v_26544;
  assign v_26542 = mux_26542(v_26543);
  assign v_26543 = ~act_1744;
  assign v_26544 = v_26545 | v_26595;
  assign v_26545 = mux_26545(v_1745);
  assign v_26547 = v_26548 | v_26550;
  assign v_26548 = mux_26548(v_26549);
  assign v_26549 = ~act_1956;
  assign v_26550 = v_26551 | v_26573;
  assign v_26551 = mux_26551(v_1957);
  assign v_26553 = v_26554 | v_26556;
  assign v_26554 = mux_26554(v_26555);
  assign v_26555 = ~act_2056;
  assign v_26556 = v_26557 | v_26565;
  assign v_26557 = mux_26557(v_2057);
  assign v_26559 = v_26560 | v_26562;
  assign v_26560 = mux_26560(v_26561);
  assign v_26561 = ~act_2100;
  assign v_26562 = v_26563 | v_26564;
  assign v_26563 = mux_26563(v_2101);
  assign v_26564 = mux_26564(v_2107);
  assign v_26565 = mux_26565(v_2087);
  assign v_26567 = v_26568 | v_26570;
  assign v_26568 = mux_26568(v_26569);
  assign v_26569 = ~act_2063;
  assign v_26570 = v_26571 | v_26572;
  assign v_26571 = mux_26571(v_2064);
  assign v_26572 = mux_26572(v_2070);
  assign v_26573 = mux_26573(v_2043);
  assign v_26575 = v_26576 | v_26578;
  assign v_26576 = mux_26576(v_26577);
  assign v_26577 = ~act_1963;
  assign v_26578 = v_26579 | v_26587;
  assign v_26579 = mux_26579(v_1964);
  assign v_26581 = v_26582 | v_26584;
  assign v_26582 = mux_26582(v_26583);
  assign v_26583 = ~act_2007;
  assign v_26584 = v_26585 | v_26586;
  assign v_26585 = mux_26585(v_2008);
  assign v_26586 = mux_26586(v_2014);
  assign v_26587 = mux_26587(v_1994);
  assign v_26589 = v_26590 | v_26592;
  assign v_26590 = mux_26590(v_26591);
  assign v_26591 = ~act_1970;
  assign v_26592 = v_26593 | v_26594;
  assign v_26593 = mux_26593(v_1971);
  assign v_26594 = mux_26594(v_1977);
  assign v_26595 = mux_26595(v_1943);
  assign v_26597 = v_26598 | v_26600;
  assign v_26598 = mux_26598(v_26599);
  assign v_26599 = ~act_1751;
  assign v_26600 = v_26601 | v_26623;
  assign v_26601 = mux_26601(v_1752);
  assign v_26603 = v_26604 | v_26606;
  assign v_26604 = mux_26604(v_26605);
  assign v_26605 = ~act_1851;
  assign v_26606 = v_26607 | v_26615;
  assign v_26607 = mux_26607(v_1852);
  assign v_26609 = v_26610 | v_26612;
  assign v_26610 = mux_26610(v_26611);
  assign v_26611 = ~act_1895;
  assign v_26612 = v_26613 | v_26614;
  assign v_26613 = mux_26613(v_1896);
  assign v_26614 = mux_26614(v_1902);
  assign v_26615 = mux_26615(v_1882);
  assign v_26617 = v_26618 | v_26620;
  assign v_26618 = mux_26618(v_26619);
  assign v_26619 = ~act_1858;
  assign v_26620 = v_26621 | v_26622;
  assign v_26621 = mux_26621(v_1859);
  assign v_26622 = mux_26622(v_1865);
  assign v_26623 = mux_26623(v_1838);
  assign v_26625 = v_26626 | v_26628;
  assign v_26626 = mux_26626(v_26627);
  assign v_26627 = ~act_1758;
  assign v_26628 = v_26629 | v_26637;
  assign v_26629 = mux_26629(v_1759);
  assign v_26631 = v_26632 | v_26634;
  assign v_26632 = mux_26632(v_26633);
  assign v_26633 = ~act_1802;
  assign v_26634 = v_26635 | v_26636;
  assign v_26635 = mux_26635(v_1803);
  assign v_26636 = mux_26636(v_1809);
  assign v_26637 = mux_26637(v_1789);
  assign v_26639 = v_26640 | v_26642;
  assign v_26640 = mux_26640(v_26641);
  assign v_26641 = ~act_1765;
  assign v_26642 = v_26643 | v_26644;
  assign v_26643 = mux_26643(v_1766);
  assign v_26644 = mux_26644(v_1772);
  assign v_26645 = mux_26645(v_4381);
  assign v_26647 = v_26648 | v_26650;
  assign v_26648 = mux_26648(v_26649);
  assign v_26649 = ~act_2621;
  assign v_26650 = v_26651 | v_26869;
  assign v_26651 = mux_26651(v_2622);
  assign v_26653 = v_26654 | v_26656;
  assign v_26654 = mux_26654(v_26655);
  assign v_26655 = ~act_3505;
  assign v_26656 = v_26657 | v_26763;
  assign v_26657 = mux_26657(v_3506);
  assign v_26659 = v_26660 | v_26662;
  assign v_26660 = mux_26660(v_26661);
  assign v_26661 = ~act_3941;
  assign v_26662 = v_26663 | v_26713;
  assign v_26663 = mux_26663(v_3942);
  assign v_26665 = v_26666 | v_26668;
  assign v_26666 = mux_26666(v_26667);
  assign v_26667 = ~act_4153;
  assign v_26668 = v_26669 | v_26691;
  assign v_26669 = mux_26669(v_4154);
  assign v_26671 = v_26672 | v_26674;
  assign v_26672 = mux_26672(v_26673);
  assign v_26673 = ~act_4253;
  assign v_26674 = v_26675 | v_26683;
  assign v_26675 = mux_26675(v_4254);
  assign v_26677 = v_26678 | v_26680;
  assign v_26678 = mux_26678(v_26679);
  assign v_26679 = ~act_4297;
  assign v_26680 = v_26681 | v_26682;
  assign v_26681 = mux_26681(v_4298);
  assign v_26682 = mux_26682(v_4304);
  assign v_26683 = mux_26683(v_4284);
  assign v_26685 = v_26686 | v_26688;
  assign v_26686 = mux_26686(v_26687);
  assign v_26687 = ~act_4260;
  assign v_26688 = v_26689 | v_26690;
  assign v_26689 = mux_26689(v_4261);
  assign v_26690 = mux_26690(v_4267);
  assign v_26691 = mux_26691(v_4240);
  assign v_26693 = v_26694 | v_26696;
  assign v_26694 = mux_26694(v_26695);
  assign v_26695 = ~act_4160;
  assign v_26696 = v_26697 | v_26705;
  assign v_26697 = mux_26697(v_4161);
  assign v_26699 = v_26700 | v_26702;
  assign v_26700 = mux_26700(v_26701);
  assign v_26701 = ~act_4204;
  assign v_26702 = v_26703 | v_26704;
  assign v_26703 = mux_26703(v_4205);
  assign v_26704 = mux_26704(v_4211);
  assign v_26705 = mux_26705(v_4191);
  assign v_26707 = v_26708 | v_26710;
  assign v_26708 = mux_26708(v_26709);
  assign v_26709 = ~act_4167;
  assign v_26710 = v_26711 | v_26712;
  assign v_26711 = mux_26711(v_4168);
  assign v_26712 = mux_26712(v_4174);
  assign v_26713 = mux_26713(v_4140);
  assign v_26715 = v_26716 | v_26718;
  assign v_26716 = mux_26716(v_26717);
  assign v_26717 = ~act_3948;
  assign v_26718 = v_26719 | v_26741;
  assign v_26719 = mux_26719(v_3949);
  assign v_26721 = v_26722 | v_26724;
  assign v_26722 = mux_26722(v_26723);
  assign v_26723 = ~act_4048;
  assign v_26724 = v_26725 | v_26733;
  assign v_26725 = mux_26725(v_4049);
  assign v_26727 = v_26728 | v_26730;
  assign v_26728 = mux_26728(v_26729);
  assign v_26729 = ~act_4092;
  assign v_26730 = v_26731 | v_26732;
  assign v_26731 = mux_26731(v_4093);
  assign v_26732 = mux_26732(v_4099);
  assign v_26733 = mux_26733(v_4079);
  assign v_26735 = v_26736 | v_26738;
  assign v_26736 = mux_26736(v_26737);
  assign v_26737 = ~act_4055;
  assign v_26738 = v_26739 | v_26740;
  assign v_26739 = mux_26739(v_4056);
  assign v_26740 = mux_26740(v_4062);
  assign v_26741 = mux_26741(v_4035);
  assign v_26743 = v_26744 | v_26746;
  assign v_26744 = mux_26744(v_26745);
  assign v_26745 = ~act_3955;
  assign v_26746 = v_26747 | v_26755;
  assign v_26747 = mux_26747(v_3956);
  assign v_26749 = v_26750 | v_26752;
  assign v_26750 = mux_26750(v_26751);
  assign v_26751 = ~act_3999;
  assign v_26752 = v_26753 | v_26754;
  assign v_26753 = mux_26753(v_4000);
  assign v_26754 = mux_26754(v_4006);
  assign v_26755 = mux_26755(v_3986);
  assign v_26757 = v_26758 | v_26760;
  assign v_26758 = mux_26758(v_26759);
  assign v_26759 = ~act_3962;
  assign v_26760 = v_26761 | v_26762;
  assign v_26761 = mux_26761(v_3963);
  assign v_26762 = mux_26762(v_3969);
  assign v_26763 = mux_26763(v_3928);
  assign v_26765 = v_26766 | v_26768;
  assign v_26766 = mux_26766(v_26767);
  assign v_26767 = ~act_3512;
  assign v_26768 = v_26769 | v_26819;
  assign v_26769 = mux_26769(v_3513);
  assign v_26771 = v_26772 | v_26774;
  assign v_26772 = mux_26772(v_26773);
  assign v_26773 = ~act_3724;
  assign v_26774 = v_26775 | v_26797;
  assign v_26775 = mux_26775(v_3725);
  assign v_26777 = v_26778 | v_26780;
  assign v_26778 = mux_26778(v_26779);
  assign v_26779 = ~act_3824;
  assign v_26780 = v_26781 | v_26789;
  assign v_26781 = mux_26781(v_3825);
  assign v_26783 = v_26784 | v_26786;
  assign v_26784 = mux_26784(v_26785);
  assign v_26785 = ~act_3868;
  assign v_26786 = v_26787 | v_26788;
  assign v_26787 = mux_26787(v_3869);
  assign v_26788 = mux_26788(v_3875);
  assign v_26789 = mux_26789(v_3855);
  assign v_26791 = v_26792 | v_26794;
  assign v_26792 = mux_26792(v_26793);
  assign v_26793 = ~act_3831;
  assign v_26794 = v_26795 | v_26796;
  assign v_26795 = mux_26795(v_3832);
  assign v_26796 = mux_26796(v_3838);
  assign v_26797 = mux_26797(v_3811);
  assign v_26799 = v_26800 | v_26802;
  assign v_26800 = mux_26800(v_26801);
  assign v_26801 = ~act_3731;
  assign v_26802 = v_26803 | v_26811;
  assign v_26803 = mux_26803(v_3732);
  assign v_26805 = v_26806 | v_26808;
  assign v_26806 = mux_26806(v_26807);
  assign v_26807 = ~act_3775;
  assign v_26808 = v_26809 | v_26810;
  assign v_26809 = mux_26809(v_3776);
  assign v_26810 = mux_26810(v_3782);
  assign v_26811 = mux_26811(v_3762);
  assign v_26813 = v_26814 | v_26816;
  assign v_26814 = mux_26814(v_26815);
  assign v_26815 = ~act_3738;
  assign v_26816 = v_26817 | v_26818;
  assign v_26817 = mux_26817(v_3739);
  assign v_26818 = mux_26818(v_3745);
  assign v_26819 = mux_26819(v_3711);
  assign v_26821 = v_26822 | v_26824;
  assign v_26822 = mux_26822(v_26823);
  assign v_26823 = ~act_3519;
  assign v_26824 = v_26825 | v_26847;
  assign v_26825 = mux_26825(v_3520);
  assign v_26827 = v_26828 | v_26830;
  assign v_26828 = mux_26828(v_26829);
  assign v_26829 = ~act_3619;
  assign v_26830 = v_26831 | v_26839;
  assign v_26831 = mux_26831(v_3620);
  assign v_26833 = v_26834 | v_26836;
  assign v_26834 = mux_26834(v_26835);
  assign v_26835 = ~act_3663;
  assign v_26836 = v_26837 | v_26838;
  assign v_26837 = mux_26837(v_3664);
  assign v_26838 = mux_26838(v_3670);
  assign v_26839 = mux_26839(v_3650);
  assign v_26841 = v_26842 | v_26844;
  assign v_26842 = mux_26842(v_26843);
  assign v_26843 = ~act_3626;
  assign v_26844 = v_26845 | v_26846;
  assign v_26845 = mux_26845(v_3627);
  assign v_26846 = mux_26846(v_3633);
  assign v_26847 = mux_26847(v_3606);
  assign v_26849 = v_26850 | v_26852;
  assign v_26850 = mux_26850(v_26851);
  assign v_26851 = ~act_3526;
  assign v_26852 = v_26853 | v_26861;
  assign v_26853 = mux_26853(v_3527);
  assign v_26855 = v_26856 | v_26858;
  assign v_26856 = mux_26856(v_26857);
  assign v_26857 = ~act_3570;
  assign v_26858 = v_26859 | v_26860;
  assign v_26859 = mux_26859(v_3571);
  assign v_26860 = mux_26860(v_3577);
  assign v_26861 = mux_26861(v_3557);
  assign v_26863 = v_26864 | v_26866;
  assign v_26864 = mux_26864(v_26865);
  assign v_26865 = ~act_3533;
  assign v_26866 = v_26867 | v_26868;
  assign v_26867 = mux_26867(v_3534);
  assign v_26868 = mux_26868(v_3540);
  assign v_26869 = mux_26869(v_3492);
  assign v_26871 = v_26872 | v_26874;
  assign v_26872 = mux_26872(v_26873);
  assign v_26873 = ~act_2628;
  assign v_26874 = v_26875 | v_26981;
  assign v_26875 = mux_26875(v_2629);
  assign v_26877 = v_26878 | v_26880;
  assign v_26878 = mux_26878(v_26879);
  assign v_26879 = ~act_3064;
  assign v_26880 = v_26881 | v_26931;
  assign v_26881 = mux_26881(v_3065);
  assign v_26883 = v_26884 | v_26886;
  assign v_26884 = mux_26884(v_26885);
  assign v_26885 = ~act_3276;
  assign v_26886 = v_26887 | v_26909;
  assign v_26887 = mux_26887(v_3277);
  assign v_26889 = v_26890 | v_26892;
  assign v_26890 = mux_26890(v_26891);
  assign v_26891 = ~act_3376;
  assign v_26892 = v_26893 | v_26901;
  assign v_26893 = mux_26893(v_3377);
  assign v_26895 = v_26896 | v_26898;
  assign v_26896 = mux_26896(v_26897);
  assign v_26897 = ~act_3420;
  assign v_26898 = v_26899 | v_26900;
  assign v_26899 = mux_26899(v_3421);
  assign v_26900 = mux_26900(v_3427);
  assign v_26901 = mux_26901(v_3407);
  assign v_26903 = v_26904 | v_26906;
  assign v_26904 = mux_26904(v_26905);
  assign v_26905 = ~act_3383;
  assign v_26906 = v_26907 | v_26908;
  assign v_26907 = mux_26907(v_3384);
  assign v_26908 = mux_26908(v_3390);
  assign v_26909 = mux_26909(v_3363);
  assign v_26911 = v_26912 | v_26914;
  assign v_26912 = mux_26912(v_26913);
  assign v_26913 = ~act_3283;
  assign v_26914 = v_26915 | v_26923;
  assign v_26915 = mux_26915(v_3284);
  assign v_26917 = v_26918 | v_26920;
  assign v_26918 = mux_26918(v_26919);
  assign v_26919 = ~act_3327;
  assign v_26920 = v_26921 | v_26922;
  assign v_26921 = mux_26921(v_3328);
  assign v_26922 = mux_26922(v_3334);
  assign v_26923 = mux_26923(v_3314);
  assign v_26925 = v_26926 | v_26928;
  assign v_26926 = mux_26926(v_26927);
  assign v_26927 = ~act_3290;
  assign v_26928 = v_26929 | v_26930;
  assign v_26929 = mux_26929(v_3291);
  assign v_26930 = mux_26930(v_3297);
  assign v_26931 = mux_26931(v_3263);
  assign v_26933 = v_26934 | v_26936;
  assign v_26934 = mux_26934(v_26935);
  assign v_26935 = ~act_3071;
  assign v_26936 = v_26937 | v_26959;
  assign v_26937 = mux_26937(v_3072);
  assign v_26939 = v_26940 | v_26942;
  assign v_26940 = mux_26940(v_26941);
  assign v_26941 = ~act_3171;
  assign v_26942 = v_26943 | v_26951;
  assign v_26943 = mux_26943(v_3172);
  assign v_26945 = v_26946 | v_26948;
  assign v_26946 = mux_26946(v_26947);
  assign v_26947 = ~act_3215;
  assign v_26948 = v_26949 | v_26950;
  assign v_26949 = mux_26949(v_3216);
  assign v_26950 = mux_26950(v_3222);
  assign v_26951 = mux_26951(v_3202);
  assign v_26953 = v_26954 | v_26956;
  assign v_26954 = mux_26954(v_26955);
  assign v_26955 = ~act_3178;
  assign v_26956 = v_26957 | v_26958;
  assign v_26957 = mux_26957(v_3179);
  assign v_26958 = mux_26958(v_3185);
  assign v_26959 = mux_26959(v_3158);
  assign v_26961 = v_26962 | v_26964;
  assign v_26962 = mux_26962(v_26963);
  assign v_26963 = ~act_3078;
  assign v_26964 = v_26965 | v_26973;
  assign v_26965 = mux_26965(v_3079);
  assign v_26967 = v_26968 | v_26970;
  assign v_26968 = mux_26968(v_26969);
  assign v_26969 = ~act_3122;
  assign v_26970 = v_26971 | v_26972;
  assign v_26971 = mux_26971(v_3123);
  assign v_26972 = mux_26972(v_3129);
  assign v_26973 = mux_26973(v_3109);
  assign v_26975 = v_26976 | v_26978;
  assign v_26976 = mux_26976(v_26977);
  assign v_26977 = ~act_3085;
  assign v_26978 = v_26979 | v_26980;
  assign v_26979 = mux_26979(v_3086);
  assign v_26980 = mux_26980(v_3092);
  assign v_26981 = mux_26981(v_3051);
  assign v_26983 = v_26984 | v_26986;
  assign v_26984 = mux_26984(v_26985);
  assign v_26985 = ~act_2635;
  assign v_26986 = v_26987 | v_27037;
  assign v_26987 = mux_26987(v_2636);
  assign v_26989 = v_26990 | v_26992;
  assign v_26990 = mux_26990(v_26991);
  assign v_26991 = ~act_2847;
  assign v_26992 = v_26993 | v_27015;
  assign v_26993 = mux_26993(v_2848);
  assign v_26995 = v_26996 | v_26998;
  assign v_26996 = mux_26996(v_26997);
  assign v_26997 = ~act_2947;
  assign v_26998 = v_26999 | v_27007;
  assign v_26999 = mux_26999(v_2948);
  assign v_27001 = v_27002 | v_27004;
  assign v_27002 = mux_27002(v_27003);
  assign v_27003 = ~act_2991;
  assign v_27004 = v_27005 | v_27006;
  assign v_27005 = mux_27005(v_2992);
  assign v_27006 = mux_27006(v_2998);
  assign v_27007 = mux_27007(v_2978);
  assign v_27009 = v_27010 | v_27012;
  assign v_27010 = mux_27010(v_27011);
  assign v_27011 = ~act_2954;
  assign v_27012 = v_27013 | v_27014;
  assign v_27013 = mux_27013(v_2955);
  assign v_27014 = mux_27014(v_2961);
  assign v_27015 = mux_27015(v_2934);
  assign v_27017 = v_27018 | v_27020;
  assign v_27018 = mux_27018(v_27019);
  assign v_27019 = ~act_2854;
  assign v_27020 = v_27021 | v_27029;
  assign v_27021 = mux_27021(v_2855);
  assign v_27023 = v_27024 | v_27026;
  assign v_27024 = mux_27024(v_27025);
  assign v_27025 = ~act_2898;
  assign v_27026 = v_27027 | v_27028;
  assign v_27027 = mux_27027(v_2899);
  assign v_27028 = mux_27028(v_2905);
  assign v_27029 = mux_27029(v_2885);
  assign v_27031 = v_27032 | v_27034;
  assign v_27032 = mux_27032(v_27033);
  assign v_27033 = ~act_2861;
  assign v_27034 = v_27035 | v_27036;
  assign v_27035 = mux_27035(v_2862);
  assign v_27036 = mux_27036(v_2868);
  assign v_27037 = mux_27037(v_2834);
  assign v_27039 = v_27040 | v_27042;
  assign v_27040 = mux_27040(v_27041);
  assign v_27041 = ~act_2642;
  assign v_27042 = v_27043 | v_27065;
  assign v_27043 = mux_27043(v_2643);
  assign v_27045 = v_27046 | v_27048;
  assign v_27046 = mux_27046(v_27047);
  assign v_27047 = ~act_2742;
  assign v_27048 = v_27049 | v_27057;
  assign v_27049 = mux_27049(v_2743);
  assign v_27051 = v_27052 | v_27054;
  assign v_27052 = mux_27052(v_27053);
  assign v_27053 = ~act_2786;
  assign v_27054 = v_27055 | v_27056;
  assign v_27055 = mux_27055(v_2787);
  assign v_27056 = mux_27056(v_2793);
  assign v_27057 = mux_27057(v_2773);
  assign v_27059 = v_27060 | v_27062;
  assign v_27060 = mux_27060(v_27061);
  assign v_27061 = ~act_2749;
  assign v_27062 = v_27063 | v_27064;
  assign v_27063 = mux_27063(v_2750);
  assign v_27064 = mux_27064(v_2756);
  assign v_27065 = mux_27065(v_2729);
  assign v_27067 = v_27068 | v_27070;
  assign v_27068 = mux_27068(v_27069);
  assign v_27069 = ~act_2649;
  assign v_27070 = v_27071 | v_27079;
  assign v_27071 = mux_27071(v_2650);
  assign v_27073 = v_27074 | v_27076;
  assign v_27074 = mux_27074(v_27075);
  assign v_27075 = ~act_2693;
  assign v_27076 = v_27077 | v_27078;
  assign v_27077 = mux_27077(v_2694);
  assign v_27078 = mux_27078(v_2700);
  assign v_27079 = mux_27079(v_2680);
  assign v_27081 = v_27082 | v_27084;
  assign v_27082 = mux_27082(v_27083);
  assign v_27083 = ~act_2656;
  assign v_27084 = v_27085 | v_27086;
  assign v_27085 = mux_27085(v_2657);
  assign v_27086 = mux_27086(v_2663);
  assign v_27087 = mux_27087(v_7953);
  assign v_27089 = v_27090 | v_27092;
  assign v_27090 = mux_27090(v_27091);
  assign v_27091 = ~act_4401;
  assign v_27092 = v_27093 | v_27535;
  assign v_27093 = mux_27093(v_4402);
  assign v_27095 = v_27096 | v_27098;
  assign v_27096 = mux_27096(v_27097);
  assign v_27097 = ~act_6181;
  assign v_27098 = v_27099 | v_27317;
  assign v_27099 = mux_27099(v_6182);
  assign v_27101 = v_27102 | v_27104;
  assign v_27102 = mux_27102(v_27103);
  assign v_27103 = ~act_7065;
  assign v_27104 = v_27105 | v_27211;
  assign v_27105 = mux_27105(v_7066);
  assign v_27107 = v_27108 | v_27110;
  assign v_27108 = mux_27108(v_27109);
  assign v_27109 = ~act_7501;
  assign v_27110 = v_27111 | v_27161;
  assign v_27111 = mux_27111(v_7502);
  assign v_27113 = v_27114 | v_27116;
  assign v_27114 = mux_27114(v_27115);
  assign v_27115 = ~act_7713;
  assign v_27116 = v_27117 | v_27139;
  assign v_27117 = mux_27117(v_7714);
  assign v_27119 = v_27120 | v_27122;
  assign v_27120 = mux_27120(v_27121);
  assign v_27121 = ~act_7813;
  assign v_27122 = v_27123 | v_27131;
  assign v_27123 = mux_27123(v_7814);
  assign v_27125 = v_27126 | v_27128;
  assign v_27126 = mux_27126(v_27127);
  assign v_27127 = ~act_7857;
  assign v_27128 = v_27129 | v_27130;
  assign v_27129 = mux_27129(v_7858);
  assign v_27130 = mux_27130(v_7864);
  assign v_27131 = mux_27131(v_7844);
  assign v_27133 = v_27134 | v_27136;
  assign v_27134 = mux_27134(v_27135);
  assign v_27135 = ~act_7820;
  assign v_27136 = v_27137 | v_27138;
  assign v_27137 = mux_27137(v_7821);
  assign v_27138 = mux_27138(v_7827);
  assign v_27139 = mux_27139(v_7800);
  assign v_27141 = v_27142 | v_27144;
  assign v_27142 = mux_27142(v_27143);
  assign v_27143 = ~act_7720;
  assign v_27144 = v_27145 | v_27153;
  assign v_27145 = mux_27145(v_7721);
  assign v_27147 = v_27148 | v_27150;
  assign v_27148 = mux_27148(v_27149);
  assign v_27149 = ~act_7764;
  assign v_27150 = v_27151 | v_27152;
  assign v_27151 = mux_27151(v_7765);
  assign v_27152 = mux_27152(v_7771);
  assign v_27153 = mux_27153(v_7751);
  assign v_27155 = v_27156 | v_27158;
  assign v_27156 = mux_27156(v_27157);
  assign v_27157 = ~act_7727;
  assign v_27158 = v_27159 | v_27160;
  assign v_27159 = mux_27159(v_7728);
  assign v_27160 = mux_27160(v_7734);
  assign v_27161 = mux_27161(v_7700);
  assign v_27163 = v_27164 | v_27166;
  assign v_27164 = mux_27164(v_27165);
  assign v_27165 = ~act_7508;
  assign v_27166 = v_27167 | v_27189;
  assign v_27167 = mux_27167(v_7509);
  assign v_27169 = v_27170 | v_27172;
  assign v_27170 = mux_27170(v_27171);
  assign v_27171 = ~act_7608;
  assign v_27172 = v_27173 | v_27181;
  assign v_27173 = mux_27173(v_7609);
  assign v_27175 = v_27176 | v_27178;
  assign v_27176 = mux_27176(v_27177);
  assign v_27177 = ~act_7652;
  assign v_27178 = v_27179 | v_27180;
  assign v_27179 = mux_27179(v_7653);
  assign v_27180 = mux_27180(v_7659);
  assign v_27181 = mux_27181(v_7639);
  assign v_27183 = v_27184 | v_27186;
  assign v_27184 = mux_27184(v_27185);
  assign v_27185 = ~act_7615;
  assign v_27186 = v_27187 | v_27188;
  assign v_27187 = mux_27187(v_7616);
  assign v_27188 = mux_27188(v_7622);
  assign v_27189 = mux_27189(v_7595);
  assign v_27191 = v_27192 | v_27194;
  assign v_27192 = mux_27192(v_27193);
  assign v_27193 = ~act_7515;
  assign v_27194 = v_27195 | v_27203;
  assign v_27195 = mux_27195(v_7516);
  assign v_27197 = v_27198 | v_27200;
  assign v_27198 = mux_27198(v_27199);
  assign v_27199 = ~act_7559;
  assign v_27200 = v_27201 | v_27202;
  assign v_27201 = mux_27201(v_7560);
  assign v_27202 = mux_27202(v_7566);
  assign v_27203 = mux_27203(v_7546);
  assign v_27205 = v_27206 | v_27208;
  assign v_27206 = mux_27206(v_27207);
  assign v_27207 = ~act_7522;
  assign v_27208 = v_27209 | v_27210;
  assign v_27209 = mux_27209(v_7523);
  assign v_27210 = mux_27210(v_7529);
  assign v_27211 = mux_27211(v_7488);
  assign v_27213 = v_27214 | v_27216;
  assign v_27214 = mux_27214(v_27215);
  assign v_27215 = ~act_7072;
  assign v_27216 = v_27217 | v_27267;
  assign v_27217 = mux_27217(v_7073);
  assign v_27219 = v_27220 | v_27222;
  assign v_27220 = mux_27220(v_27221);
  assign v_27221 = ~act_7284;
  assign v_27222 = v_27223 | v_27245;
  assign v_27223 = mux_27223(v_7285);
  assign v_27225 = v_27226 | v_27228;
  assign v_27226 = mux_27226(v_27227);
  assign v_27227 = ~act_7384;
  assign v_27228 = v_27229 | v_27237;
  assign v_27229 = mux_27229(v_7385);
  assign v_27231 = v_27232 | v_27234;
  assign v_27232 = mux_27232(v_27233);
  assign v_27233 = ~act_7428;
  assign v_27234 = v_27235 | v_27236;
  assign v_27235 = mux_27235(v_7429);
  assign v_27236 = mux_27236(v_7435);
  assign v_27237 = mux_27237(v_7415);
  assign v_27239 = v_27240 | v_27242;
  assign v_27240 = mux_27240(v_27241);
  assign v_27241 = ~act_7391;
  assign v_27242 = v_27243 | v_27244;
  assign v_27243 = mux_27243(v_7392);
  assign v_27244 = mux_27244(v_7398);
  assign v_27245 = mux_27245(v_7371);
  assign v_27247 = v_27248 | v_27250;
  assign v_27248 = mux_27248(v_27249);
  assign v_27249 = ~act_7291;
  assign v_27250 = v_27251 | v_27259;
  assign v_27251 = mux_27251(v_7292);
  assign v_27253 = v_27254 | v_27256;
  assign v_27254 = mux_27254(v_27255);
  assign v_27255 = ~act_7335;
  assign v_27256 = v_27257 | v_27258;
  assign v_27257 = mux_27257(v_7336);
  assign v_27258 = mux_27258(v_7342);
  assign v_27259 = mux_27259(v_7322);
  assign v_27261 = v_27262 | v_27264;
  assign v_27262 = mux_27262(v_27263);
  assign v_27263 = ~act_7298;
  assign v_27264 = v_27265 | v_27266;
  assign v_27265 = mux_27265(v_7299);
  assign v_27266 = mux_27266(v_7305);
  assign v_27267 = mux_27267(v_7271);
  assign v_27269 = v_27270 | v_27272;
  assign v_27270 = mux_27270(v_27271);
  assign v_27271 = ~act_7079;
  assign v_27272 = v_27273 | v_27295;
  assign v_27273 = mux_27273(v_7080);
  assign v_27275 = v_27276 | v_27278;
  assign v_27276 = mux_27276(v_27277);
  assign v_27277 = ~act_7179;
  assign v_27278 = v_27279 | v_27287;
  assign v_27279 = mux_27279(v_7180);
  assign v_27281 = v_27282 | v_27284;
  assign v_27282 = mux_27282(v_27283);
  assign v_27283 = ~act_7223;
  assign v_27284 = v_27285 | v_27286;
  assign v_27285 = mux_27285(v_7224);
  assign v_27286 = mux_27286(v_7230);
  assign v_27287 = mux_27287(v_7210);
  assign v_27289 = v_27290 | v_27292;
  assign v_27290 = mux_27290(v_27291);
  assign v_27291 = ~act_7186;
  assign v_27292 = v_27293 | v_27294;
  assign v_27293 = mux_27293(v_7187);
  assign v_27294 = mux_27294(v_7193);
  assign v_27295 = mux_27295(v_7166);
  assign v_27297 = v_27298 | v_27300;
  assign v_27298 = mux_27298(v_27299);
  assign v_27299 = ~act_7086;
  assign v_27300 = v_27301 | v_27309;
  assign v_27301 = mux_27301(v_7087);
  assign v_27303 = v_27304 | v_27306;
  assign v_27304 = mux_27304(v_27305);
  assign v_27305 = ~act_7130;
  assign v_27306 = v_27307 | v_27308;
  assign v_27307 = mux_27307(v_7131);
  assign v_27308 = mux_27308(v_7137);
  assign v_27309 = mux_27309(v_7117);
  assign v_27311 = v_27312 | v_27314;
  assign v_27312 = mux_27312(v_27313);
  assign v_27313 = ~act_7093;
  assign v_27314 = v_27315 | v_27316;
  assign v_27315 = mux_27315(v_7094);
  assign v_27316 = mux_27316(v_7100);
  assign v_27317 = mux_27317(v_7052);
  assign v_27319 = v_27320 | v_27322;
  assign v_27320 = mux_27320(v_27321);
  assign v_27321 = ~act_6188;
  assign v_27322 = v_27323 | v_27429;
  assign v_27323 = mux_27323(v_6189);
  assign v_27325 = v_27326 | v_27328;
  assign v_27326 = mux_27326(v_27327);
  assign v_27327 = ~act_6624;
  assign v_27328 = v_27329 | v_27379;
  assign v_27329 = mux_27329(v_6625);
  assign v_27331 = v_27332 | v_27334;
  assign v_27332 = mux_27332(v_27333);
  assign v_27333 = ~act_6836;
  assign v_27334 = v_27335 | v_27357;
  assign v_27335 = mux_27335(v_6837);
  assign v_27337 = v_27338 | v_27340;
  assign v_27338 = mux_27338(v_27339);
  assign v_27339 = ~act_6936;
  assign v_27340 = v_27341 | v_27349;
  assign v_27341 = mux_27341(v_6937);
  assign v_27343 = v_27344 | v_27346;
  assign v_27344 = mux_27344(v_27345);
  assign v_27345 = ~act_6980;
  assign v_27346 = v_27347 | v_27348;
  assign v_27347 = mux_27347(v_6981);
  assign v_27348 = mux_27348(v_6987);
  assign v_27349 = mux_27349(v_6967);
  assign v_27351 = v_27352 | v_27354;
  assign v_27352 = mux_27352(v_27353);
  assign v_27353 = ~act_6943;
  assign v_27354 = v_27355 | v_27356;
  assign v_27355 = mux_27355(v_6944);
  assign v_27356 = mux_27356(v_6950);
  assign v_27357 = mux_27357(v_6923);
  assign v_27359 = v_27360 | v_27362;
  assign v_27360 = mux_27360(v_27361);
  assign v_27361 = ~act_6843;
  assign v_27362 = v_27363 | v_27371;
  assign v_27363 = mux_27363(v_6844);
  assign v_27365 = v_27366 | v_27368;
  assign v_27366 = mux_27366(v_27367);
  assign v_27367 = ~act_6887;
  assign v_27368 = v_27369 | v_27370;
  assign v_27369 = mux_27369(v_6888);
  assign v_27370 = mux_27370(v_6894);
  assign v_27371 = mux_27371(v_6874);
  assign v_27373 = v_27374 | v_27376;
  assign v_27374 = mux_27374(v_27375);
  assign v_27375 = ~act_6850;
  assign v_27376 = v_27377 | v_27378;
  assign v_27377 = mux_27377(v_6851);
  assign v_27378 = mux_27378(v_6857);
  assign v_27379 = mux_27379(v_6823);
  assign v_27381 = v_27382 | v_27384;
  assign v_27382 = mux_27382(v_27383);
  assign v_27383 = ~act_6631;
  assign v_27384 = v_27385 | v_27407;
  assign v_27385 = mux_27385(v_6632);
  assign v_27387 = v_27388 | v_27390;
  assign v_27388 = mux_27388(v_27389);
  assign v_27389 = ~act_6731;
  assign v_27390 = v_27391 | v_27399;
  assign v_27391 = mux_27391(v_6732);
  assign v_27393 = v_27394 | v_27396;
  assign v_27394 = mux_27394(v_27395);
  assign v_27395 = ~act_6775;
  assign v_27396 = v_27397 | v_27398;
  assign v_27397 = mux_27397(v_6776);
  assign v_27398 = mux_27398(v_6782);
  assign v_27399 = mux_27399(v_6762);
  assign v_27401 = v_27402 | v_27404;
  assign v_27402 = mux_27402(v_27403);
  assign v_27403 = ~act_6738;
  assign v_27404 = v_27405 | v_27406;
  assign v_27405 = mux_27405(v_6739);
  assign v_27406 = mux_27406(v_6745);
  assign v_27407 = mux_27407(v_6718);
  assign v_27409 = v_27410 | v_27412;
  assign v_27410 = mux_27410(v_27411);
  assign v_27411 = ~act_6638;
  assign v_27412 = v_27413 | v_27421;
  assign v_27413 = mux_27413(v_6639);
  assign v_27415 = v_27416 | v_27418;
  assign v_27416 = mux_27416(v_27417);
  assign v_27417 = ~act_6682;
  assign v_27418 = v_27419 | v_27420;
  assign v_27419 = mux_27419(v_6683);
  assign v_27420 = mux_27420(v_6689);
  assign v_27421 = mux_27421(v_6669);
  assign v_27423 = v_27424 | v_27426;
  assign v_27424 = mux_27424(v_27425);
  assign v_27425 = ~act_6645;
  assign v_27426 = v_27427 | v_27428;
  assign v_27427 = mux_27427(v_6646);
  assign v_27428 = mux_27428(v_6652);
  assign v_27429 = mux_27429(v_6611);
  assign v_27431 = v_27432 | v_27434;
  assign v_27432 = mux_27432(v_27433);
  assign v_27433 = ~act_6195;
  assign v_27434 = v_27435 | v_27485;
  assign v_27435 = mux_27435(v_6196);
  assign v_27437 = v_27438 | v_27440;
  assign v_27438 = mux_27438(v_27439);
  assign v_27439 = ~act_6407;
  assign v_27440 = v_27441 | v_27463;
  assign v_27441 = mux_27441(v_6408);
  assign v_27443 = v_27444 | v_27446;
  assign v_27444 = mux_27444(v_27445);
  assign v_27445 = ~act_6507;
  assign v_27446 = v_27447 | v_27455;
  assign v_27447 = mux_27447(v_6508);
  assign v_27449 = v_27450 | v_27452;
  assign v_27450 = mux_27450(v_27451);
  assign v_27451 = ~act_6551;
  assign v_27452 = v_27453 | v_27454;
  assign v_27453 = mux_27453(v_6552);
  assign v_27454 = mux_27454(v_6558);
  assign v_27455 = mux_27455(v_6538);
  assign v_27457 = v_27458 | v_27460;
  assign v_27458 = mux_27458(v_27459);
  assign v_27459 = ~act_6514;
  assign v_27460 = v_27461 | v_27462;
  assign v_27461 = mux_27461(v_6515);
  assign v_27462 = mux_27462(v_6521);
  assign v_27463 = mux_27463(v_6494);
  assign v_27465 = v_27466 | v_27468;
  assign v_27466 = mux_27466(v_27467);
  assign v_27467 = ~act_6414;
  assign v_27468 = v_27469 | v_27477;
  assign v_27469 = mux_27469(v_6415);
  assign v_27471 = v_27472 | v_27474;
  assign v_27472 = mux_27472(v_27473);
  assign v_27473 = ~act_6458;
  assign v_27474 = v_27475 | v_27476;
  assign v_27475 = mux_27475(v_6459);
  assign v_27476 = mux_27476(v_6465);
  assign v_27477 = mux_27477(v_6445);
  assign v_27479 = v_27480 | v_27482;
  assign v_27480 = mux_27480(v_27481);
  assign v_27481 = ~act_6421;
  assign v_27482 = v_27483 | v_27484;
  assign v_27483 = mux_27483(v_6422);
  assign v_27484 = mux_27484(v_6428);
  assign v_27485 = mux_27485(v_6394);
  assign v_27487 = v_27488 | v_27490;
  assign v_27488 = mux_27488(v_27489);
  assign v_27489 = ~act_6202;
  assign v_27490 = v_27491 | v_27513;
  assign v_27491 = mux_27491(v_6203);
  assign v_27493 = v_27494 | v_27496;
  assign v_27494 = mux_27494(v_27495);
  assign v_27495 = ~act_6302;
  assign v_27496 = v_27497 | v_27505;
  assign v_27497 = mux_27497(v_6303);
  assign v_27499 = v_27500 | v_27502;
  assign v_27500 = mux_27500(v_27501);
  assign v_27501 = ~act_6346;
  assign v_27502 = v_27503 | v_27504;
  assign v_27503 = mux_27503(v_6347);
  assign v_27504 = mux_27504(v_6353);
  assign v_27505 = mux_27505(v_6333);
  assign v_27507 = v_27508 | v_27510;
  assign v_27508 = mux_27508(v_27509);
  assign v_27509 = ~act_6309;
  assign v_27510 = v_27511 | v_27512;
  assign v_27511 = mux_27511(v_6310);
  assign v_27512 = mux_27512(v_6316);
  assign v_27513 = mux_27513(v_6289);
  assign v_27515 = v_27516 | v_27518;
  assign v_27516 = mux_27516(v_27517);
  assign v_27517 = ~act_6209;
  assign v_27518 = v_27519 | v_27527;
  assign v_27519 = mux_27519(v_6210);
  assign v_27521 = v_27522 | v_27524;
  assign v_27522 = mux_27522(v_27523);
  assign v_27523 = ~act_6253;
  assign v_27524 = v_27525 | v_27526;
  assign v_27525 = mux_27525(v_6254);
  assign v_27526 = mux_27526(v_6260);
  assign v_27527 = mux_27527(v_6240);
  assign v_27529 = v_27530 | v_27532;
  assign v_27530 = mux_27530(v_27531);
  assign v_27531 = ~act_6216;
  assign v_27532 = v_27533 | v_27534;
  assign v_27533 = mux_27533(v_6217);
  assign v_27534 = mux_27534(v_6223);
  assign v_27535 = mux_27535(v_6168);
  assign v_27537 = v_27538 | v_27540;
  assign v_27538 = mux_27538(v_27539);
  assign v_27539 = ~act_4408;
  assign v_27540 = v_27541 | v_27759;
  assign v_27541 = mux_27541(v_4409);
  assign v_27543 = v_27544 | v_27546;
  assign v_27544 = mux_27544(v_27545);
  assign v_27545 = ~act_5292;
  assign v_27546 = v_27547 | v_27653;
  assign v_27547 = mux_27547(v_5293);
  assign v_27549 = v_27550 | v_27552;
  assign v_27550 = mux_27550(v_27551);
  assign v_27551 = ~act_5728;
  assign v_27552 = v_27553 | v_27603;
  assign v_27553 = mux_27553(v_5729);
  assign v_27555 = v_27556 | v_27558;
  assign v_27556 = mux_27556(v_27557);
  assign v_27557 = ~act_5940;
  assign v_27558 = v_27559 | v_27581;
  assign v_27559 = mux_27559(v_5941);
  assign v_27561 = v_27562 | v_27564;
  assign v_27562 = mux_27562(v_27563);
  assign v_27563 = ~act_6040;
  assign v_27564 = v_27565 | v_27573;
  assign v_27565 = mux_27565(v_6041);
  assign v_27567 = v_27568 | v_27570;
  assign v_27568 = mux_27568(v_27569);
  assign v_27569 = ~act_6084;
  assign v_27570 = v_27571 | v_27572;
  assign v_27571 = mux_27571(v_6085);
  assign v_27572 = mux_27572(v_6091);
  assign v_27573 = mux_27573(v_6071);
  assign v_27575 = v_27576 | v_27578;
  assign v_27576 = mux_27576(v_27577);
  assign v_27577 = ~act_6047;
  assign v_27578 = v_27579 | v_27580;
  assign v_27579 = mux_27579(v_6048);
  assign v_27580 = mux_27580(v_6054);
  assign v_27581 = mux_27581(v_6027);
  assign v_27583 = v_27584 | v_27586;
  assign v_27584 = mux_27584(v_27585);
  assign v_27585 = ~act_5947;
  assign v_27586 = v_27587 | v_27595;
  assign v_27587 = mux_27587(v_5948);
  assign v_27589 = v_27590 | v_27592;
  assign v_27590 = mux_27590(v_27591);
  assign v_27591 = ~act_5991;
  assign v_27592 = v_27593 | v_27594;
  assign v_27593 = mux_27593(v_5992);
  assign v_27594 = mux_27594(v_5998);
  assign v_27595 = mux_27595(v_5978);
  assign v_27597 = v_27598 | v_27600;
  assign v_27598 = mux_27598(v_27599);
  assign v_27599 = ~act_5954;
  assign v_27600 = v_27601 | v_27602;
  assign v_27601 = mux_27601(v_5955);
  assign v_27602 = mux_27602(v_5961);
  assign v_27603 = mux_27603(v_5927);
  assign v_27605 = v_27606 | v_27608;
  assign v_27606 = mux_27606(v_27607);
  assign v_27607 = ~act_5735;
  assign v_27608 = v_27609 | v_27631;
  assign v_27609 = mux_27609(v_5736);
  assign v_27611 = v_27612 | v_27614;
  assign v_27612 = mux_27612(v_27613);
  assign v_27613 = ~act_5835;
  assign v_27614 = v_27615 | v_27623;
  assign v_27615 = mux_27615(v_5836);
  assign v_27617 = v_27618 | v_27620;
  assign v_27618 = mux_27618(v_27619);
  assign v_27619 = ~act_5879;
  assign v_27620 = v_27621 | v_27622;
  assign v_27621 = mux_27621(v_5880);
  assign v_27622 = mux_27622(v_5886);
  assign v_27623 = mux_27623(v_5866);
  assign v_27625 = v_27626 | v_27628;
  assign v_27626 = mux_27626(v_27627);
  assign v_27627 = ~act_5842;
  assign v_27628 = v_27629 | v_27630;
  assign v_27629 = mux_27629(v_5843);
  assign v_27630 = mux_27630(v_5849);
  assign v_27631 = mux_27631(v_5822);
  assign v_27633 = v_27634 | v_27636;
  assign v_27634 = mux_27634(v_27635);
  assign v_27635 = ~act_5742;
  assign v_27636 = v_27637 | v_27645;
  assign v_27637 = mux_27637(v_5743);
  assign v_27639 = v_27640 | v_27642;
  assign v_27640 = mux_27640(v_27641);
  assign v_27641 = ~act_5786;
  assign v_27642 = v_27643 | v_27644;
  assign v_27643 = mux_27643(v_5787);
  assign v_27644 = mux_27644(v_5793);
  assign v_27645 = mux_27645(v_5773);
  assign v_27647 = v_27648 | v_27650;
  assign v_27648 = mux_27648(v_27649);
  assign v_27649 = ~act_5749;
  assign v_27650 = v_27651 | v_27652;
  assign v_27651 = mux_27651(v_5750);
  assign v_27652 = mux_27652(v_5756);
  assign v_27653 = mux_27653(v_5715);
  assign v_27655 = v_27656 | v_27658;
  assign v_27656 = mux_27656(v_27657);
  assign v_27657 = ~act_5299;
  assign v_27658 = v_27659 | v_27709;
  assign v_27659 = mux_27659(v_5300);
  assign v_27661 = v_27662 | v_27664;
  assign v_27662 = mux_27662(v_27663);
  assign v_27663 = ~act_5511;
  assign v_27664 = v_27665 | v_27687;
  assign v_27665 = mux_27665(v_5512);
  assign v_27667 = v_27668 | v_27670;
  assign v_27668 = mux_27668(v_27669);
  assign v_27669 = ~act_5611;
  assign v_27670 = v_27671 | v_27679;
  assign v_27671 = mux_27671(v_5612);
  assign v_27673 = v_27674 | v_27676;
  assign v_27674 = mux_27674(v_27675);
  assign v_27675 = ~act_5655;
  assign v_27676 = v_27677 | v_27678;
  assign v_27677 = mux_27677(v_5656);
  assign v_27678 = mux_27678(v_5662);
  assign v_27679 = mux_27679(v_5642);
  assign v_27681 = v_27682 | v_27684;
  assign v_27682 = mux_27682(v_27683);
  assign v_27683 = ~act_5618;
  assign v_27684 = v_27685 | v_27686;
  assign v_27685 = mux_27685(v_5619);
  assign v_27686 = mux_27686(v_5625);
  assign v_27687 = mux_27687(v_5598);
  assign v_27689 = v_27690 | v_27692;
  assign v_27690 = mux_27690(v_27691);
  assign v_27691 = ~act_5518;
  assign v_27692 = v_27693 | v_27701;
  assign v_27693 = mux_27693(v_5519);
  assign v_27695 = v_27696 | v_27698;
  assign v_27696 = mux_27696(v_27697);
  assign v_27697 = ~act_5562;
  assign v_27698 = v_27699 | v_27700;
  assign v_27699 = mux_27699(v_5563);
  assign v_27700 = mux_27700(v_5569);
  assign v_27701 = mux_27701(v_5549);
  assign v_27703 = v_27704 | v_27706;
  assign v_27704 = mux_27704(v_27705);
  assign v_27705 = ~act_5525;
  assign v_27706 = v_27707 | v_27708;
  assign v_27707 = mux_27707(v_5526);
  assign v_27708 = mux_27708(v_5532);
  assign v_27709 = mux_27709(v_5498);
  assign v_27711 = v_27712 | v_27714;
  assign v_27712 = mux_27712(v_27713);
  assign v_27713 = ~act_5306;
  assign v_27714 = v_27715 | v_27737;
  assign v_27715 = mux_27715(v_5307);
  assign v_27717 = v_27718 | v_27720;
  assign v_27718 = mux_27718(v_27719);
  assign v_27719 = ~act_5406;
  assign v_27720 = v_27721 | v_27729;
  assign v_27721 = mux_27721(v_5407);
  assign v_27723 = v_27724 | v_27726;
  assign v_27724 = mux_27724(v_27725);
  assign v_27725 = ~act_5450;
  assign v_27726 = v_27727 | v_27728;
  assign v_27727 = mux_27727(v_5451);
  assign v_27728 = mux_27728(v_5457);
  assign v_27729 = mux_27729(v_5437);
  assign v_27731 = v_27732 | v_27734;
  assign v_27732 = mux_27732(v_27733);
  assign v_27733 = ~act_5413;
  assign v_27734 = v_27735 | v_27736;
  assign v_27735 = mux_27735(v_5414);
  assign v_27736 = mux_27736(v_5420);
  assign v_27737 = mux_27737(v_5393);
  assign v_27739 = v_27740 | v_27742;
  assign v_27740 = mux_27740(v_27741);
  assign v_27741 = ~act_5313;
  assign v_27742 = v_27743 | v_27751;
  assign v_27743 = mux_27743(v_5314);
  assign v_27745 = v_27746 | v_27748;
  assign v_27746 = mux_27746(v_27747);
  assign v_27747 = ~act_5357;
  assign v_27748 = v_27749 | v_27750;
  assign v_27749 = mux_27749(v_5358);
  assign v_27750 = mux_27750(v_5364);
  assign v_27751 = mux_27751(v_5344);
  assign v_27753 = v_27754 | v_27756;
  assign v_27754 = mux_27754(v_27755);
  assign v_27755 = ~act_5320;
  assign v_27756 = v_27757 | v_27758;
  assign v_27757 = mux_27757(v_5321);
  assign v_27758 = mux_27758(v_5327);
  assign v_27759 = mux_27759(v_5279);
  assign v_27761 = v_27762 | v_27764;
  assign v_27762 = mux_27762(v_27763);
  assign v_27763 = ~act_4415;
  assign v_27764 = v_27765 | v_27871;
  assign v_27765 = mux_27765(v_4416);
  assign v_27767 = v_27768 | v_27770;
  assign v_27768 = mux_27768(v_27769);
  assign v_27769 = ~act_4851;
  assign v_27770 = v_27771 | v_27821;
  assign v_27771 = mux_27771(v_4852);
  assign v_27773 = v_27774 | v_27776;
  assign v_27774 = mux_27774(v_27775);
  assign v_27775 = ~act_5063;
  assign v_27776 = v_27777 | v_27799;
  assign v_27777 = mux_27777(v_5064);
  assign v_27779 = v_27780 | v_27782;
  assign v_27780 = mux_27780(v_27781);
  assign v_27781 = ~act_5163;
  assign v_27782 = v_27783 | v_27791;
  assign v_27783 = mux_27783(v_5164);
  assign v_27785 = v_27786 | v_27788;
  assign v_27786 = mux_27786(v_27787);
  assign v_27787 = ~act_5207;
  assign v_27788 = v_27789 | v_27790;
  assign v_27789 = mux_27789(v_5208);
  assign v_27790 = mux_27790(v_5214);
  assign v_27791 = mux_27791(v_5194);
  assign v_27793 = v_27794 | v_27796;
  assign v_27794 = mux_27794(v_27795);
  assign v_27795 = ~act_5170;
  assign v_27796 = v_27797 | v_27798;
  assign v_27797 = mux_27797(v_5171);
  assign v_27798 = mux_27798(v_5177);
  assign v_27799 = mux_27799(v_5150);
  assign v_27801 = v_27802 | v_27804;
  assign v_27802 = mux_27802(v_27803);
  assign v_27803 = ~act_5070;
  assign v_27804 = v_27805 | v_27813;
  assign v_27805 = mux_27805(v_5071);
  assign v_27807 = v_27808 | v_27810;
  assign v_27808 = mux_27808(v_27809);
  assign v_27809 = ~act_5114;
  assign v_27810 = v_27811 | v_27812;
  assign v_27811 = mux_27811(v_5115);
  assign v_27812 = mux_27812(v_5121);
  assign v_27813 = mux_27813(v_5101);
  assign v_27815 = v_27816 | v_27818;
  assign v_27816 = mux_27816(v_27817);
  assign v_27817 = ~act_5077;
  assign v_27818 = v_27819 | v_27820;
  assign v_27819 = mux_27819(v_5078);
  assign v_27820 = mux_27820(v_5084);
  assign v_27821 = mux_27821(v_5050);
  assign v_27823 = v_27824 | v_27826;
  assign v_27824 = mux_27824(v_27825);
  assign v_27825 = ~act_4858;
  assign v_27826 = v_27827 | v_27849;
  assign v_27827 = mux_27827(v_4859);
  assign v_27829 = v_27830 | v_27832;
  assign v_27830 = mux_27830(v_27831);
  assign v_27831 = ~act_4958;
  assign v_27832 = v_27833 | v_27841;
  assign v_27833 = mux_27833(v_4959);
  assign v_27835 = v_27836 | v_27838;
  assign v_27836 = mux_27836(v_27837);
  assign v_27837 = ~act_5002;
  assign v_27838 = v_27839 | v_27840;
  assign v_27839 = mux_27839(v_5003);
  assign v_27840 = mux_27840(v_5009);
  assign v_27841 = mux_27841(v_4989);
  assign v_27843 = v_27844 | v_27846;
  assign v_27844 = mux_27844(v_27845);
  assign v_27845 = ~act_4965;
  assign v_27846 = v_27847 | v_27848;
  assign v_27847 = mux_27847(v_4966);
  assign v_27848 = mux_27848(v_4972);
  assign v_27849 = mux_27849(v_4945);
  assign v_27851 = v_27852 | v_27854;
  assign v_27852 = mux_27852(v_27853);
  assign v_27853 = ~act_4865;
  assign v_27854 = v_27855 | v_27863;
  assign v_27855 = mux_27855(v_4866);
  assign v_27857 = v_27858 | v_27860;
  assign v_27858 = mux_27858(v_27859);
  assign v_27859 = ~act_4909;
  assign v_27860 = v_27861 | v_27862;
  assign v_27861 = mux_27861(v_4910);
  assign v_27862 = mux_27862(v_4916);
  assign v_27863 = mux_27863(v_4896);
  assign v_27865 = v_27866 | v_27868;
  assign v_27866 = mux_27866(v_27867);
  assign v_27867 = ~act_4872;
  assign v_27868 = v_27869 | v_27870;
  assign v_27869 = mux_27869(v_4873);
  assign v_27870 = mux_27870(v_4879);
  assign v_27871 = mux_27871(v_4838);
  assign v_27873 = v_27874 | v_27876;
  assign v_27874 = mux_27874(v_27875);
  assign v_27875 = ~act_4422;
  assign v_27876 = v_27877 | v_27927;
  assign v_27877 = mux_27877(v_4423);
  assign v_27879 = v_27880 | v_27882;
  assign v_27880 = mux_27880(v_27881);
  assign v_27881 = ~act_4634;
  assign v_27882 = v_27883 | v_27905;
  assign v_27883 = mux_27883(v_4635);
  assign v_27885 = v_27886 | v_27888;
  assign v_27886 = mux_27886(v_27887);
  assign v_27887 = ~act_4734;
  assign v_27888 = v_27889 | v_27897;
  assign v_27889 = mux_27889(v_4735);
  assign v_27891 = v_27892 | v_27894;
  assign v_27892 = mux_27892(v_27893);
  assign v_27893 = ~act_4778;
  assign v_27894 = v_27895 | v_27896;
  assign v_27895 = mux_27895(v_4779);
  assign v_27896 = mux_27896(v_4785);
  assign v_27897 = mux_27897(v_4765);
  assign v_27899 = v_27900 | v_27902;
  assign v_27900 = mux_27900(v_27901);
  assign v_27901 = ~act_4741;
  assign v_27902 = v_27903 | v_27904;
  assign v_27903 = mux_27903(v_4742);
  assign v_27904 = mux_27904(v_4748);
  assign v_27905 = mux_27905(v_4721);
  assign v_27907 = v_27908 | v_27910;
  assign v_27908 = mux_27908(v_27909);
  assign v_27909 = ~act_4641;
  assign v_27910 = v_27911 | v_27919;
  assign v_27911 = mux_27911(v_4642);
  assign v_27913 = v_27914 | v_27916;
  assign v_27914 = mux_27914(v_27915);
  assign v_27915 = ~act_4685;
  assign v_27916 = v_27917 | v_27918;
  assign v_27917 = mux_27917(v_4686);
  assign v_27918 = mux_27918(v_4692);
  assign v_27919 = mux_27919(v_4672);
  assign v_27921 = v_27922 | v_27924;
  assign v_27922 = mux_27922(v_27923);
  assign v_27923 = ~act_4648;
  assign v_27924 = v_27925 | v_27926;
  assign v_27925 = mux_27925(v_4649);
  assign v_27926 = mux_27926(v_4655);
  assign v_27927 = mux_27927(v_4621);
  assign v_27929 = v_27930 | v_27932;
  assign v_27930 = mux_27930(v_27931);
  assign v_27931 = ~act_4429;
  assign v_27932 = v_27933 | v_27955;
  assign v_27933 = mux_27933(v_4430);
  assign v_27935 = v_27936 | v_27938;
  assign v_27936 = mux_27936(v_27937);
  assign v_27937 = ~act_4529;
  assign v_27938 = v_27939 | v_27947;
  assign v_27939 = mux_27939(v_4530);
  assign v_27941 = v_27942 | v_27944;
  assign v_27942 = mux_27942(v_27943);
  assign v_27943 = ~act_4573;
  assign v_27944 = v_27945 | v_27946;
  assign v_27945 = mux_27945(v_4574);
  assign v_27946 = mux_27946(v_4580);
  assign v_27947 = mux_27947(v_4560);
  assign v_27949 = v_27950 | v_27952;
  assign v_27950 = mux_27950(v_27951);
  assign v_27951 = ~act_4536;
  assign v_27952 = v_27953 | v_27954;
  assign v_27953 = mux_27953(v_4537);
  assign v_27954 = mux_27954(v_4543);
  assign v_27955 = mux_27955(v_4516);
  assign v_27957 = v_27958 | v_27960;
  assign v_27958 = mux_27958(v_27959);
  assign v_27959 = ~act_4436;
  assign v_27960 = v_27961 | v_27969;
  assign v_27961 = mux_27961(v_4437);
  assign v_27963 = v_27964 | v_27966;
  assign v_27964 = mux_27964(v_27965);
  assign v_27965 = ~act_4480;
  assign v_27966 = v_27967 | v_27968;
  assign v_27967 = mux_27967(v_4481);
  assign v_27968 = mux_27968(v_4487);
  assign v_27969 = mux_27969(v_4467);
  assign v_27971 = v_27972 | v_27974;
  assign v_27972 = mux_27972(v_27973);
  assign v_27973 = ~act_4443;
  assign v_27974 = v_27975 | v_27976;
  assign v_27975 = mux_27975(v_4444);
  assign v_27976 = mux_27976(v_4450);
  assign v_27977 = in0_canPeek;
  assign v_27978 = in0_peek;
  // Always block
  //////////////////////////////////////////////////////////////////////////////
  always @(posedge clock) begin
    if (reset) begin
      v_7 <= 1'h0;
      v_29 <= 1'h0;
      v_36 <= 1'h0;
      v_79 <= 1'h0;
      v_86 <= 1'h0;
      v_93 <= 1'h0;
      v_130 <= 1'h0;
      v_185 <= 1'h0;
      v_192 <= 1'h0;
      v_199 <= 1'h0;
      v_206 <= 1'h0;
      v_243 <= 1'h0;
      v_292 <= 1'h0;
      v_299 <= 1'h0;
      v_336 <= 1'h0;
      v_403 <= 1'h0;
      v_410 <= 1'h0;
      v_417 <= 1'h0;
      v_424 <= 1'h0;
      v_431 <= 1'h0;
      v_468 <= 1'h0;
      v_517 <= 1'h0;
      v_524 <= 1'h0;
      v_561 <= 1'h0;
      v_622 <= 1'h0;
      v_629 <= 1'h0;
      v_636 <= 1'h0;
      v_673 <= 1'h0;
      v_722 <= 1'h0;
      v_729 <= 1'h0;
      v_766 <= 1'h0;
      v_845 <= 1'h0;
      v_852 <= 1'h0;
      v_859 <= 1'h0;
      v_866 <= 1'h0;
      v_873 <= 1'h0;
      v_880 <= 1'h0;
      v_917 <= 1'h0;
      v_966 <= 1'h0;
      v_973 <= 1'h0;
      v_1010 <= 1'h0;
      v_1071 <= 1'h0;
      v_1078 <= 1'h0;
      v_1085 <= 1'h0;
      v_1122 <= 1'h0;
      v_1171 <= 1'h0;
      v_1178 <= 1'h0;
      v_1215 <= 1'h0;
      v_1288 <= 1'h0;
      v_1295 <= 1'h0;
      v_1302 <= 1'h0;
      v_1309 <= 1'h0;
      v_1346 <= 1'h0;
      v_1395 <= 1'h0;
      v_1402 <= 1'h0;
      v_1439 <= 1'h0;
      v_1500 <= 1'h0;
      v_1507 <= 1'h0;
      v_1514 <= 1'h0;
      v_1551 <= 1'h0;
      v_1600 <= 1'h0;
      v_1607 <= 1'h0;
      v_1644 <= 1'h0;
      v_1734 <= 1'h0;
      v_1741 <= 1'h0;
      v_1748 <= 1'h0;
      v_1755 <= 1'h0;
      v_1762 <= 1'h0;
      v_1799 <= 1'h0;
      v_1848 <= 1'h0;
      v_1855 <= 1'h0;
      v_1892 <= 1'h0;
      v_1953 <= 1'h0;
      v_1960 <= 1'h0;
      v_1967 <= 1'h0;
      v_2004 <= 1'h0;
      v_2053 <= 1'h0;
      v_2060 <= 1'h0;
      v_2097 <= 1'h0;
      v_2170 <= 1'h0;
      v_2177 <= 1'h0;
      v_2184 <= 1'h0;
      v_2191 <= 1'h0;
      v_2228 <= 1'h0;
      v_2277 <= 1'h0;
      v_2284 <= 1'h0;
      v_2321 <= 1'h0;
      v_2382 <= 1'h0;
      v_2389 <= 1'h0;
      v_2396 <= 1'h0;
      v_2433 <= 1'h0;
      v_2482 <= 1'h0;
      v_2489 <= 1'h0;
      v_2526 <= 1'h0;
      v_2605 <= 1'h0;
      v_2618 <= 1'h0;
      v_2625 <= 1'h0;
      v_2632 <= 1'h0;
      v_2639 <= 1'h0;
      v_2646 <= 1'h0;
      v_2653 <= 1'h0;
      v_2690 <= 1'h0;
      v_2739 <= 1'h0;
      v_2746 <= 1'h0;
      v_2783 <= 1'h0;
      v_2844 <= 1'h0;
      v_2851 <= 1'h0;
      v_2858 <= 1'h0;
      v_2895 <= 1'h0;
      v_2944 <= 1'h0;
      v_2951 <= 1'h0;
      v_2988 <= 1'h0;
      v_3061 <= 1'h0;
      v_3068 <= 1'h0;
      v_3075 <= 1'h0;
      v_3082 <= 1'h0;
      v_3119 <= 1'h0;
      v_3168 <= 1'h0;
      v_3175 <= 1'h0;
      v_3212 <= 1'h0;
      v_3273 <= 1'h0;
      v_3280 <= 1'h0;
      v_3287 <= 1'h0;
      v_3324 <= 1'h0;
      v_3373 <= 1'h0;
      v_3380 <= 1'h0;
      v_3417 <= 1'h0;
      v_3502 <= 1'h0;
      v_3509 <= 1'h0;
      v_3516 <= 1'h0;
      v_3523 <= 1'h0;
      v_3530 <= 1'h0;
      v_3567 <= 1'h0;
      v_3616 <= 1'h0;
      v_3623 <= 1'h0;
      v_3660 <= 1'h0;
      v_3721 <= 1'h0;
      v_3728 <= 1'h0;
      v_3735 <= 1'h0;
      v_3772 <= 1'h0;
      v_3821 <= 1'h0;
      v_3828 <= 1'h0;
      v_3865 <= 1'h0;
      v_3938 <= 1'h0;
      v_3945 <= 1'h0;
      v_3952 <= 1'h0;
      v_3959 <= 1'h0;
      v_3996 <= 1'h0;
      v_4045 <= 1'h0;
      v_4052 <= 1'h0;
      v_4089 <= 1'h0;
      v_4150 <= 1'h0;
      v_4157 <= 1'h0;
      v_4164 <= 1'h0;
      v_4201 <= 1'h0;
      v_4250 <= 1'h0;
      v_4257 <= 1'h0;
      v_4294 <= 1'h0;
      v_4385 <= 1'h0;
      v_4398 <= 1'h0;
      v_4405 <= 1'h0;
      v_4412 <= 1'h0;
      v_4419 <= 1'h0;
      v_4426 <= 1'h0;
      v_4433 <= 1'h0;
      v_4440 <= 1'h0;
      v_4477 <= 1'h0;
      v_4526 <= 1'h0;
      v_4533 <= 1'h0;
      v_4570 <= 1'h0;
      v_4631 <= 1'h0;
      v_4638 <= 1'h0;
      v_4645 <= 1'h0;
      v_4682 <= 1'h0;
      v_4731 <= 1'h0;
      v_4738 <= 1'h0;
      v_4775 <= 1'h0;
      v_4848 <= 1'h0;
      v_4855 <= 1'h0;
      v_4862 <= 1'h0;
      v_4869 <= 1'h0;
      v_4906 <= 1'h0;
      v_4955 <= 1'h0;
      v_4962 <= 1'h0;
      v_4999 <= 1'h0;
      v_5060 <= 1'h0;
      v_5067 <= 1'h0;
      v_5074 <= 1'h0;
      v_5111 <= 1'h0;
      v_5160 <= 1'h0;
      v_5167 <= 1'h0;
      v_5204 <= 1'h0;
      v_5289 <= 1'h0;
      v_5296 <= 1'h0;
      v_5303 <= 1'h0;
      v_5310 <= 1'h0;
      v_5317 <= 1'h0;
      v_5354 <= 1'h0;
      v_5403 <= 1'h0;
      v_5410 <= 1'h0;
      v_5447 <= 1'h0;
      v_5508 <= 1'h0;
      v_5515 <= 1'h0;
      v_5522 <= 1'h0;
      v_5559 <= 1'h0;
      v_5608 <= 1'h0;
      v_5615 <= 1'h0;
      v_5652 <= 1'h0;
      v_5725 <= 1'h0;
      v_5732 <= 1'h0;
      v_5739 <= 1'h0;
      v_5746 <= 1'h0;
      v_5783 <= 1'h0;
      v_5832 <= 1'h0;
      v_5839 <= 1'h0;
      v_5876 <= 1'h0;
      v_5937 <= 1'h0;
      v_5944 <= 1'h0;
      v_5951 <= 1'h0;
      v_5988 <= 1'h0;
      v_6037 <= 1'h0;
      v_6044 <= 1'h0;
      v_6081 <= 1'h0;
      v_6178 <= 1'h0;
      v_6185 <= 1'h0;
      v_6192 <= 1'h0;
      v_6199 <= 1'h0;
      v_6206 <= 1'h0;
      v_6213 <= 1'h0;
      v_6250 <= 1'h0;
      v_6299 <= 1'h0;
      v_6306 <= 1'h0;
      v_6343 <= 1'h0;
      v_6404 <= 1'h0;
      v_6411 <= 1'h0;
      v_6418 <= 1'h0;
      v_6455 <= 1'h0;
      v_6504 <= 1'h0;
      v_6511 <= 1'h0;
      v_6548 <= 1'h0;
      v_6621 <= 1'h0;
      v_6628 <= 1'h0;
      v_6635 <= 1'h0;
      v_6642 <= 1'h0;
      v_6679 <= 1'h0;
      v_6728 <= 1'h0;
      v_6735 <= 1'h0;
      v_6772 <= 1'h0;
      v_6833 <= 1'h0;
      v_6840 <= 1'h0;
      v_6847 <= 1'h0;
      v_6884 <= 1'h0;
      v_6933 <= 1'h0;
      v_6940 <= 1'h0;
      v_6977 <= 1'h0;
      v_7062 <= 1'h0;
      v_7069 <= 1'h0;
      v_7076 <= 1'h0;
      v_7083 <= 1'h0;
      v_7090 <= 1'h0;
      v_7127 <= 1'h0;
      v_7176 <= 1'h0;
      v_7183 <= 1'h0;
      v_7220 <= 1'h0;
      v_7281 <= 1'h0;
      v_7288 <= 1'h0;
      v_7295 <= 1'h0;
      v_7332 <= 1'h0;
      v_7381 <= 1'h0;
      v_7388 <= 1'h0;
      v_7425 <= 1'h0;
      v_7498 <= 1'h0;
      v_7505 <= 1'h0;
      v_7512 <= 1'h0;
      v_7519 <= 1'h0;
      v_7556 <= 1'h0;
      v_7605 <= 1'h0;
      v_7612 <= 1'h0;
      v_7649 <= 1'h0;
      v_7710 <= 1'h0;
      v_7717 <= 1'h0;
      v_7724 <= 1'h0;
      v_7761 <= 1'h0;
      v_7810 <= 1'h0;
      v_7817 <= 1'h0;
      v_7854 <= 1'h0;
      v_7957 <= 1'h0;
      v_7971 <= 1'h0;
      v_7978 <= 1'h0;
      v_7985 <= 1'h0;
      v_7992 <= 1'h0;
      v_7999 <= 1'h0;
      v_8006 <= 1'h0;
      v_8013 <= 1'h0;
      v_8020 <= 1'h0;
      v_8027 <= 1'h0;
      v_8034 <= 1'h0;
      v_8071 <= 1'h0;
      v_8120 <= 1'h0;
      v_8127 <= 1'h0;
      v_8164 <= 1'h0;
      v_8225 <= 1'h0;
      v_8232 <= 1'h0;
      v_8239 <= 1'h0;
      v_8276 <= 1'h0;
      v_8325 <= 1'h0;
      v_8332 <= 1'h0;
      v_8369 <= 1'h0;
      v_8442 <= 1'h0;
      v_8449 <= 1'h0;
      v_8456 <= 1'h0;
      v_8463 <= 1'h0;
      v_8500 <= 1'h0;
      v_8549 <= 1'h0;
      v_8556 <= 1'h0;
      v_8593 <= 1'h0;
      v_8654 <= 1'h0;
      v_8661 <= 1'h0;
      v_8668 <= 1'h0;
      v_8705 <= 1'h0;
      v_8754 <= 1'h0;
      v_8761 <= 1'h0;
      v_8798 <= 1'h0;
      v_8883 <= 1'h0;
      v_8890 <= 1'h0;
      v_8897 <= 1'h0;
      v_8904 <= 1'h0;
      v_8911 <= 1'h0;
      v_8948 <= 1'h0;
      v_8997 <= 1'h0;
      v_9004 <= 1'h0;
      v_9041 <= 1'h0;
      v_9102 <= 1'h0;
      v_9109 <= 1'h0;
      v_9116 <= 1'h0;
      v_9153 <= 1'h0;
      v_9202 <= 1'h0;
      v_9209 <= 1'h0;
      v_9246 <= 1'h0;
      v_9319 <= 1'h0;
      v_9326 <= 1'h0;
      v_9333 <= 1'h0;
      v_9340 <= 1'h0;
      v_9377 <= 1'h0;
      v_9426 <= 1'h0;
      v_9433 <= 1'h0;
      v_9470 <= 1'h0;
      v_9531 <= 1'h0;
      v_9538 <= 1'h0;
      v_9545 <= 1'h0;
      v_9582 <= 1'h0;
      v_9631 <= 1'h0;
      v_9638 <= 1'h0;
      v_9675 <= 1'h0;
      v_9772 <= 1'h0;
      v_9779 <= 1'h0;
      v_9786 <= 1'h0;
      v_9793 <= 1'h0;
      v_9800 <= 1'h0;
      v_9807 <= 1'h0;
      v_9844 <= 1'h0;
      v_9893 <= 1'h0;
      v_9900 <= 1'h0;
      v_9937 <= 1'h0;
      v_9998 <= 1'h0;
      v_10005 <= 1'h0;
      v_10012 <= 1'h0;
      v_10049 <= 1'h0;
      v_10098 <= 1'h0;
      v_10105 <= 1'h0;
      v_10142 <= 1'h0;
      v_10215 <= 1'h0;
      v_10222 <= 1'h0;
      v_10229 <= 1'h0;
      v_10236 <= 1'h0;
      v_10273 <= 1'h0;
      v_10322 <= 1'h0;
      v_10329 <= 1'h0;
      v_10366 <= 1'h0;
      v_10427 <= 1'h0;
      v_10434 <= 1'h0;
      v_10441 <= 1'h0;
      v_10478 <= 1'h0;
      v_10527 <= 1'h0;
      v_10534 <= 1'h0;
      v_10571 <= 1'h0;
      v_10656 <= 1'h0;
      v_10663 <= 1'h0;
      v_10670 <= 1'h0;
      v_10677 <= 1'h0;
      v_10684 <= 1'h0;
      v_10721 <= 1'h0;
      v_10770 <= 1'h0;
      v_10777 <= 1'h0;
      v_10814 <= 1'h0;
      v_10875 <= 1'h0;
      v_10882 <= 1'h0;
      v_10889 <= 1'h0;
      v_10926 <= 1'h0;
      v_10975 <= 1'h0;
      v_10982 <= 1'h0;
      v_11019 <= 1'h0;
      v_11092 <= 1'h0;
      v_11099 <= 1'h0;
      v_11106 <= 1'h0;
      v_11113 <= 1'h0;
      v_11150 <= 1'h0;
      v_11199 <= 1'h0;
      v_11206 <= 1'h0;
      v_11243 <= 1'h0;
      v_11304 <= 1'h0;
      v_11311 <= 1'h0;
      v_11318 <= 1'h0;
      v_11355 <= 1'h0;
      v_11404 <= 1'h0;
      v_11411 <= 1'h0;
      v_11448 <= 1'h0;
      v_11557 <= 1'h0;
      v_11564 <= 1'h0;
      v_11571 <= 1'h0;
      v_11578 <= 1'h0;
      v_11585 <= 1'h0;
      v_11592 <= 1'h0;
      v_11599 <= 1'h0;
      v_11636 <= 1'h0;
      v_11685 <= 1'h0;
      v_11692 <= 1'h0;
      v_11729 <= 1'h0;
      v_11790 <= 1'h0;
      v_11797 <= 1'h0;
      v_11804 <= 1'h0;
      v_11841 <= 1'h0;
      v_11890 <= 1'h0;
      v_11897 <= 1'h0;
      v_11934 <= 1'h0;
      v_12007 <= 1'h0;
      v_12014 <= 1'h0;
      v_12021 <= 1'h0;
      v_12028 <= 1'h0;
      v_12065 <= 1'h0;
      v_12114 <= 1'h0;
      v_12121 <= 1'h0;
      v_12158 <= 1'h0;
      v_12219 <= 1'h0;
      v_12226 <= 1'h0;
      v_12233 <= 1'h0;
      v_12270 <= 1'h0;
      v_12319 <= 1'h0;
      v_12326 <= 1'h0;
      v_12363 <= 1'h0;
      v_12448 <= 1'h0;
      v_12455 <= 1'h0;
      v_12462 <= 1'h0;
      v_12469 <= 1'h0;
      v_12476 <= 1'h0;
      v_12513 <= 1'h0;
      v_12562 <= 1'h0;
      v_12569 <= 1'h0;
      v_12606 <= 1'h0;
      v_12667 <= 1'h0;
      v_12674 <= 1'h0;
      v_12681 <= 1'h0;
      v_12718 <= 1'h0;
      v_12767 <= 1'h0;
      v_12774 <= 1'h0;
      v_12811 <= 1'h0;
      v_12884 <= 1'h0;
      v_12891 <= 1'h0;
      v_12898 <= 1'h0;
      v_12905 <= 1'h0;
      v_12942 <= 1'h0;
      v_12991 <= 1'h0;
      v_12998 <= 1'h0;
      v_13035 <= 1'h0;
      v_13096 <= 1'h0;
      v_13103 <= 1'h0;
      v_13110 <= 1'h0;
      v_13147 <= 1'h0;
      v_13196 <= 1'h0;
      v_13203 <= 1'h0;
      v_13240 <= 1'h0;
      v_13337 <= 1'h0;
      v_13344 <= 1'h0;
      v_13351 <= 1'h0;
      v_13358 <= 1'h0;
      v_13365 <= 1'h0;
      v_13372 <= 1'h0;
      v_13409 <= 1'h0;
      v_13458 <= 1'h0;
      v_13465 <= 1'h0;
      v_13502 <= 1'h0;
      v_13563 <= 1'h0;
      v_13570 <= 1'h0;
      v_13577 <= 1'h0;
      v_13614 <= 1'h0;
      v_13663 <= 1'h0;
      v_13670 <= 1'h0;
      v_13707 <= 1'h0;
      v_13780 <= 1'h0;
      v_13787 <= 1'h0;
      v_13794 <= 1'h0;
      v_13801 <= 1'h0;
      v_13838 <= 1'h0;
      v_13887 <= 1'h0;
      v_13894 <= 1'h0;
      v_13931 <= 1'h0;
      v_13992 <= 1'h0;
      v_13999 <= 1'h0;
      v_14006 <= 1'h0;
      v_14043 <= 1'h0;
      v_14092 <= 1'h0;
      v_14099 <= 1'h0;
      v_14136 <= 1'h0;
      v_14221 <= 1'h0;
      v_14228 <= 1'h0;
      v_14235 <= 1'h0;
      v_14242 <= 1'h0;
      v_14249 <= 1'h0;
      v_14286 <= 1'h0;
      v_14335 <= 1'h0;
      v_14342 <= 1'h0;
      v_14379 <= 1'h0;
      v_14440 <= 1'h0;
      v_14447 <= 1'h0;
      v_14454 <= 1'h0;
      v_14491 <= 1'h0;
      v_14540 <= 1'h0;
      v_14547 <= 1'h0;
      v_14584 <= 1'h0;
      v_14657 <= 1'h0;
      v_14664 <= 1'h0;
      v_14671 <= 1'h0;
      v_14678 <= 1'h0;
      v_14715 <= 1'h0;
      v_14764 <= 1'h0;
      v_14771 <= 1'h0;
      v_14808 <= 1'h0;
      v_14869 <= 1'h0;
      v_14876 <= 1'h0;
      v_14883 <= 1'h0;
      v_14920 <= 1'h0;
      v_14969 <= 1'h0;
      v_14976 <= 1'h0;
      v_15013 <= 1'h0;
      v_15134 <= 1'h0;
      v_15141 <= 1'h0;
      v_15148 <= 1'h0;
      v_15155 <= 1'h0;
      v_15162 <= 1'h0;
      v_15169 <= 1'h0;
      v_15176 <= 1'h0;
      v_15183 <= 1'h0;
      v_15220 <= 1'h0;
      v_15269 <= 1'h0;
      v_15276 <= 1'h0;
      v_15313 <= 1'h0;
      v_15374 <= 1'h0;
      v_15381 <= 1'h0;
      v_15388 <= 1'h0;
      v_15425 <= 1'h0;
      v_15474 <= 1'h0;
      v_15481 <= 1'h0;
      v_15518 <= 1'h0;
      v_15591 <= 1'h0;
      v_15598 <= 1'h0;
      v_15605 <= 1'h0;
      v_15612 <= 1'h0;
      v_15649 <= 1'h0;
      v_15698 <= 1'h0;
      v_15705 <= 1'h0;
      v_15742 <= 1'h0;
      v_15803 <= 1'h0;
      v_15810 <= 1'h0;
      v_15817 <= 1'h0;
      v_15854 <= 1'h0;
      v_15903 <= 1'h0;
      v_15910 <= 1'h0;
      v_15947 <= 1'h0;
      v_16032 <= 1'h0;
      v_16039 <= 1'h0;
      v_16046 <= 1'h0;
      v_16053 <= 1'h0;
      v_16060 <= 1'h0;
      v_16097 <= 1'h0;
      v_16146 <= 1'h0;
      v_16153 <= 1'h0;
      v_16190 <= 1'h0;
      v_16251 <= 1'h0;
      v_16258 <= 1'h0;
      v_16265 <= 1'h0;
      v_16302 <= 1'h0;
      v_16351 <= 1'h0;
      v_16358 <= 1'h0;
      v_16395 <= 1'h0;
      v_16468 <= 1'h0;
      v_16475 <= 1'h0;
      v_16482 <= 1'h0;
      v_16489 <= 1'h0;
      v_16526 <= 1'h0;
      v_16575 <= 1'h0;
      v_16582 <= 1'h0;
      v_16619 <= 1'h0;
      v_16680 <= 1'h0;
      v_16687 <= 1'h0;
      v_16694 <= 1'h0;
      v_16731 <= 1'h0;
      v_16780 <= 1'h0;
      v_16787 <= 1'h0;
      v_16824 <= 1'h0;
      v_16921 <= 1'h0;
      v_16928 <= 1'h0;
      v_16935 <= 1'h0;
      v_16942 <= 1'h0;
      v_16949 <= 1'h0;
      v_16956 <= 1'h0;
      v_16993 <= 1'h0;
      v_17042 <= 1'h0;
      v_17049 <= 1'h0;
      v_17086 <= 1'h0;
      v_17147 <= 1'h0;
      v_17154 <= 1'h0;
      v_17161 <= 1'h0;
      v_17198 <= 1'h0;
      v_17247 <= 1'h0;
      v_17254 <= 1'h0;
      v_17291 <= 1'h0;
      v_17364 <= 1'h0;
      v_17371 <= 1'h0;
      v_17378 <= 1'h0;
      v_17385 <= 1'h0;
      v_17422 <= 1'h0;
      v_17471 <= 1'h0;
      v_17478 <= 1'h0;
      v_17515 <= 1'h0;
      v_17576 <= 1'h0;
      v_17583 <= 1'h0;
      v_17590 <= 1'h0;
      v_17627 <= 1'h0;
      v_17676 <= 1'h0;
      v_17683 <= 1'h0;
      v_17720 <= 1'h0;
      v_17805 <= 1'h0;
      v_17812 <= 1'h0;
      v_17819 <= 1'h0;
      v_17826 <= 1'h0;
      v_17833 <= 1'h0;
      v_17870 <= 1'h0;
      v_17919 <= 1'h0;
      v_17926 <= 1'h0;
      v_17963 <= 1'h0;
      v_18024 <= 1'h0;
      v_18031 <= 1'h0;
      v_18038 <= 1'h0;
      v_18075 <= 1'h0;
      v_18124 <= 1'h0;
      v_18131 <= 1'h0;
      v_18168 <= 1'h0;
      v_18241 <= 1'h0;
      v_18248 <= 1'h0;
      v_18255 <= 1'h0;
      v_18262 <= 1'h0;
      v_18299 <= 1'h0;
      v_18348 <= 1'h0;
      v_18355 <= 1'h0;
      v_18392 <= 1'h0;
      v_18453 <= 1'h0;
      v_18460 <= 1'h0;
      v_18467 <= 1'h0;
      v_18504 <= 1'h0;
      v_18553 <= 1'h0;
      v_18560 <= 1'h0;
      v_18597 <= 1'h0;
      v_18706 <= 1'h0;
      v_18713 <= 1'h0;
      v_18720 <= 1'h0;
      v_18727 <= 1'h0;
      v_18734 <= 1'h0;
      v_18741 <= 1'h0;
      v_18748 <= 1'h0;
      v_18785 <= 1'h0;
      v_18834 <= 1'h0;
      v_18841 <= 1'h0;
      v_18878 <= 1'h0;
      v_18939 <= 1'h0;
      v_18946 <= 1'h0;
      v_18953 <= 1'h0;
      v_18990 <= 1'h0;
      v_19039 <= 1'h0;
      v_19046 <= 1'h0;
      v_19083 <= 1'h0;
      v_19156 <= 1'h0;
      v_19163 <= 1'h0;
      v_19170 <= 1'h0;
      v_19177 <= 1'h0;
      v_19214 <= 1'h0;
      v_19263 <= 1'h0;
      v_19270 <= 1'h0;
      v_19307 <= 1'h0;
      v_19368 <= 1'h0;
      v_19375 <= 1'h0;
      v_19382 <= 1'h0;
      v_19419 <= 1'h0;
      v_19468 <= 1'h0;
      v_19475 <= 1'h0;
      v_19512 <= 1'h0;
      v_19597 <= 1'h0;
      v_19604 <= 1'h0;
      v_19611 <= 1'h0;
      v_19618 <= 1'h0;
      v_19625 <= 1'h0;
      v_19662 <= 1'h0;
      v_19711 <= 1'h0;
      v_19718 <= 1'h0;
      v_19755 <= 1'h0;
      v_19816 <= 1'h0;
      v_19823 <= 1'h0;
      v_19830 <= 1'h0;
      v_19867 <= 1'h0;
      v_19916 <= 1'h0;
      v_19923 <= 1'h0;
      v_19960 <= 1'h0;
      v_20033 <= 1'h0;
      v_20040 <= 1'h0;
      v_20047 <= 1'h0;
      v_20054 <= 1'h0;
      v_20091 <= 1'h0;
      v_20140 <= 1'h0;
      v_20147 <= 1'h0;
      v_20184 <= 1'h0;
      v_20245 <= 1'h0;
      v_20252 <= 1'h0;
      v_20259 <= 1'h0;
      v_20296 <= 1'h0;
      v_20345 <= 1'h0;
      v_20352 <= 1'h0;
      v_20389 <= 1'h0;
      v_20486 <= 1'h0;
      v_20493 <= 1'h0;
      v_20500 <= 1'h0;
      v_20507 <= 1'h0;
      v_20514 <= 1'h0;
      v_20521 <= 1'h0;
      v_20558 <= 1'h0;
      v_20607 <= 1'h0;
      v_20614 <= 1'h0;
      v_20651 <= 1'h0;
      v_20712 <= 1'h0;
      v_20719 <= 1'h0;
      v_20726 <= 1'h0;
      v_20763 <= 1'h0;
      v_20812 <= 1'h0;
      v_20819 <= 1'h0;
      v_20856 <= 1'h0;
      v_20929 <= 1'h0;
      v_20936 <= 1'h0;
      v_20943 <= 1'h0;
      v_20950 <= 1'h0;
      v_20987 <= 1'h0;
      v_21036 <= 1'h0;
      v_21043 <= 1'h0;
      v_21080 <= 1'h0;
      v_21141 <= 1'h0;
      v_21148 <= 1'h0;
      v_21155 <= 1'h0;
      v_21192 <= 1'h0;
      v_21241 <= 1'h0;
      v_21248 <= 1'h0;
      v_21285 <= 1'h0;
      v_21370 <= 1'h0;
      v_21377 <= 1'h0;
      v_21384 <= 1'h0;
      v_21391 <= 1'h0;
      v_21398 <= 1'h0;
      v_21435 <= 1'h0;
      v_21484 <= 1'h0;
      v_21491 <= 1'h0;
      v_21528 <= 1'h0;
      v_21589 <= 1'h0;
      v_21596 <= 1'h0;
      v_21603 <= 1'h0;
      v_21640 <= 1'h0;
      v_21689 <= 1'h0;
      v_21696 <= 1'h0;
      v_21733 <= 1'h0;
      v_21806 <= 1'h0;
      v_21813 <= 1'h0;
      v_21820 <= 1'h0;
      v_21827 <= 1'h0;
      v_21864 <= 1'h0;
      v_21913 <= 1'h0;
      v_21920 <= 1'h0;
      v_21957 <= 1'h0;
      v_22018 <= 1'h0;
      v_22025 <= 1'h0;
      v_22032 <= 1'h0;
      v_22069 <= 1'h0;
      v_22118 <= 1'h0;
      v_22125 <= 1'h0;
      v_22162 <= 1'h0;
      v_22384 <= 8'h0;
      v_22390 <= 8'h0;
      v_22396 <= 8'h0;
      v_22402 <= 8'h0;
      v_22408 <= 8'h0;
      v_22414 <= 8'h0;
      v_22420 <= 8'h0;
      v_22426 <= 8'h0;
      v_22432 <= 8'h0;
      v_22438 <= 8'h0;
      v_22446 <= 8'h0;
      v_22454 <= 8'h0;
      v_22460 <= 8'h0;
      v_22468 <= 8'h0;
      v_22476 <= 8'h0;
      v_22482 <= 8'h0;
      v_22488 <= 8'h0;
      v_22496 <= 8'h0;
      v_22504 <= 8'h0;
      v_22510 <= 8'h0;
      v_22518 <= 8'h0;
      v_22526 <= 8'h0;
      v_22532 <= 8'h0;
      v_22538 <= 8'h0;
      v_22544 <= 8'h0;
      v_22552 <= 8'h0;
      v_22560 <= 8'h0;
      v_22566 <= 8'h0;
      v_22574 <= 8'h0;
      v_22582 <= 8'h0;
      v_22588 <= 8'h0;
      v_22594 <= 8'h0;
      v_22602 <= 8'h0;
      v_22610 <= 8'h0;
      v_22616 <= 8'h0;
      v_22624 <= 8'h0;
      v_22632 <= 8'h0;
      v_22638 <= 8'h0;
      v_22644 <= 8'h0;
      v_22650 <= 8'h0;
      v_22656 <= 8'h0;
      v_22664 <= 8'h0;
      v_22672 <= 8'h0;
      v_22678 <= 8'h0;
      v_22686 <= 8'h0;
      v_22694 <= 8'h0;
      v_22700 <= 8'h0;
      v_22706 <= 8'h0;
      v_22714 <= 8'h0;
      v_22722 <= 8'h0;
      v_22728 <= 8'h0;
      v_22736 <= 8'h0;
      v_22744 <= 8'h0;
      v_22750 <= 8'h0;
      v_22756 <= 8'h0;
      v_22762 <= 8'h0;
      v_22770 <= 8'h0;
      v_22778 <= 8'h0;
      v_22784 <= 8'h0;
      v_22792 <= 8'h0;
      v_22800 <= 8'h0;
      v_22806 <= 8'h0;
      v_22812 <= 8'h0;
      v_22820 <= 8'h0;
      v_22828 <= 8'h0;
      v_22834 <= 8'h0;
      v_22842 <= 8'h0;
      v_22850 <= 8'h0;
      v_22856 <= 8'h0;
      v_22862 <= 8'h0;
      v_22868 <= 8'h0;
      v_22874 <= 8'h0;
      v_22880 <= 8'h0;
      v_22888 <= 8'h0;
      v_22896 <= 8'h0;
      v_22902 <= 8'h0;
      v_22910 <= 8'h0;
      v_22918 <= 8'h0;
      v_22924 <= 8'h0;
      v_22930 <= 8'h0;
      v_22938 <= 8'h0;
      v_22946 <= 8'h0;
      v_22952 <= 8'h0;
      v_22960 <= 8'h0;
      v_22968 <= 8'h0;
      v_22974 <= 8'h0;
      v_22980 <= 8'h0;
      v_22986 <= 8'h0;
      v_22994 <= 8'h0;
      v_23002 <= 8'h0;
      v_23008 <= 8'h0;
      v_23016 <= 8'h0;
      v_23024 <= 8'h0;
      v_23030 <= 8'h0;
      v_23036 <= 8'h0;
      v_23044 <= 8'h0;
      v_23052 <= 8'h0;
      v_23058 <= 8'h0;
      v_23066 <= 8'h0;
      v_23074 <= 8'h0;
      v_23080 <= 8'h0;
      v_23086 <= 8'h0;
      v_23092 <= 8'h0;
      v_23098 <= 8'h0;
      v_23106 <= 8'h0;
      v_23114 <= 8'h0;
      v_23120 <= 8'h0;
      v_23128 <= 8'h0;
      v_23136 <= 8'h0;
      v_23142 <= 8'h0;
      v_23148 <= 8'h0;
      v_23156 <= 8'h0;
      v_23164 <= 8'h0;
      v_23170 <= 8'h0;
      v_23178 <= 8'h0;
      v_23186 <= 8'h0;
      v_23192 <= 8'h0;
      v_23198 <= 8'h0;
      v_23204 <= 8'h0;
      v_23212 <= 8'h0;
      v_23220 <= 8'h0;
      v_23226 <= 8'h0;
      v_23234 <= 8'h0;
      v_23242 <= 8'h0;
      v_23248 <= 8'h0;
      v_23254 <= 8'h0;
      v_23262 <= 8'h0;
      v_23270 <= 8'h0;
      v_23276 <= 8'h0;
      v_23284 <= 8'h0;
      v_23292 <= 8'h0;
      v_23298 <= 8'h0;
      v_23304 <= 8'h0;
      v_23310 <= 8'h0;
      v_23316 <= 8'h0;
      v_23322 <= 8'h0;
      v_23328 <= 8'h0;
      v_23336 <= 8'h0;
      v_23344 <= 8'h0;
      v_23350 <= 8'h0;
      v_23358 <= 8'h0;
      v_23366 <= 8'h0;
      v_23372 <= 8'h0;
      v_23378 <= 8'h0;
      v_23386 <= 8'h0;
      v_23394 <= 8'h0;
      v_23400 <= 8'h0;
      v_23408 <= 8'h0;
      v_23416 <= 8'h0;
      v_23422 <= 8'h0;
      v_23428 <= 8'h0;
      v_23434 <= 8'h0;
      v_23442 <= 8'h0;
      v_23450 <= 8'h0;
      v_23456 <= 8'h0;
      v_23464 <= 8'h0;
      v_23472 <= 8'h0;
      v_23478 <= 8'h0;
      v_23484 <= 8'h0;
      v_23492 <= 8'h0;
      v_23500 <= 8'h0;
      v_23506 <= 8'h0;
      v_23514 <= 8'h0;
      v_23522 <= 8'h0;
      v_23528 <= 8'h0;
      v_23534 <= 8'h0;
      v_23540 <= 8'h0;
      v_23546 <= 8'h0;
      v_23554 <= 8'h0;
      v_23562 <= 8'h0;
      v_23568 <= 8'h0;
      v_23576 <= 8'h0;
      v_23584 <= 8'h0;
      v_23590 <= 8'h0;
      v_23596 <= 8'h0;
      v_23604 <= 8'h0;
      v_23612 <= 8'h0;
      v_23618 <= 8'h0;
      v_23626 <= 8'h0;
      v_23634 <= 8'h0;
      v_23640 <= 8'h0;
      v_23646 <= 8'h0;
      v_23652 <= 8'h0;
      v_23660 <= 8'h0;
      v_23668 <= 8'h0;
      v_23674 <= 8'h0;
      v_23682 <= 8'h0;
      v_23690 <= 8'h0;
      v_23696 <= 8'h0;
      v_23702 <= 8'h0;
      v_23710 <= 8'h0;
      v_23718 <= 8'h0;
      v_23724 <= 8'h0;
      v_23732 <= 8'h0;
      v_23740 <= 8'h0;
      v_23746 <= 8'h0;
      v_23752 <= 8'h0;
      v_23758 <= 8'h0;
      v_23764 <= 8'h0;
      v_23770 <= 8'h0;
      v_23778 <= 8'h0;
      v_23786 <= 8'h0;
      v_23792 <= 8'h0;
      v_23800 <= 8'h0;
      v_23808 <= 8'h0;
      v_23814 <= 8'h0;
      v_23820 <= 8'h0;
      v_23828 <= 8'h0;
      v_23836 <= 8'h0;
      v_23842 <= 8'h0;
      v_23850 <= 8'h0;
      v_23858 <= 8'h0;
      v_23864 <= 8'h0;
      v_23870 <= 8'h0;
      v_23876 <= 8'h0;
      v_23884 <= 8'h0;
      v_23892 <= 8'h0;
      v_23898 <= 8'h0;
      v_23906 <= 8'h0;
      v_23914 <= 8'h0;
      v_23920 <= 8'h0;
      v_23926 <= 8'h0;
      v_23934 <= 8'h0;
      v_23942 <= 8'h0;
      v_23948 <= 8'h0;
      v_23956 <= 8'h0;
      v_23964 <= 8'h0;
      v_23970 <= 8'h0;
      v_23976 <= 8'h0;
      v_23982 <= 8'h0;
      v_23988 <= 8'h0;
      v_23996 <= 8'h0;
      v_24004 <= 8'h0;
      v_24010 <= 8'h0;
      v_24018 <= 8'h0;
      v_24026 <= 8'h0;
      v_24032 <= 8'h0;
      v_24038 <= 8'h0;
      v_24046 <= 8'h0;
      v_24054 <= 8'h0;
      v_24060 <= 8'h0;
      v_24068 <= 8'h0;
      v_24076 <= 8'h0;
      v_24082 <= 8'h0;
      v_24088 <= 8'h0;
      v_24094 <= 8'h0;
      v_24102 <= 8'h0;
      v_24110 <= 8'h0;
      v_24116 <= 8'h0;
      v_24124 <= 8'h0;
      v_24132 <= 8'h0;
      v_24138 <= 8'h0;
      v_24144 <= 8'h0;
      v_24152 <= 8'h0;
      v_24160 <= 8'h0;
      v_24166 <= 8'h0;
      v_24174 <= 8'h0;
      v_24182 <= 8'h0;
      v_24188 <= 8'h0;
      v_24194 <= 8'h0;
      v_24200 <= 8'h0;
      v_24206 <= 8'h0;
      v_24212 <= 8'h0;
      v_24218 <= 8'h0;
      v_24224 <= 8'h0;
      v_24232 <= 8'h0;
      v_24240 <= 8'h0;
      v_24246 <= 8'h0;
      v_24254 <= 8'h0;
      v_24262 <= 8'h0;
      v_24268 <= 8'h0;
      v_24274 <= 8'h0;
      v_24282 <= 8'h0;
      v_24290 <= 8'h0;
      v_24296 <= 8'h0;
      v_24304 <= 8'h0;
      v_24312 <= 8'h0;
      v_24318 <= 8'h0;
      v_24324 <= 8'h0;
      v_24330 <= 8'h0;
      v_24338 <= 8'h0;
      v_24346 <= 8'h0;
      v_24352 <= 8'h0;
      v_24360 <= 8'h0;
      v_24368 <= 8'h0;
      v_24374 <= 8'h0;
      v_24380 <= 8'h0;
      v_24388 <= 8'h0;
      v_24396 <= 8'h0;
      v_24402 <= 8'h0;
      v_24410 <= 8'h0;
      v_24418 <= 8'h0;
      v_24424 <= 8'h0;
      v_24430 <= 8'h0;
      v_24436 <= 8'h0;
      v_24442 <= 8'h0;
      v_24450 <= 8'h0;
      v_24458 <= 8'h0;
      v_24464 <= 8'h0;
      v_24472 <= 8'h0;
      v_24480 <= 8'h0;
      v_24486 <= 8'h0;
      v_24492 <= 8'h0;
      v_24500 <= 8'h0;
      v_24508 <= 8'h0;
      v_24514 <= 8'h0;
      v_24522 <= 8'h0;
      v_24530 <= 8'h0;
      v_24536 <= 8'h0;
      v_24542 <= 8'h0;
      v_24548 <= 8'h0;
      v_24556 <= 8'h0;
      v_24564 <= 8'h0;
      v_24570 <= 8'h0;
      v_24578 <= 8'h0;
      v_24586 <= 8'h0;
      v_24592 <= 8'h0;
      v_24598 <= 8'h0;
      v_24606 <= 8'h0;
      v_24614 <= 8'h0;
      v_24620 <= 8'h0;
      v_24628 <= 8'h0;
      v_24636 <= 8'h0;
      v_24642 <= 8'h0;
      v_24648 <= 8'h0;
      v_24654 <= 8'h0;
      v_24660 <= 8'h0;
      v_24666 <= 8'h0;
      v_24674 <= 8'h0;
      v_24682 <= 8'h0;
      v_24688 <= 8'h0;
      v_24696 <= 8'h0;
      v_24704 <= 8'h0;
      v_24710 <= 8'h0;
      v_24716 <= 8'h0;
      v_24724 <= 8'h0;
      v_24732 <= 8'h0;
      v_24738 <= 8'h0;
      v_24746 <= 8'h0;
      v_24754 <= 8'h0;
      v_24760 <= 8'h0;
      v_24766 <= 8'h0;
      v_24772 <= 8'h0;
      v_24780 <= 8'h0;
      v_24788 <= 8'h0;
      v_24794 <= 8'h0;
      v_24802 <= 8'h0;
      v_24810 <= 8'h0;
      v_24816 <= 8'h0;
      v_24822 <= 8'h0;
      v_24830 <= 8'h0;
      v_24838 <= 8'h0;
      v_24844 <= 8'h0;
      v_24852 <= 8'h0;
      v_24860 <= 8'h0;
      v_24866 <= 8'h0;
      v_24872 <= 8'h0;
      v_24878 <= 8'h0;
      v_24884 <= 8'h0;
      v_24892 <= 8'h0;
      v_24900 <= 8'h0;
      v_24906 <= 8'h0;
      v_24914 <= 8'h0;
      v_24922 <= 8'h0;
      v_24928 <= 8'h0;
      v_24934 <= 8'h0;
      v_24942 <= 8'h0;
      v_24950 <= 8'h0;
      v_24956 <= 8'h0;
      v_24964 <= 8'h0;
      v_24972 <= 8'h0;
      v_24978 <= 8'h0;
      v_24984 <= 8'h0;
      v_24990 <= 8'h0;
      v_24998 <= 8'h0;
      v_25006 <= 8'h0;
      v_25012 <= 8'h0;
      v_25020 <= 8'h0;
      v_25028 <= 8'h0;
      v_25034 <= 8'h0;
      v_25040 <= 8'h0;
      v_25048 <= 8'h0;
      v_25056 <= 8'h0;
      v_25062 <= 8'h0;
      v_25070 <= 8'h0;
      v_25078 <= 8'h0;
      v_25084 <= 8'h0;
      v_25090 <= 8'h0;
      v_25096 <= 8'h0;
      v_25102 <= 8'h0;
      v_25108 <= 8'h0;
      v_25114 <= 8'h0;
      v_25122 <= 8'h0;
      v_25130 <= 8'h0;
      v_25136 <= 8'h0;
      v_25144 <= 8'h0;
      v_25152 <= 8'h0;
      v_25158 <= 8'h0;
      v_25164 <= 8'h0;
      v_25172 <= 8'h0;
      v_25180 <= 8'h0;
      v_25186 <= 8'h0;
      v_25194 <= 8'h0;
      v_25202 <= 8'h0;
      v_25208 <= 8'h0;
      v_25214 <= 8'h0;
      v_25220 <= 8'h0;
      v_25228 <= 8'h0;
      v_25236 <= 8'h0;
      v_25242 <= 8'h0;
      v_25250 <= 8'h0;
      v_25258 <= 8'h0;
      v_25264 <= 8'h0;
      v_25270 <= 8'h0;
      v_25278 <= 8'h0;
      v_25286 <= 8'h0;
      v_25292 <= 8'h0;
      v_25300 <= 8'h0;
      v_25308 <= 8'h0;
      v_25314 <= 8'h0;
      v_25320 <= 8'h0;
      v_25326 <= 8'h0;
      v_25332 <= 8'h0;
      v_25340 <= 8'h0;
      v_25348 <= 8'h0;
      v_25354 <= 8'h0;
      v_25362 <= 8'h0;
      v_25370 <= 8'h0;
      v_25376 <= 8'h0;
      v_25382 <= 8'h0;
      v_25390 <= 8'h0;
      v_25398 <= 8'h0;
      v_25404 <= 8'h0;
      v_25412 <= 8'h0;
      v_25420 <= 8'h0;
      v_25426 <= 8'h0;
      v_25432 <= 8'h0;
      v_25438 <= 8'h0;
      v_25446 <= 8'h0;
      v_25454 <= 8'h0;
      v_25460 <= 8'h0;
      v_25468 <= 8'h0;
      v_25476 <= 8'h0;
      v_25482 <= 8'h0;
      v_25488 <= 8'h0;
      v_25496 <= 8'h0;
      v_25504 <= 8'h0;
      v_25510 <= 8'h0;
      v_25518 <= 8'h0;
      v_25526 <= 8'h0;
      v_25532 <= 8'h0;
      v_25538 <= 8'h0;
      v_25544 <= 8'h0;
      v_25550 <= 8'h0;
      v_25556 <= 8'h0;
      v_25564 <= 8'h0;
      v_25572 <= 8'h0;
      v_25578 <= 8'h0;
      v_25586 <= 8'h0;
      v_25594 <= 8'h0;
      v_25600 <= 8'h0;
      v_25606 <= 8'h0;
      v_25614 <= 8'h0;
      v_25622 <= 8'h0;
      v_25628 <= 8'h0;
      v_25636 <= 8'h0;
      v_25644 <= 8'h0;
      v_25650 <= 8'h0;
      v_25656 <= 8'h0;
      v_25662 <= 8'h0;
      v_25670 <= 8'h0;
      v_25678 <= 8'h0;
      v_25684 <= 8'h0;
      v_25692 <= 8'h0;
      v_25700 <= 8'h0;
      v_25706 <= 8'h0;
      v_25712 <= 8'h0;
      v_25720 <= 8'h0;
      v_25728 <= 8'h0;
      v_25734 <= 8'h0;
      v_25742 <= 8'h0;
      v_25750 <= 8'h0;
      v_25756 <= 8'h0;
      v_25762 <= 8'h0;
      v_25768 <= 8'h0;
      v_25774 <= 8'h0;
      v_25782 <= 8'h0;
      v_25790 <= 8'h0;
      v_25796 <= 8'h0;
      v_25804 <= 8'h0;
      v_25812 <= 8'h0;
      v_25818 <= 8'h0;
      v_25824 <= 8'h0;
      v_25832 <= 8'h0;
      v_25840 <= 8'h0;
      v_25846 <= 8'h0;
      v_25854 <= 8'h0;
      v_25862 <= 8'h0;
      v_25868 <= 8'h0;
      v_25874 <= 8'h0;
      v_25880 <= 8'h0;
      v_25888 <= 8'h0;
      v_25896 <= 8'h0;
      v_25902 <= 8'h0;
      v_25910 <= 8'h0;
      v_25918 <= 8'h0;
      v_25924 <= 8'h0;
      v_25930 <= 8'h0;
      v_25938 <= 8'h0;
      v_25946 <= 8'h0;
      v_25952 <= 8'h0;
      v_25960 <= 8'h0;
      v_25968 <= 8'h0;
      v_25974 <= 8'h0;
      v_25980 <= 8'h0;
      v_25986 <= 8'h0;
      v_25992 <= 8'h0;
      v_25998 <= 8'h0;
      v_26004 <= 8'h0;
      v_26010 <= 8'h0;
      v_26016 <= 8'h0;
      v_26024 <= 8'h0;
      v_26032 <= 8'h0;
      v_26038 <= 8'h0;
      v_26046 <= 8'h0;
      v_26054 <= 8'h0;
      v_26060 <= 8'h0;
      v_26066 <= 8'h0;
      v_26074 <= 8'h0;
      v_26082 <= 8'h0;
      v_26088 <= 8'h0;
      v_26096 <= 8'h0;
      v_26104 <= 8'h0;
      v_26110 <= 8'h0;
      v_26116 <= 8'h0;
      v_26122 <= 8'h0;
      v_26130 <= 8'h0;
      v_26138 <= 8'h0;
      v_26144 <= 8'h0;
      v_26152 <= 8'h0;
      v_26160 <= 8'h0;
      v_26166 <= 8'h0;
      v_26172 <= 8'h0;
      v_26180 <= 8'h0;
      v_26188 <= 8'h0;
      v_26194 <= 8'h0;
      v_26202 <= 8'h0;
      v_26210 <= 8'h0;
      v_26216 <= 8'h0;
      v_26222 <= 8'h0;
      v_26228 <= 8'h0;
      v_26234 <= 8'h0;
      v_26242 <= 8'h0;
      v_26250 <= 8'h0;
      v_26256 <= 8'h0;
      v_26264 <= 8'h0;
      v_26272 <= 8'h0;
      v_26278 <= 8'h0;
      v_26284 <= 8'h0;
      v_26292 <= 8'h0;
      v_26300 <= 8'h0;
      v_26306 <= 8'h0;
      v_26314 <= 8'h0;
      v_26322 <= 8'h0;
      v_26328 <= 8'h0;
      v_26334 <= 8'h0;
      v_26340 <= 8'h0;
      v_26348 <= 8'h0;
      v_26356 <= 8'h0;
      v_26362 <= 8'h0;
      v_26370 <= 8'h0;
      v_26378 <= 8'h0;
      v_26384 <= 8'h0;
      v_26390 <= 8'h0;
      v_26398 <= 8'h0;
      v_26406 <= 8'h0;
      v_26412 <= 8'h0;
      v_26420 <= 8'h0;
      v_26428 <= 8'h0;
      v_26434 <= 8'h0;
      v_26440 <= 8'h0;
      v_26446 <= 8'h0;
      v_26452 <= 8'h0;
      v_26460 <= 8'h0;
      v_26468 <= 8'h0;
      v_26474 <= 8'h0;
      v_26482 <= 8'h0;
      v_26490 <= 8'h0;
      v_26496 <= 8'h0;
      v_26502 <= 8'h0;
      v_26510 <= 8'h0;
      v_26518 <= 8'h0;
      v_26524 <= 8'h0;
      v_26532 <= 8'h0;
      v_26540 <= 8'h0;
      v_26546 <= 8'h0;
      v_26552 <= 8'h0;
      v_26558 <= 8'h0;
      v_26566 <= 8'h0;
      v_26574 <= 8'h0;
      v_26580 <= 8'h0;
      v_26588 <= 8'h0;
      v_26596 <= 8'h0;
      v_26602 <= 8'h0;
      v_26608 <= 8'h0;
      v_26616 <= 8'h0;
      v_26624 <= 8'h0;
      v_26630 <= 8'h0;
      v_26638 <= 8'h0;
      v_26646 <= 8'h0;
      v_26652 <= 8'h0;
      v_26658 <= 8'h0;
      v_26664 <= 8'h0;
      v_26670 <= 8'h0;
      v_26676 <= 8'h0;
      v_26684 <= 8'h0;
      v_26692 <= 8'h0;
      v_26698 <= 8'h0;
      v_26706 <= 8'h0;
      v_26714 <= 8'h0;
      v_26720 <= 8'h0;
      v_26726 <= 8'h0;
      v_26734 <= 8'h0;
      v_26742 <= 8'h0;
      v_26748 <= 8'h0;
      v_26756 <= 8'h0;
      v_26764 <= 8'h0;
      v_26770 <= 8'h0;
      v_26776 <= 8'h0;
      v_26782 <= 8'h0;
      v_26790 <= 8'h0;
      v_26798 <= 8'h0;
      v_26804 <= 8'h0;
      v_26812 <= 8'h0;
      v_26820 <= 8'h0;
      v_26826 <= 8'h0;
      v_26832 <= 8'h0;
      v_26840 <= 8'h0;
      v_26848 <= 8'h0;
      v_26854 <= 8'h0;
      v_26862 <= 8'h0;
      v_26870 <= 8'h0;
      v_26876 <= 8'h0;
      v_26882 <= 8'h0;
      v_26888 <= 8'h0;
      v_26894 <= 8'h0;
      v_26902 <= 8'h0;
      v_26910 <= 8'h0;
      v_26916 <= 8'h0;
      v_26924 <= 8'h0;
      v_26932 <= 8'h0;
      v_26938 <= 8'h0;
      v_26944 <= 8'h0;
      v_26952 <= 8'h0;
      v_26960 <= 8'h0;
      v_26966 <= 8'h0;
      v_26974 <= 8'h0;
      v_26982 <= 8'h0;
      v_26988 <= 8'h0;
      v_26994 <= 8'h0;
      v_27000 <= 8'h0;
      v_27008 <= 8'h0;
      v_27016 <= 8'h0;
      v_27022 <= 8'h0;
      v_27030 <= 8'h0;
      v_27038 <= 8'h0;
      v_27044 <= 8'h0;
      v_27050 <= 8'h0;
      v_27058 <= 8'h0;
      v_27066 <= 8'h0;
      v_27072 <= 8'h0;
      v_27080 <= 8'h0;
      v_27088 <= 8'h0;
      v_27094 <= 8'h0;
      v_27100 <= 8'h0;
      v_27106 <= 8'h0;
      v_27112 <= 8'h0;
      v_27118 <= 8'h0;
      v_27124 <= 8'h0;
      v_27132 <= 8'h0;
      v_27140 <= 8'h0;
      v_27146 <= 8'h0;
      v_27154 <= 8'h0;
      v_27162 <= 8'h0;
      v_27168 <= 8'h0;
      v_27174 <= 8'h0;
      v_27182 <= 8'h0;
      v_27190 <= 8'h0;
      v_27196 <= 8'h0;
      v_27204 <= 8'h0;
      v_27212 <= 8'h0;
      v_27218 <= 8'h0;
      v_27224 <= 8'h0;
      v_27230 <= 8'h0;
      v_27238 <= 8'h0;
      v_27246 <= 8'h0;
      v_27252 <= 8'h0;
      v_27260 <= 8'h0;
      v_27268 <= 8'h0;
      v_27274 <= 8'h0;
      v_27280 <= 8'h0;
      v_27288 <= 8'h0;
      v_27296 <= 8'h0;
      v_27302 <= 8'h0;
      v_27310 <= 8'h0;
      v_27318 <= 8'h0;
      v_27324 <= 8'h0;
      v_27330 <= 8'h0;
      v_27336 <= 8'h0;
      v_27342 <= 8'h0;
      v_27350 <= 8'h0;
      v_27358 <= 8'h0;
      v_27364 <= 8'h0;
      v_27372 <= 8'h0;
      v_27380 <= 8'h0;
      v_27386 <= 8'h0;
      v_27392 <= 8'h0;
      v_27400 <= 8'h0;
      v_27408 <= 8'h0;
      v_27414 <= 8'h0;
      v_27422 <= 8'h0;
      v_27430 <= 8'h0;
      v_27436 <= 8'h0;
      v_27442 <= 8'h0;
      v_27448 <= 8'h0;
      v_27456 <= 8'h0;
      v_27464 <= 8'h0;
      v_27470 <= 8'h0;
      v_27478 <= 8'h0;
      v_27486 <= 8'h0;
      v_27492 <= 8'h0;
      v_27498 <= 8'h0;
      v_27506 <= 8'h0;
      v_27514 <= 8'h0;
      v_27520 <= 8'h0;
      v_27528 <= 8'h0;
      v_27536 <= 8'h0;
      v_27542 <= 8'h0;
      v_27548 <= 8'h0;
      v_27554 <= 8'h0;
      v_27560 <= 8'h0;
      v_27566 <= 8'h0;
      v_27574 <= 8'h0;
      v_27582 <= 8'h0;
      v_27588 <= 8'h0;
      v_27596 <= 8'h0;
      v_27604 <= 8'h0;
      v_27610 <= 8'h0;
      v_27616 <= 8'h0;
      v_27624 <= 8'h0;
      v_27632 <= 8'h0;
      v_27638 <= 8'h0;
      v_27646 <= 8'h0;
      v_27654 <= 8'h0;
      v_27660 <= 8'h0;
      v_27666 <= 8'h0;
      v_27672 <= 8'h0;
      v_27680 <= 8'h0;
      v_27688 <= 8'h0;
      v_27694 <= 8'h0;
      v_27702 <= 8'h0;
      v_27710 <= 8'h0;
      v_27716 <= 8'h0;
      v_27722 <= 8'h0;
      v_27730 <= 8'h0;
      v_27738 <= 8'h0;
      v_27744 <= 8'h0;
      v_27752 <= 8'h0;
      v_27760 <= 8'h0;
      v_27766 <= 8'h0;
      v_27772 <= 8'h0;
      v_27778 <= 8'h0;
      v_27784 <= 8'h0;
      v_27792 <= 8'h0;
      v_27800 <= 8'h0;
      v_27806 <= 8'h0;
      v_27814 <= 8'h0;
      v_27822 <= 8'h0;
      v_27828 <= 8'h0;
      v_27834 <= 8'h0;
      v_27842 <= 8'h0;
      v_27850 <= 8'h0;
      v_27856 <= 8'h0;
      v_27864 <= 8'h0;
      v_27872 <= 8'h0;
      v_27878 <= 8'h0;
      v_27884 <= 8'h0;
      v_27890 <= 8'h0;
      v_27898 <= 8'h0;
      v_27906 <= 8'h0;
      v_27912 <= 8'h0;
      v_27920 <= 8'h0;
      v_27928 <= 8'h0;
      v_27934 <= 8'h0;
      v_27940 <= 8'h0;
      v_27948 <= 8'h0;
      v_27956 <= 8'h0;
      v_27962 <= 8'h0;
      v_27970 <= 8'h0;
    end else begin
      if (v_8 == 1) v_7 <= v_22374;
      if (v_30 == 1) v_29 <= v_22368;
      if (v_37 == 1) v_36 <= v_66;
      if (v_80 == 1) v_79 <= v_22362;
      if (v_87 == 1) v_86 <= v_172;
      if (v_94 == 1) v_93 <= v_127;
      if (v_131 == 1) v_130 <= v_160;
      if (v_186 == 1) v_185 <= v_22356;
      if (v_193 == 1) v_192 <= v_390;
      if (v_200 == 1) v_199 <= v_289;
      if (v_207 == 1) v_206 <= v_240;
      if (v_244 == 1) v_243 <= v_273;
      if (v_293 == 1) v_292 <= v_378;
      if (v_300 == 1) v_299 <= v_333;
      if (v_337 == 1) v_336 <= v_366;
      if (v_404 == 1) v_403 <= v_22350;
      if (v_411 == 1) v_410 <= v_832;
      if (v_418 == 1) v_417 <= v_619;
      if (v_425 == 1) v_424 <= v_514;
      if (v_432 == 1) v_431 <= v_465;
      if (v_469 == 1) v_468 <= v_498;
      if (v_518 == 1) v_517 <= v_603;
      if (v_525 == 1) v_524 <= v_558;
      if (v_562 == 1) v_561 <= v_591;
      if (v_623 == 1) v_622 <= v_820;
      if (v_630 == 1) v_629 <= v_719;
      if (v_637 == 1) v_636 <= v_670;
      if (v_674 == 1) v_673 <= v_703;
      if (v_723 == 1) v_722 <= v_808;
      if (v_730 == 1) v_729 <= v_763;
      if (v_767 == 1) v_766 <= v_796;
      if (v_846 == 1) v_845 <= v_22344;
      if (v_853 == 1) v_852 <= v_1722;
      if (v_860 == 1) v_859 <= v_1285;
      if (v_867 == 1) v_866 <= v_1068;
      if (v_874 == 1) v_873 <= v_963;
      if (v_881 == 1) v_880 <= v_914;
      if (v_918 == 1) v_917 <= v_947;
      if (v_967 == 1) v_966 <= v_1052;
      if (v_974 == 1) v_973 <= v_1007;
      if (v_1011 == 1) v_1010 <= v_1040;
      if (v_1072 == 1) v_1071 <= v_1269;
      if (v_1079 == 1) v_1078 <= v_1168;
      if (v_1086 == 1) v_1085 <= v_1119;
      if (v_1123 == 1) v_1122 <= v_1152;
      if (v_1172 == 1) v_1171 <= v_1257;
      if (v_1179 == 1) v_1178 <= v_1212;
      if (v_1216 == 1) v_1215 <= v_1245;
      if (v_1289 == 1) v_1288 <= v_1710;
      if (v_1296 == 1) v_1295 <= v_1497;
      if (v_1303 == 1) v_1302 <= v_1392;
      if (v_1310 == 1) v_1309 <= v_1343;
      if (v_1347 == 1) v_1346 <= v_1376;
      if (v_1396 == 1) v_1395 <= v_1481;
      if (v_1403 == 1) v_1402 <= v_1436;
      if (v_1440 == 1) v_1439 <= v_1469;
      if (v_1501 == 1) v_1500 <= v_1698;
      if (v_1508 == 1) v_1507 <= v_1597;
      if (v_1515 == 1) v_1514 <= v_1548;
      if (v_1552 == 1) v_1551 <= v_1581;
      if (v_1601 == 1) v_1600 <= v_1686;
      if (v_1608 == 1) v_1607 <= v_1641;
      if (v_1645 == 1) v_1644 <= v_1674;
      if (v_1735 == 1) v_1734 <= v_22338;
      if (v_1742 == 1) v_1741 <= v_2167;
      if (v_1749 == 1) v_1748 <= v_1950;
      if (v_1756 == 1) v_1755 <= v_1845;
      if (v_1763 == 1) v_1762 <= v_1796;
      if (v_1800 == 1) v_1799 <= v_1829;
      if (v_1849 == 1) v_1848 <= v_1934;
      if (v_1856 == 1) v_1855 <= v_1889;
      if (v_1893 == 1) v_1892 <= v_1922;
      if (v_1954 == 1) v_1953 <= v_2151;
      if (v_1961 == 1) v_1960 <= v_2050;
      if (v_1968 == 1) v_1967 <= v_2001;
      if (v_2005 == 1) v_2004 <= v_2034;
      if (v_2054 == 1) v_2053 <= v_2139;
      if (v_2061 == 1) v_2060 <= v_2094;
      if (v_2098 == 1) v_2097 <= v_2127;
      if (v_2171 == 1) v_2170 <= v_2592;
      if (v_2178 == 1) v_2177 <= v_2379;
      if (v_2185 == 1) v_2184 <= v_2274;
      if (v_2192 == 1) v_2191 <= v_2225;
      if (v_2229 == 1) v_2228 <= v_2258;
      if (v_2278 == 1) v_2277 <= v_2363;
      if (v_2285 == 1) v_2284 <= v_2318;
      if (v_2322 == 1) v_2321 <= v_2351;
      if (v_2383 == 1) v_2382 <= v_2580;
      if (v_2390 == 1) v_2389 <= v_2479;
      if (v_2397 == 1) v_2396 <= v_2430;
      if (v_2434 == 1) v_2433 <= v_2463;
      if (v_2483 == 1) v_2482 <= v_2568;
      if (v_2490 == 1) v_2489 <= v_2523;
      if (v_2527 == 1) v_2526 <= v_2556;
      if (v_2606 == 1) v_2605 <= v_22332;
      if (v_2619 == 1) v_2618 <= v_22326;
      if (v_2626 == 1) v_2625 <= v_3499;
      if (v_2633 == 1) v_2632 <= v_3058;
      if (v_2640 == 1) v_2639 <= v_2841;
      if (v_2647 == 1) v_2646 <= v_2736;
      if (v_2654 == 1) v_2653 <= v_2687;
      if (v_2691 == 1) v_2690 <= v_2720;
      if (v_2740 == 1) v_2739 <= v_2825;
      if (v_2747 == 1) v_2746 <= v_2780;
      if (v_2784 == 1) v_2783 <= v_2813;
      if (v_2845 == 1) v_2844 <= v_3042;
      if (v_2852 == 1) v_2851 <= v_2941;
      if (v_2859 == 1) v_2858 <= v_2892;
      if (v_2896 == 1) v_2895 <= v_2925;
      if (v_2945 == 1) v_2944 <= v_3030;
      if (v_2952 == 1) v_2951 <= v_2985;
      if (v_2989 == 1) v_2988 <= v_3018;
      if (v_3062 == 1) v_3061 <= v_3483;
      if (v_3069 == 1) v_3068 <= v_3270;
      if (v_3076 == 1) v_3075 <= v_3165;
      if (v_3083 == 1) v_3082 <= v_3116;
      if (v_3120 == 1) v_3119 <= v_3149;
      if (v_3169 == 1) v_3168 <= v_3254;
      if (v_3176 == 1) v_3175 <= v_3209;
      if (v_3213 == 1) v_3212 <= v_3242;
      if (v_3274 == 1) v_3273 <= v_3471;
      if (v_3281 == 1) v_3280 <= v_3370;
      if (v_3288 == 1) v_3287 <= v_3321;
      if (v_3325 == 1) v_3324 <= v_3354;
      if (v_3374 == 1) v_3373 <= v_3459;
      if (v_3381 == 1) v_3380 <= v_3414;
      if (v_3418 == 1) v_3417 <= v_3447;
      if (v_3503 == 1) v_3502 <= v_4372;
      if (v_3510 == 1) v_3509 <= v_3935;
      if (v_3517 == 1) v_3516 <= v_3718;
      if (v_3524 == 1) v_3523 <= v_3613;
      if (v_3531 == 1) v_3530 <= v_3564;
      if (v_3568 == 1) v_3567 <= v_3597;
      if (v_3617 == 1) v_3616 <= v_3702;
      if (v_3624 == 1) v_3623 <= v_3657;
      if (v_3661 == 1) v_3660 <= v_3690;
      if (v_3722 == 1) v_3721 <= v_3919;
      if (v_3729 == 1) v_3728 <= v_3818;
      if (v_3736 == 1) v_3735 <= v_3769;
      if (v_3773 == 1) v_3772 <= v_3802;
      if (v_3822 == 1) v_3821 <= v_3907;
      if (v_3829 == 1) v_3828 <= v_3862;
      if (v_3866 == 1) v_3865 <= v_3895;
      if (v_3939 == 1) v_3938 <= v_4360;
      if (v_3946 == 1) v_3945 <= v_4147;
      if (v_3953 == 1) v_3952 <= v_4042;
      if (v_3960 == 1) v_3959 <= v_3993;
      if (v_3997 == 1) v_3996 <= v_4026;
      if (v_4046 == 1) v_4045 <= v_4131;
      if (v_4053 == 1) v_4052 <= v_4086;
      if (v_4090 == 1) v_4089 <= v_4119;
      if (v_4151 == 1) v_4150 <= v_4348;
      if (v_4158 == 1) v_4157 <= v_4247;
      if (v_4165 == 1) v_4164 <= v_4198;
      if (v_4202 == 1) v_4201 <= v_4231;
      if (v_4251 == 1) v_4250 <= v_4336;
      if (v_4258 == 1) v_4257 <= v_4291;
      if (v_4295 == 1) v_4294 <= v_4324;
      if (v_4386 == 1) v_4385 <= v_22320;
      if (v_4399 == 1) v_4398 <= v_22314;
      if (v_4406 == 1) v_4405 <= v_6175;
      if (v_4413 == 1) v_4412 <= v_5286;
      if (v_4420 == 1) v_4419 <= v_4845;
      if (v_4427 == 1) v_4426 <= v_4628;
      if (v_4434 == 1) v_4433 <= v_4523;
      if (v_4441 == 1) v_4440 <= v_4474;
      if (v_4478 == 1) v_4477 <= v_4507;
      if (v_4527 == 1) v_4526 <= v_4612;
      if (v_4534 == 1) v_4533 <= v_4567;
      if (v_4571 == 1) v_4570 <= v_4600;
      if (v_4632 == 1) v_4631 <= v_4829;
      if (v_4639 == 1) v_4638 <= v_4728;
      if (v_4646 == 1) v_4645 <= v_4679;
      if (v_4683 == 1) v_4682 <= v_4712;
      if (v_4732 == 1) v_4731 <= v_4817;
      if (v_4739 == 1) v_4738 <= v_4772;
      if (v_4776 == 1) v_4775 <= v_4805;
      if (v_4849 == 1) v_4848 <= v_5270;
      if (v_4856 == 1) v_4855 <= v_5057;
      if (v_4863 == 1) v_4862 <= v_4952;
      if (v_4870 == 1) v_4869 <= v_4903;
      if (v_4907 == 1) v_4906 <= v_4936;
      if (v_4956 == 1) v_4955 <= v_5041;
      if (v_4963 == 1) v_4962 <= v_4996;
      if (v_5000 == 1) v_4999 <= v_5029;
      if (v_5061 == 1) v_5060 <= v_5258;
      if (v_5068 == 1) v_5067 <= v_5157;
      if (v_5075 == 1) v_5074 <= v_5108;
      if (v_5112 == 1) v_5111 <= v_5141;
      if (v_5161 == 1) v_5160 <= v_5246;
      if (v_5168 == 1) v_5167 <= v_5201;
      if (v_5205 == 1) v_5204 <= v_5234;
      if (v_5290 == 1) v_5289 <= v_6159;
      if (v_5297 == 1) v_5296 <= v_5722;
      if (v_5304 == 1) v_5303 <= v_5505;
      if (v_5311 == 1) v_5310 <= v_5400;
      if (v_5318 == 1) v_5317 <= v_5351;
      if (v_5355 == 1) v_5354 <= v_5384;
      if (v_5404 == 1) v_5403 <= v_5489;
      if (v_5411 == 1) v_5410 <= v_5444;
      if (v_5448 == 1) v_5447 <= v_5477;
      if (v_5509 == 1) v_5508 <= v_5706;
      if (v_5516 == 1) v_5515 <= v_5605;
      if (v_5523 == 1) v_5522 <= v_5556;
      if (v_5560 == 1) v_5559 <= v_5589;
      if (v_5609 == 1) v_5608 <= v_5694;
      if (v_5616 == 1) v_5615 <= v_5649;
      if (v_5653 == 1) v_5652 <= v_5682;
      if (v_5726 == 1) v_5725 <= v_6147;
      if (v_5733 == 1) v_5732 <= v_5934;
      if (v_5740 == 1) v_5739 <= v_5829;
      if (v_5747 == 1) v_5746 <= v_5780;
      if (v_5784 == 1) v_5783 <= v_5813;
      if (v_5833 == 1) v_5832 <= v_5918;
      if (v_5840 == 1) v_5839 <= v_5873;
      if (v_5877 == 1) v_5876 <= v_5906;
      if (v_5938 == 1) v_5937 <= v_6135;
      if (v_5945 == 1) v_5944 <= v_6034;
      if (v_5952 == 1) v_5951 <= v_5985;
      if (v_5989 == 1) v_5988 <= v_6018;
      if (v_6038 == 1) v_6037 <= v_6123;
      if (v_6045 == 1) v_6044 <= v_6078;
      if (v_6082 == 1) v_6081 <= v_6111;
      if (v_6179 == 1) v_6178 <= v_7944;
      if (v_6186 == 1) v_6185 <= v_7059;
      if (v_6193 == 1) v_6192 <= v_6618;
      if (v_6200 == 1) v_6199 <= v_6401;
      if (v_6207 == 1) v_6206 <= v_6296;
      if (v_6214 == 1) v_6213 <= v_6247;
      if (v_6251 == 1) v_6250 <= v_6280;
      if (v_6300 == 1) v_6299 <= v_6385;
      if (v_6307 == 1) v_6306 <= v_6340;
      if (v_6344 == 1) v_6343 <= v_6373;
      if (v_6405 == 1) v_6404 <= v_6602;
      if (v_6412 == 1) v_6411 <= v_6501;
      if (v_6419 == 1) v_6418 <= v_6452;
      if (v_6456 == 1) v_6455 <= v_6485;
      if (v_6505 == 1) v_6504 <= v_6590;
      if (v_6512 == 1) v_6511 <= v_6545;
      if (v_6549 == 1) v_6548 <= v_6578;
      if (v_6622 == 1) v_6621 <= v_7043;
      if (v_6629 == 1) v_6628 <= v_6830;
      if (v_6636 == 1) v_6635 <= v_6725;
      if (v_6643 == 1) v_6642 <= v_6676;
      if (v_6680 == 1) v_6679 <= v_6709;
      if (v_6729 == 1) v_6728 <= v_6814;
      if (v_6736 == 1) v_6735 <= v_6769;
      if (v_6773 == 1) v_6772 <= v_6802;
      if (v_6834 == 1) v_6833 <= v_7031;
      if (v_6841 == 1) v_6840 <= v_6930;
      if (v_6848 == 1) v_6847 <= v_6881;
      if (v_6885 == 1) v_6884 <= v_6914;
      if (v_6934 == 1) v_6933 <= v_7019;
      if (v_6941 == 1) v_6940 <= v_6974;
      if (v_6978 == 1) v_6977 <= v_7007;
      if (v_7063 == 1) v_7062 <= v_7932;
      if (v_7070 == 1) v_7069 <= v_7495;
      if (v_7077 == 1) v_7076 <= v_7278;
      if (v_7084 == 1) v_7083 <= v_7173;
      if (v_7091 == 1) v_7090 <= v_7124;
      if (v_7128 == 1) v_7127 <= v_7157;
      if (v_7177 == 1) v_7176 <= v_7262;
      if (v_7184 == 1) v_7183 <= v_7217;
      if (v_7221 == 1) v_7220 <= v_7250;
      if (v_7282 == 1) v_7281 <= v_7479;
      if (v_7289 == 1) v_7288 <= v_7378;
      if (v_7296 == 1) v_7295 <= v_7329;
      if (v_7333 == 1) v_7332 <= v_7362;
      if (v_7382 == 1) v_7381 <= v_7467;
      if (v_7389 == 1) v_7388 <= v_7422;
      if (v_7426 == 1) v_7425 <= v_7455;
      if (v_7499 == 1) v_7498 <= v_7920;
      if (v_7506 == 1) v_7505 <= v_7707;
      if (v_7513 == 1) v_7512 <= v_7602;
      if (v_7520 == 1) v_7519 <= v_7553;
      if (v_7557 == 1) v_7556 <= v_7586;
      if (v_7606 == 1) v_7605 <= v_7691;
      if (v_7613 == 1) v_7612 <= v_7646;
      if (v_7650 == 1) v_7649 <= v_7679;
      if (v_7711 == 1) v_7710 <= v_7908;
      if (v_7718 == 1) v_7717 <= v_7807;
      if (v_7725 == 1) v_7724 <= v_7758;
      if (v_7762 == 1) v_7761 <= v_7791;
      if (v_7811 == 1) v_7810 <= v_7896;
      if (v_7818 == 1) v_7817 <= v_7851;
      if (v_7855 == 1) v_7854 <= v_7884;
      if (v_7958 == 1) v_7957 <= v_22308;
      if (v_7972 == 1) v_7971 <= v_22302;
      if (v_7979 == 1) v_7978 <= v_22288;
      if (v_7986 == 1) v_7985 <= v_15131;
      if (v_7993 == 1) v_7992 <= v_11554;
      if (v_8000 == 1) v_7999 <= v_9769;
      if (v_8007 == 1) v_8006 <= v_8880;
      if (v_8014 == 1) v_8013 <= v_8439;
      if (v_8021 == 1) v_8020 <= v_8222;
      if (v_8028 == 1) v_8027 <= v_8117;
      if (v_8035 == 1) v_8034 <= v_8068;
      if (v_8072 == 1) v_8071 <= v_8101;
      if (v_8121 == 1) v_8120 <= v_8206;
      if (v_8128 == 1) v_8127 <= v_8161;
      if (v_8165 == 1) v_8164 <= v_8194;
      if (v_8226 == 1) v_8225 <= v_8423;
      if (v_8233 == 1) v_8232 <= v_8322;
      if (v_8240 == 1) v_8239 <= v_8273;
      if (v_8277 == 1) v_8276 <= v_8306;
      if (v_8326 == 1) v_8325 <= v_8411;
      if (v_8333 == 1) v_8332 <= v_8366;
      if (v_8370 == 1) v_8369 <= v_8399;
      if (v_8443 == 1) v_8442 <= v_8864;
      if (v_8450 == 1) v_8449 <= v_8651;
      if (v_8457 == 1) v_8456 <= v_8546;
      if (v_8464 == 1) v_8463 <= v_8497;
      if (v_8501 == 1) v_8500 <= v_8530;
      if (v_8550 == 1) v_8549 <= v_8635;
      if (v_8557 == 1) v_8556 <= v_8590;
      if (v_8594 == 1) v_8593 <= v_8623;
      if (v_8655 == 1) v_8654 <= v_8852;
      if (v_8662 == 1) v_8661 <= v_8751;
      if (v_8669 == 1) v_8668 <= v_8702;
      if (v_8706 == 1) v_8705 <= v_8735;
      if (v_8755 == 1) v_8754 <= v_8840;
      if (v_8762 == 1) v_8761 <= v_8795;
      if (v_8799 == 1) v_8798 <= v_8828;
      if (v_8884 == 1) v_8883 <= v_9753;
      if (v_8891 == 1) v_8890 <= v_9316;
      if (v_8898 == 1) v_8897 <= v_9099;
      if (v_8905 == 1) v_8904 <= v_8994;
      if (v_8912 == 1) v_8911 <= v_8945;
      if (v_8949 == 1) v_8948 <= v_8978;
      if (v_8998 == 1) v_8997 <= v_9083;
      if (v_9005 == 1) v_9004 <= v_9038;
      if (v_9042 == 1) v_9041 <= v_9071;
      if (v_9103 == 1) v_9102 <= v_9300;
      if (v_9110 == 1) v_9109 <= v_9199;
      if (v_9117 == 1) v_9116 <= v_9150;
      if (v_9154 == 1) v_9153 <= v_9183;
      if (v_9203 == 1) v_9202 <= v_9288;
      if (v_9210 == 1) v_9209 <= v_9243;
      if (v_9247 == 1) v_9246 <= v_9276;
      if (v_9320 == 1) v_9319 <= v_9741;
      if (v_9327 == 1) v_9326 <= v_9528;
      if (v_9334 == 1) v_9333 <= v_9423;
      if (v_9341 == 1) v_9340 <= v_9374;
      if (v_9378 == 1) v_9377 <= v_9407;
      if (v_9427 == 1) v_9426 <= v_9512;
      if (v_9434 == 1) v_9433 <= v_9467;
      if (v_9471 == 1) v_9470 <= v_9500;
      if (v_9532 == 1) v_9531 <= v_9729;
      if (v_9539 == 1) v_9538 <= v_9628;
      if (v_9546 == 1) v_9545 <= v_9579;
      if (v_9583 == 1) v_9582 <= v_9612;
      if (v_9632 == 1) v_9631 <= v_9717;
      if (v_9639 == 1) v_9638 <= v_9672;
      if (v_9676 == 1) v_9675 <= v_9705;
      if (v_9773 == 1) v_9772 <= v_11538;
      if (v_9780 == 1) v_9779 <= v_10653;
      if (v_9787 == 1) v_9786 <= v_10212;
      if (v_9794 == 1) v_9793 <= v_9995;
      if (v_9801 == 1) v_9800 <= v_9890;
      if (v_9808 == 1) v_9807 <= v_9841;
      if (v_9845 == 1) v_9844 <= v_9874;
      if (v_9894 == 1) v_9893 <= v_9979;
      if (v_9901 == 1) v_9900 <= v_9934;
      if (v_9938 == 1) v_9937 <= v_9967;
      if (v_9999 == 1) v_9998 <= v_10196;
      if (v_10006 == 1) v_10005 <= v_10095;
      if (v_10013 == 1) v_10012 <= v_10046;
      if (v_10050 == 1) v_10049 <= v_10079;
      if (v_10099 == 1) v_10098 <= v_10184;
      if (v_10106 == 1) v_10105 <= v_10139;
      if (v_10143 == 1) v_10142 <= v_10172;
      if (v_10216 == 1) v_10215 <= v_10637;
      if (v_10223 == 1) v_10222 <= v_10424;
      if (v_10230 == 1) v_10229 <= v_10319;
      if (v_10237 == 1) v_10236 <= v_10270;
      if (v_10274 == 1) v_10273 <= v_10303;
      if (v_10323 == 1) v_10322 <= v_10408;
      if (v_10330 == 1) v_10329 <= v_10363;
      if (v_10367 == 1) v_10366 <= v_10396;
      if (v_10428 == 1) v_10427 <= v_10625;
      if (v_10435 == 1) v_10434 <= v_10524;
      if (v_10442 == 1) v_10441 <= v_10475;
      if (v_10479 == 1) v_10478 <= v_10508;
      if (v_10528 == 1) v_10527 <= v_10613;
      if (v_10535 == 1) v_10534 <= v_10568;
      if (v_10572 == 1) v_10571 <= v_10601;
      if (v_10657 == 1) v_10656 <= v_11526;
      if (v_10664 == 1) v_10663 <= v_11089;
      if (v_10671 == 1) v_10670 <= v_10872;
      if (v_10678 == 1) v_10677 <= v_10767;
      if (v_10685 == 1) v_10684 <= v_10718;
      if (v_10722 == 1) v_10721 <= v_10751;
      if (v_10771 == 1) v_10770 <= v_10856;
      if (v_10778 == 1) v_10777 <= v_10811;
      if (v_10815 == 1) v_10814 <= v_10844;
      if (v_10876 == 1) v_10875 <= v_11073;
      if (v_10883 == 1) v_10882 <= v_10972;
      if (v_10890 == 1) v_10889 <= v_10923;
      if (v_10927 == 1) v_10926 <= v_10956;
      if (v_10976 == 1) v_10975 <= v_11061;
      if (v_10983 == 1) v_10982 <= v_11016;
      if (v_11020 == 1) v_11019 <= v_11049;
      if (v_11093 == 1) v_11092 <= v_11514;
      if (v_11100 == 1) v_11099 <= v_11301;
      if (v_11107 == 1) v_11106 <= v_11196;
      if (v_11114 == 1) v_11113 <= v_11147;
      if (v_11151 == 1) v_11150 <= v_11180;
      if (v_11200 == 1) v_11199 <= v_11285;
      if (v_11207 == 1) v_11206 <= v_11240;
      if (v_11244 == 1) v_11243 <= v_11273;
      if (v_11305 == 1) v_11304 <= v_11502;
      if (v_11312 == 1) v_11311 <= v_11401;
      if (v_11319 == 1) v_11318 <= v_11352;
      if (v_11356 == 1) v_11355 <= v_11385;
      if (v_11405 == 1) v_11404 <= v_11490;
      if (v_11412 == 1) v_11411 <= v_11445;
      if (v_11449 == 1) v_11448 <= v_11478;
      if (v_11558 == 1) v_11557 <= v_15115;
      if (v_11565 == 1) v_11564 <= v_13334;
      if (v_11572 == 1) v_11571 <= v_12445;
      if (v_11579 == 1) v_11578 <= v_12004;
      if (v_11586 == 1) v_11585 <= v_11787;
      if (v_11593 == 1) v_11592 <= v_11682;
      if (v_11600 == 1) v_11599 <= v_11633;
      if (v_11637 == 1) v_11636 <= v_11666;
      if (v_11686 == 1) v_11685 <= v_11771;
      if (v_11693 == 1) v_11692 <= v_11726;
      if (v_11730 == 1) v_11729 <= v_11759;
      if (v_11791 == 1) v_11790 <= v_11988;
      if (v_11798 == 1) v_11797 <= v_11887;
      if (v_11805 == 1) v_11804 <= v_11838;
      if (v_11842 == 1) v_11841 <= v_11871;
      if (v_11891 == 1) v_11890 <= v_11976;
      if (v_11898 == 1) v_11897 <= v_11931;
      if (v_11935 == 1) v_11934 <= v_11964;
      if (v_12008 == 1) v_12007 <= v_12429;
      if (v_12015 == 1) v_12014 <= v_12216;
      if (v_12022 == 1) v_12021 <= v_12111;
      if (v_12029 == 1) v_12028 <= v_12062;
      if (v_12066 == 1) v_12065 <= v_12095;
      if (v_12115 == 1) v_12114 <= v_12200;
      if (v_12122 == 1) v_12121 <= v_12155;
      if (v_12159 == 1) v_12158 <= v_12188;
      if (v_12220 == 1) v_12219 <= v_12417;
      if (v_12227 == 1) v_12226 <= v_12316;
      if (v_12234 == 1) v_12233 <= v_12267;
      if (v_12271 == 1) v_12270 <= v_12300;
      if (v_12320 == 1) v_12319 <= v_12405;
      if (v_12327 == 1) v_12326 <= v_12360;
      if (v_12364 == 1) v_12363 <= v_12393;
      if (v_12449 == 1) v_12448 <= v_13318;
      if (v_12456 == 1) v_12455 <= v_12881;
      if (v_12463 == 1) v_12462 <= v_12664;
      if (v_12470 == 1) v_12469 <= v_12559;
      if (v_12477 == 1) v_12476 <= v_12510;
      if (v_12514 == 1) v_12513 <= v_12543;
      if (v_12563 == 1) v_12562 <= v_12648;
      if (v_12570 == 1) v_12569 <= v_12603;
      if (v_12607 == 1) v_12606 <= v_12636;
      if (v_12668 == 1) v_12667 <= v_12865;
      if (v_12675 == 1) v_12674 <= v_12764;
      if (v_12682 == 1) v_12681 <= v_12715;
      if (v_12719 == 1) v_12718 <= v_12748;
      if (v_12768 == 1) v_12767 <= v_12853;
      if (v_12775 == 1) v_12774 <= v_12808;
      if (v_12812 == 1) v_12811 <= v_12841;
      if (v_12885 == 1) v_12884 <= v_13306;
      if (v_12892 == 1) v_12891 <= v_13093;
      if (v_12899 == 1) v_12898 <= v_12988;
      if (v_12906 == 1) v_12905 <= v_12939;
      if (v_12943 == 1) v_12942 <= v_12972;
      if (v_12992 == 1) v_12991 <= v_13077;
      if (v_12999 == 1) v_12998 <= v_13032;
      if (v_13036 == 1) v_13035 <= v_13065;
      if (v_13097 == 1) v_13096 <= v_13294;
      if (v_13104 == 1) v_13103 <= v_13193;
      if (v_13111 == 1) v_13110 <= v_13144;
      if (v_13148 == 1) v_13147 <= v_13177;
      if (v_13197 == 1) v_13196 <= v_13282;
      if (v_13204 == 1) v_13203 <= v_13237;
      if (v_13241 == 1) v_13240 <= v_13270;
      if (v_13338 == 1) v_13337 <= v_15103;
      if (v_13345 == 1) v_13344 <= v_14218;
      if (v_13352 == 1) v_13351 <= v_13777;
      if (v_13359 == 1) v_13358 <= v_13560;
      if (v_13366 == 1) v_13365 <= v_13455;
      if (v_13373 == 1) v_13372 <= v_13406;
      if (v_13410 == 1) v_13409 <= v_13439;
      if (v_13459 == 1) v_13458 <= v_13544;
      if (v_13466 == 1) v_13465 <= v_13499;
      if (v_13503 == 1) v_13502 <= v_13532;
      if (v_13564 == 1) v_13563 <= v_13761;
      if (v_13571 == 1) v_13570 <= v_13660;
      if (v_13578 == 1) v_13577 <= v_13611;
      if (v_13615 == 1) v_13614 <= v_13644;
      if (v_13664 == 1) v_13663 <= v_13749;
      if (v_13671 == 1) v_13670 <= v_13704;
      if (v_13708 == 1) v_13707 <= v_13737;
      if (v_13781 == 1) v_13780 <= v_14202;
      if (v_13788 == 1) v_13787 <= v_13989;
      if (v_13795 == 1) v_13794 <= v_13884;
      if (v_13802 == 1) v_13801 <= v_13835;
      if (v_13839 == 1) v_13838 <= v_13868;
      if (v_13888 == 1) v_13887 <= v_13973;
      if (v_13895 == 1) v_13894 <= v_13928;
      if (v_13932 == 1) v_13931 <= v_13961;
      if (v_13993 == 1) v_13992 <= v_14190;
      if (v_14000 == 1) v_13999 <= v_14089;
      if (v_14007 == 1) v_14006 <= v_14040;
      if (v_14044 == 1) v_14043 <= v_14073;
      if (v_14093 == 1) v_14092 <= v_14178;
      if (v_14100 == 1) v_14099 <= v_14133;
      if (v_14137 == 1) v_14136 <= v_14166;
      if (v_14222 == 1) v_14221 <= v_15091;
      if (v_14229 == 1) v_14228 <= v_14654;
      if (v_14236 == 1) v_14235 <= v_14437;
      if (v_14243 == 1) v_14242 <= v_14332;
      if (v_14250 == 1) v_14249 <= v_14283;
      if (v_14287 == 1) v_14286 <= v_14316;
      if (v_14336 == 1) v_14335 <= v_14421;
      if (v_14343 == 1) v_14342 <= v_14376;
      if (v_14380 == 1) v_14379 <= v_14409;
      if (v_14441 == 1) v_14440 <= v_14638;
      if (v_14448 == 1) v_14447 <= v_14537;
      if (v_14455 == 1) v_14454 <= v_14488;
      if (v_14492 == 1) v_14491 <= v_14521;
      if (v_14541 == 1) v_14540 <= v_14626;
      if (v_14548 == 1) v_14547 <= v_14581;
      if (v_14585 == 1) v_14584 <= v_14614;
      if (v_14658 == 1) v_14657 <= v_15079;
      if (v_14665 == 1) v_14664 <= v_14866;
      if (v_14672 == 1) v_14671 <= v_14761;
      if (v_14679 == 1) v_14678 <= v_14712;
      if (v_14716 == 1) v_14715 <= v_14745;
      if (v_14765 == 1) v_14764 <= v_14850;
      if (v_14772 == 1) v_14771 <= v_14805;
      if (v_14809 == 1) v_14808 <= v_14838;
      if (v_14870 == 1) v_14869 <= v_15067;
      if (v_14877 == 1) v_14876 <= v_14966;
      if (v_14884 == 1) v_14883 <= v_14917;
      if (v_14921 == 1) v_14920 <= v_14950;
      if (v_14970 == 1) v_14969 <= v_15055;
      if (v_14977 == 1) v_14976 <= v_15010;
      if (v_15014 == 1) v_15013 <= v_15043;
      if (v_15135 == 1) v_15134 <= v_22276;
      if (v_15142 == 1) v_15141 <= v_18703;
      if (v_15149 == 1) v_15148 <= v_16918;
      if (v_15156 == 1) v_15155 <= v_16029;
      if (v_15163 == 1) v_15162 <= v_15588;
      if (v_15170 == 1) v_15169 <= v_15371;
      if (v_15177 == 1) v_15176 <= v_15266;
      if (v_15184 == 1) v_15183 <= v_15217;
      if (v_15221 == 1) v_15220 <= v_15250;
      if (v_15270 == 1) v_15269 <= v_15355;
      if (v_15277 == 1) v_15276 <= v_15310;
      if (v_15314 == 1) v_15313 <= v_15343;
      if (v_15375 == 1) v_15374 <= v_15572;
      if (v_15382 == 1) v_15381 <= v_15471;
      if (v_15389 == 1) v_15388 <= v_15422;
      if (v_15426 == 1) v_15425 <= v_15455;
      if (v_15475 == 1) v_15474 <= v_15560;
      if (v_15482 == 1) v_15481 <= v_15515;
      if (v_15519 == 1) v_15518 <= v_15548;
      if (v_15592 == 1) v_15591 <= v_16013;
      if (v_15599 == 1) v_15598 <= v_15800;
      if (v_15606 == 1) v_15605 <= v_15695;
      if (v_15613 == 1) v_15612 <= v_15646;
      if (v_15650 == 1) v_15649 <= v_15679;
      if (v_15699 == 1) v_15698 <= v_15784;
      if (v_15706 == 1) v_15705 <= v_15739;
      if (v_15743 == 1) v_15742 <= v_15772;
      if (v_15804 == 1) v_15803 <= v_16001;
      if (v_15811 == 1) v_15810 <= v_15900;
      if (v_15818 == 1) v_15817 <= v_15851;
      if (v_15855 == 1) v_15854 <= v_15884;
      if (v_15904 == 1) v_15903 <= v_15989;
      if (v_15911 == 1) v_15910 <= v_15944;
      if (v_15948 == 1) v_15947 <= v_15977;
      if (v_16033 == 1) v_16032 <= v_16902;
      if (v_16040 == 1) v_16039 <= v_16465;
      if (v_16047 == 1) v_16046 <= v_16248;
      if (v_16054 == 1) v_16053 <= v_16143;
      if (v_16061 == 1) v_16060 <= v_16094;
      if (v_16098 == 1) v_16097 <= v_16127;
      if (v_16147 == 1) v_16146 <= v_16232;
      if (v_16154 == 1) v_16153 <= v_16187;
      if (v_16191 == 1) v_16190 <= v_16220;
      if (v_16252 == 1) v_16251 <= v_16449;
      if (v_16259 == 1) v_16258 <= v_16348;
      if (v_16266 == 1) v_16265 <= v_16299;
      if (v_16303 == 1) v_16302 <= v_16332;
      if (v_16352 == 1) v_16351 <= v_16437;
      if (v_16359 == 1) v_16358 <= v_16392;
      if (v_16396 == 1) v_16395 <= v_16425;
      if (v_16469 == 1) v_16468 <= v_16890;
      if (v_16476 == 1) v_16475 <= v_16677;
      if (v_16483 == 1) v_16482 <= v_16572;
      if (v_16490 == 1) v_16489 <= v_16523;
      if (v_16527 == 1) v_16526 <= v_16556;
      if (v_16576 == 1) v_16575 <= v_16661;
      if (v_16583 == 1) v_16582 <= v_16616;
      if (v_16620 == 1) v_16619 <= v_16649;
      if (v_16681 == 1) v_16680 <= v_16878;
      if (v_16688 == 1) v_16687 <= v_16777;
      if (v_16695 == 1) v_16694 <= v_16728;
      if (v_16732 == 1) v_16731 <= v_16761;
      if (v_16781 == 1) v_16780 <= v_16866;
      if (v_16788 == 1) v_16787 <= v_16821;
      if (v_16825 == 1) v_16824 <= v_16854;
      if (v_16922 == 1) v_16921 <= v_18687;
      if (v_16929 == 1) v_16928 <= v_17802;
      if (v_16936 == 1) v_16935 <= v_17361;
      if (v_16943 == 1) v_16942 <= v_17144;
      if (v_16950 == 1) v_16949 <= v_17039;
      if (v_16957 == 1) v_16956 <= v_16990;
      if (v_16994 == 1) v_16993 <= v_17023;
      if (v_17043 == 1) v_17042 <= v_17128;
      if (v_17050 == 1) v_17049 <= v_17083;
      if (v_17087 == 1) v_17086 <= v_17116;
      if (v_17148 == 1) v_17147 <= v_17345;
      if (v_17155 == 1) v_17154 <= v_17244;
      if (v_17162 == 1) v_17161 <= v_17195;
      if (v_17199 == 1) v_17198 <= v_17228;
      if (v_17248 == 1) v_17247 <= v_17333;
      if (v_17255 == 1) v_17254 <= v_17288;
      if (v_17292 == 1) v_17291 <= v_17321;
      if (v_17365 == 1) v_17364 <= v_17786;
      if (v_17372 == 1) v_17371 <= v_17573;
      if (v_17379 == 1) v_17378 <= v_17468;
      if (v_17386 == 1) v_17385 <= v_17419;
      if (v_17423 == 1) v_17422 <= v_17452;
      if (v_17472 == 1) v_17471 <= v_17557;
      if (v_17479 == 1) v_17478 <= v_17512;
      if (v_17516 == 1) v_17515 <= v_17545;
      if (v_17577 == 1) v_17576 <= v_17774;
      if (v_17584 == 1) v_17583 <= v_17673;
      if (v_17591 == 1) v_17590 <= v_17624;
      if (v_17628 == 1) v_17627 <= v_17657;
      if (v_17677 == 1) v_17676 <= v_17762;
      if (v_17684 == 1) v_17683 <= v_17717;
      if (v_17721 == 1) v_17720 <= v_17750;
      if (v_17806 == 1) v_17805 <= v_18675;
      if (v_17813 == 1) v_17812 <= v_18238;
      if (v_17820 == 1) v_17819 <= v_18021;
      if (v_17827 == 1) v_17826 <= v_17916;
      if (v_17834 == 1) v_17833 <= v_17867;
      if (v_17871 == 1) v_17870 <= v_17900;
      if (v_17920 == 1) v_17919 <= v_18005;
      if (v_17927 == 1) v_17926 <= v_17960;
      if (v_17964 == 1) v_17963 <= v_17993;
      if (v_18025 == 1) v_18024 <= v_18222;
      if (v_18032 == 1) v_18031 <= v_18121;
      if (v_18039 == 1) v_18038 <= v_18072;
      if (v_18076 == 1) v_18075 <= v_18105;
      if (v_18125 == 1) v_18124 <= v_18210;
      if (v_18132 == 1) v_18131 <= v_18165;
      if (v_18169 == 1) v_18168 <= v_18198;
      if (v_18242 == 1) v_18241 <= v_18663;
      if (v_18249 == 1) v_18248 <= v_18450;
      if (v_18256 == 1) v_18255 <= v_18345;
      if (v_18263 == 1) v_18262 <= v_18296;
      if (v_18300 == 1) v_18299 <= v_18329;
      if (v_18349 == 1) v_18348 <= v_18434;
      if (v_18356 == 1) v_18355 <= v_18389;
      if (v_18393 == 1) v_18392 <= v_18422;
      if (v_18454 == 1) v_18453 <= v_18651;
      if (v_18461 == 1) v_18460 <= v_18550;
      if (v_18468 == 1) v_18467 <= v_18501;
      if (v_18505 == 1) v_18504 <= v_18534;
      if (v_18554 == 1) v_18553 <= v_18639;
      if (v_18561 == 1) v_18560 <= v_18594;
      if (v_18598 == 1) v_18597 <= v_18627;
      if (v_18707 == 1) v_18706 <= v_22264;
      if (v_18714 == 1) v_18713 <= v_20483;
      if (v_18721 == 1) v_18720 <= v_19594;
      if (v_18728 == 1) v_18727 <= v_19153;
      if (v_18735 == 1) v_18734 <= v_18936;
      if (v_18742 == 1) v_18741 <= v_18831;
      if (v_18749 == 1) v_18748 <= v_18782;
      if (v_18786 == 1) v_18785 <= v_18815;
      if (v_18835 == 1) v_18834 <= v_18920;
      if (v_18842 == 1) v_18841 <= v_18875;
      if (v_18879 == 1) v_18878 <= v_18908;
      if (v_18940 == 1) v_18939 <= v_19137;
      if (v_18947 == 1) v_18946 <= v_19036;
      if (v_18954 == 1) v_18953 <= v_18987;
      if (v_18991 == 1) v_18990 <= v_19020;
      if (v_19040 == 1) v_19039 <= v_19125;
      if (v_19047 == 1) v_19046 <= v_19080;
      if (v_19084 == 1) v_19083 <= v_19113;
      if (v_19157 == 1) v_19156 <= v_19578;
      if (v_19164 == 1) v_19163 <= v_19365;
      if (v_19171 == 1) v_19170 <= v_19260;
      if (v_19178 == 1) v_19177 <= v_19211;
      if (v_19215 == 1) v_19214 <= v_19244;
      if (v_19264 == 1) v_19263 <= v_19349;
      if (v_19271 == 1) v_19270 <= v_19304;
      if (v_19308 == 1) v_19307 <= v_19337;
      if (v_19369 == 1) v_19368 <= v_19566;
      if (v_19376 == 1) v_19375 <= v_19465;
      if (v_19383 == 1) v_19382 <= v_19416;
      if (v_19420 == 1) v_19419 <= v_19449;
      if (v_19469 == 1) v_19468 <= v_19554;
      if (v_19476 == 1) v_19475 <= v_19509;
      if (v_19513 == 1) v_19512 <= v_19542;
      if (v_19598 == 1) v_19597 <= v_20467;
      if (v_19605 == 1) v_19604 <= v_20030;
      if (v_19612 == 1) v_19611 <= v_19813;
      if (v_19619 == 1) v_19618 <= v_19708;
      if (v_19626 == 1) v_19625 <= v_19659;
      if (v_19663 == 1) v_19662 <= v_19692;
      if (v_19712 == 1) v_19711 <= v_19797;
      if (v_19719 == 1) v_19718 <= v_19752;
      if (v_19756 == 1) v_19755 <= v_19785;
      if (v_19817 == 1) v_19816 <= v_20014;
      if (v_19824 == 1) v_19823 <= v_19913;
      if (v_19831 == 1) v_19830 <= v_19864;
      if (v_19868 == 1) v_19867 <= v_19897;
      if (v_19917 == 1) v_19916 <= v_20002;
      if (v_19924 == 1) v_19923 <= v_19957;
      if (v_19961 == 1) v_19960 <= v_19990;
      if (v_20034 == 1) v_20033 <= v_20455;
      if (v_20041 == 1) v_20040 <= v_20242;
      if (v_20048 == 1) v_20047 <= v_20137;
      if (v_20055 == 1) v_20054 <= v_20088;
      if (v_20092 == 1) v_20091 <= v_20121;
      if (v_20141 == 1) v_20140 <= v_20226;
      if (v_20148 == 1) v_20147 <= v_20181;
      if (v_20185 == 1) v_20184 <= v_20214;
      if (v_20246 == 1) v_20245 <= v_20443;
      if (v_20253 == 1) v_20252 <= v_20342;
      if (v_20260 == 1) v_20259 <= v_20293;
      if (v_20297 == 1) v_20296 <= v_20326;
      if (v_20346 == 1) v_20345 <= v_20431;
      if (v_20353 == 1) v_20352 <= v_20386;
      if (v_20390 == 1) v_20389 <= v_20419;
      if (v_20487 == 1) v_20486 <= v_22252;
      if (v_20494 == 1) v_20493 <= v_21367;
      if (v_20501 == 1) v_20500 <= v_20926;
      if (v_20508 == 1) v_20507 <= v_20709;
      if (v_20515 == 1) v_20514 <= v_20604;
      if (v_20522 == 1) v_20521 <= v_20555;
      if (v_20559 == 1) v_20558 <= v_20588;
      if (v_20608 == 1) v_20607 <= v_20693;
      if (v_20615 == 1) v_20614 <= v_20648;
      if (v_20652 == 1) v_20651 <= v_20681;
      if (v_20713 == 1) v_20712 <= v_20910;
      if (v_20720 == 1) v_20719 <= v_20809;
      if (v_20727 == 1) v_20726 <= v_20760;
      if (v_20764 == 1) v_20763 <= v_20793;
      if (v_20813 == 1) v_20812 <= v_20898;
      if (v_20820 == 1) v_20819 <= v_20853;
      if (v_20857 == 1) v_20856 <= v_20886;
      if (v_20930 == 1) v_20929 <= v_21351;
      if (v_20937 == 1) v_20936 <= v_21138;
      if (v_20944 == 1) v_20943 <= v_21033;
      if (v_20951 == 1) v_20950 <= v_20984;
      if (v_20988 == 1) v_20987 <= v_21017;
      if (v_21037 == 1) v_21036 <= v_21122;
      if (v_21044 == 1) v_21043 <= v_21077;
      if (v_21081 == 1) v_21080 <= v_21110;
      if (v_21142 == 1) v_21141 <= v_21339;
      if (v_21149 == 1) v_21148 <= v_21238;
      if (v_21156 == 1) v_21155 <= v_21189;
      if (v_21193 == 1) v_21192 <= v_21222;
      if (v_21242 == 1) v_21241 <= v_21327;
      if (v_21249 == 1) v_21248 <= v_21282;
      if (v_21286 == 1) v_21285 <= v_21315;
      if (v_21371 == 1) v_21370 <= v_22240;
      if (v_21378 == 1) v_21377 <= v_21803;
      if (v_21385 == 1) v_21384 <= v_21586;
      if (v_21392 == 1) v_21391 <= v_21481;
      if (v_21399 == 1) v_21398 <= v_21432;
      if (v_21436 == 1) v_21435 <= v_21465;
      if (v_21485 == 1) v_21484 <= v_21570;
      if (v_21492 == 1) v_21491 <= v_21525;
      if (v_21529 == 1) v_21528 <= v_21558;
      if (v_21590 == 1) v_21589 <= v_21787;
      if (v_21597 == 1) v_21596 <= v_21686;
      if (v_21604 == 1) v_21603 <= v_21637;
      if (v_21641 == 1) v_21640 <= v_21670;
      if (v_21690 == 1) v_21689 <= v_21775;
      if (v_21697 == 1) v_21696 <= v_21730;
      if (v_21734 == 1) v_21733 <= v_21763;
      if (v_21807 == 1) v_21806 <= v_22228;
      if (v_21814 == 1) v_21813 <= v_22015;
      if (v_21821 == 1) v_21820 <= v_21910;
      if (v_21828 == 1) v_21827 <= v_21861;
      if (v_21865 == 1) v_21864 <= v_21894;
      if (v_21914 == 1) v_21913 <= v_21999;
      if (v_21921 == 1) v_21920 <= v_21954;
      if (v_21958 == 1) v_21957 <= v_21987;
      if (v_22019 == 1) v_22018 <= v_22216;
      if (v_22026 == 1) v_22025 <= v_22115;
      if (v_22033 == 1) v_22032 <= v_22066;
      if (v_22070 == 1) v_22069 <= v_22099;
      if (v_22119 == 1) v_22118 <= v_22204;
      if (v_22126 == 1) v_22125 <= v_22159;
      if (v_22163 == 1) v_22162 <= v_22192;
      if (v_7973 == 1) v_22384 <= v_22385;
      if (v_7980 == 1) v_22390 <= v_22391;
      if (v_15136 == 1) v_22396 <= v_22397;
      if (v_18708 == 1) v_22402 <= v_22403;
      if (v_20488 == 1) v_22408 <= v_22409;
      if (v_21372 == 1) v_22414 <= v_22415;
      if (v_21808 == 1) v_22420 <= v_22421;
      if (v_22020 == 1) v_22426 <= v_22427;
      if (v_22120 == 1) v_22432 <= v_22433;
      if (v_22164 == 1) v_22438 <= v_22439;
      if (v_22127 == 1) v_22446 <= v_22447;
      if (v_22027 == 1) v_22454 <= v_22455;
      if (v_22071 == 1) v_22460 <= v_22461;
      if (v_22034 == 1) v_22468 <= v_22469;
      if (v_21815 == 1) v_22476 <= v_22477;
      if (v_21915 == 1) v_22482 <= v_22483;
      if (v_21959 == 1) v_22488 <= v_22489;
      if (v_21922 == 1) v_22496 <= v_22497;
      if (v_21822 == 1) v_22504 <= v_22505;
      if (v_21866 == 1) v_22510 <= v_22511;
      if (v_21829 == 1) v_22518 <= v_22519;
      if (v_21379 == 1) v_22526 <= v_22527;
      if (v_21591 == 1) v_22532 <= v_22533;
      if (v_21691 == 1) v_22538 <= v_22539;
      if (v_21735 == 1) v_22544 <= v_22545;
      if (v_21698 == 1) v_22552 <= v_22553;
      if (v_21598 == 1) v_22560 <= v_22561;
      if (v_21642 == 1) v_22566 <= v_22567;
      if (v_21605 == 1) v_22574 <= v_22575;
      if (v_21386 == 1) v_22582 <= v_22583;
      if (v_21486 == 1) v_22588 <= v_22589;
      if (v_21530 == 1) v_22594 <= v_22595;
      if (v_21493 == 1) v_22602 <= v_22603;
      if (v_21393 == 1) v_22610 <= v_22611;
      if (v_21437 == 1) v_22616 <= v_22617;
      if (v_21400 == 1) v_22624 <= v_22625;
      if (v_20495 == 1) v_22632 <= v_22633;
      if (v_20931 == 1) v_22638 <= v_22639;
      if (v_21143 == 1) v_22644 <= v_22645;
      if (v_21243 == 1) v_22650 <= v_22651;
      if (v_21287 == 1) v_22656 <= v_22657;
      if (v_21250 == 1) v_22664 <= v_22665;
      if (v_21150 == 1) v_22672 <= v_22673;
      if (v_21194 == 1) v_22678 <= v_22679;
      if (v_21157 == 1) v_22686 <= v_22687;
      if (v_20938 == 1) v_22694 <= v_22695;
      if (v_21038 == 1) v_22700 <= v_22701;
      if (v_21082 == 1) v_22706 <= v_22707;
      if (v_21045 == 1) v_22714 <= v_22715;
      if (v_20945 == 1) v_22722 <= v_22723;
      if (v_20989 == 1) v_22728 <= v_22729;
      if (v_20952 == 1) v_22736 <= v_22737;
      if (v_20502 == 1) v_22744 <= v_22745;
      if (v_20714 == 1) v_22750 <= v_22751;
      if (v_20814 == 1) v_22756 <= v_22757;
      if (v_20858 == 1) v_22762 <= v_22763;
      if (v_20821 == 1) v_22770 <= v_22771;
      if (v_20721 == 1) v_22778 <= v_22779;
      if (v_20765 == 1) v_22784 <= v_22785;
      if (v_20728 == 1) v_22792 <= v_22793;
      if (v_20509 == 1) v_22800 <= v_22801;
      if (v_20609 == 1) v_22806 <= v_22807;
      if (v_20653 == 1) v_22812 <= v_22813;
      if (v_20616 == 1) v_22820 <= v_22821;
      if (v_20516 == 1) v_22828 <= v_22829;
      if (v_20560 == 1) v_22834 <= v_22835;
      if (v_20523 == 1) v_22842 <= v_22843;
      if (v_18715 == 1) v_22850 <= v_22851;
      if (v_19599 == 1) v_22856 <= v_22857;
      if (v_20035 == 1) v_22862 <= v_22863;
      if (v_20247 == 1) v_22868 <= v_22869;
      if (v_20347 == 1) v_22874 <= v_22875;
      if (v_20391 == 1) v_22880 <= v_22881;
      if (v_20354 == 1) v_22888 <= v_22889;
      if (v_20254 == 1) v_22896 <= v_22897;
      if (v_20298 == 1) v_22902 <= v_22903;
      if (v_20261 == 1) v_22910 <= v_22911;
      if (v_20042 == 1) v_22918 <= v_22919;
      if (v_20142 == 1) v_22924 <= v_22925;
      if (v_20186 == 1) v_22930 <= v_22931;
      if (v_20149 == 1) v_22938 <= v_22939;
      if (v_20049 == 1) v_22946 <= v_22947;
      if (v_20093 == 1) v_22952 <= v_22953;
      if (v_20056 == 1) v_22960 <= v_22961;
      if (v_19606 == 1) v_22968 <= v_22969;
      if (v_19818 == 1) v_22974 <= v_22975;
      if (v_19918 == 1) v_22980 <= v_22981;
      if (v_19962 == 1) v_22986 <= v_22987;
      if (v_19925 == 1) v_22994 <= v_22995;
      if (v_19825 == 1) v_23002 <= v_23003;
      if (v_19869 == 1) v_23008 <= v_23009;
      if (v_19832 == 1) v_23016 <= v_23017;
      if (v_19613 == 1) v_23024 <= v_23025;
      if (v_19713 == 1) v_23030 <= v_23031;
      if (v_19757 == 1) v_23036 <= v_23037;
      if (v_19720 == 1) v_23044 <= v_23045;
      if (v_19620 == 1) v_23052 <= v_23053;
      if (v_19664 == 1) v_23058 <= v_23059;
      if (v_19627 == 1) v_23066 <= v_23067;
      if (v_18722 == 1) v_23074 <= v_23075;
      if (v_19158 == 1) v_23080 <= v_23081;
      if (v_19370 == 1) v_23086 <= v_23087;
      if (v_19470 == 1) v_23092 <= v_23093;
      if (v_19514 == 1) v_23098 <= v_23099;
      if (v_19477 == 1) v_23106 <= v_23107;
      if (v_19377 == 1) v_23114 <= v_23115;
      if (v_19421 == 1) v_23120 <= v_23121;
      if (v_19384 == 1) v_23128 <= v_23129;
      if (v_19165 == 1) v_23136 <= v_23137;
      if (v_19265 == 1) v_23142 <= v_23143;
      if (v_19309 == 1) v_23148 <= v_23149;
      if (v_19272 == 1) v_23156 <= v_23157;
      if (v_19172 == 1) v_23164 <= v_23165;
      if (v_19216 == 1) v_23170 <= v_23171;
      if (v_19179 == 1) v_23178 <= v_23179;
      if (v_18729 == 1) v_23186 <= v_23187;
      if (v_18941 == 1) v_23192 <= v_23193;
      if (v_19041 == 1) v_23198 <= v_23199;
      if (v_19085 == 1) v_23204 <= v_23205;
      if (v_19048 == 1) v_23212 <= v_23213;
      if (v_18948 == 1) v_23220 <= v_23221;
      if (v_18992 == 1) v_23226 <= v_23227;
      if (v_18955 == 1) v_23234 <= v_23235;
      if (v_18736 == 1) v_23242 <= v_23243;
      if (v_18836 == 1) v_23248 <= v_23249;
      if (v_18880 == 1) v_23254 <= v_23255;
      if (v_18843 == 1) v_23262 <= v_23263;
      if (v_18743 == 1) v_23270 <= v_23271;
      if (v_18787 == 1) v_23276 <= v_23277;
      if (v_18750 == 1) v_23284 <= v_23285;
      if (v_15143 == 1) v_23292 <= v_23293;
      if (v_16923 == 1) v_23298 <= v_23299;
      if (v_17807 == 1) v_23304 <= v_23305;
      if (v_18243 == 1) v_23310 <= v_23311;
      if (v_18455 == 1) v_23316 <= v_23317;
      if (v_18555 == 1) v_23322 <= v_23323;
      if (v_18599 == 1) v_23328 <= v_23329;
      if (v_18562 == 1) v_23336 <= v_23337;
      if (v_18462 == 1) v_23344 <= v_23345;
      if (v_18506 == 1) v_23350 <= v_23351;
      if (v_18469 == 1) v_23358 <= v_23359;
      if (v_18250 == 1) v_23366 <= v_23367;
      if (v_18350 == 1) v_23372 <= v_23373;
      if (v_18394 == 1) v_23378 <= v_23379;
      if (v_18357 == 1) v_23386 <= v_23387;
      if (v_18257 == 1) v_23394 <= v_23395;
      if (v_18301 == 1) v_23400 <= v_23401;
      if (v_18264 == 1) v_23408 <= v_23409;
      if (v_17814 == 1) v_23416 <= v_23417;
      if (v_18026 == 1) v_23422 <= v_23423;
      if (v_18126 == 1) v_23428 <= v_23429;
      if (v_18170 == 1) v_23434 <= v_23435;
      if (v_18133 == 1) v_23442 <= v_23443;
      if (v_18033 == 1) v_23450 <= v_23451;
      if (v_18077 == 1) v_23456 <= v_23457;
      if (v_18040 == 1) v_23464 <= v_23465;
      if (v_17821 == 1) v_23472 <= v_23473;
      if (v_17921 == 1) v_23478 <= v_23479;
      if (v_17965 == 1) v_23484 <= v_23485;
      if (v_17928 == 1) v_23492 <= v_23493;
      if (v_17828 == 1) v_23500 <= v_23501;
      if (v_17872 == 1) v_23506 <= v_23507;
      if (v_17835 == 1) v_23514 <= v_23515;
      if (v_16930 == 1) v_23522 <= v_23523;
      if (v_17366 == 1) v_23528 <= v_23529;
      if (v_17578 == 1) v_23534 <= v_23535;
      if (v_17678 == 1) v_23540 <= v_23541;
      if (v_17722 == 1) v_23546 <= v_23547;
      if (v_17685 == 1) v_23554 <= v_23555;
      if (v_17585 == 1) v_23562 <= v_23563;
      if (v_17629 == 1) v_23568 <= v_23569;
      if (v_17592 == 1) v_23576 <= v_23577;
      if (v_17373 == 1) v_23584 <= v_23585;
      if (v_17473 == 1) v_23590 <= v_23591;
      if (v_17517 == 1) v_23596 <= v_23597;
      if (v_17480 == 1) v_23604 <= v_23605;
      if (v_17380 == 1) v_23612 <= v_23613;
      if (v_17424 == 1) v_23618 <= v_23619;
      if (v_17387 == 1) v_23626 <= v_23627;
      if (v_16937 == 1) v_23634 <= v_23635;
      if (v_17149 == 1) v_23640 <= v_23641;
      if (v_17249 == 1) v_23646 <= v_23647;
      if (v_17293 == 1) v_23652 <= v_23653;
      if (v_17256 == 1) v_23660 <= v_23661;
      if (v_17156 == 1) v_23668 <= v_23669;
      if (v_17200 == 1) v_23674 <= v_23675;
      if (v_17163 == 1) v_23682 <= v_23683;
      if (v_16944 == 1) v_23690 <= v_23691;
      if (v_17044 == 1) v_23696 <= v_23697;
      if (v_17088 == 1) v_23702 <= v_23703;
      if (v_17051 == 1) v_23710 <= v_23711;
      if (v_16951 == 1) v_23718 <= v_23719;
      if (v_16995 == 1) v_23724 <= v_23725;
      if (v_16958 == 1) v_23732 <= v_23733;
      if (v_15150 == 1) v_23740 <= v_23741;
      if (v_16034 == 1) v_23746 <= v_23747;
      if (v_16470 == 1) v_23752 <= v_23753;
      if (v_16682 == 1) v_23758 <= v_23759;
      if (v_16782 == 1) v_23764 <= v_23765;
      if (v_16826 == 1) v_23770 <= v_23771;
      if (v_16789 == 1) v_23778 <= v_23779;
      if (v_16689 == 1) v_23786 <= v_23787;
      if (v_16733 == 1) v_23792 <= v_23793;
      if (v_16696 == 1) v_23800 <= v_23801;
      if (v_16477 == 1) v_23808 <= v_23809;
      if (v_16577 == 1) v_23814 <= v_23815;
      if (v_16621 == 1) v_23820 <= v_23821;
      if (v_16584 == 1) v_23828 <= v_23829;
      if (v_16484 == 1) v_23836 <= v_23837;
      if (v_16528 == 1) v_23842 <= v_23843;
      if (v_16491 == 1) v_23850 <= v_23851;
      if (v_16041 == 1) v_23858 <= v_23859;
      if (v_16253 == 1) v_23864 <= v_23865;
      if (v_16353 == 1) v_23870 <= v_23871;
      if (v_16397 == 1) v_23876 <= v_23877;
      if (v_16360 == 1) v_23884 <= v_23885;
      if (v_16260 == 1) v_23892 <= v_23893;
      if (v_16304 == 1) v_23898 <= v_23899;
      if (v_16267 == 1) v_23906 <= v_23907;
      if (v_16048 == 1) v_23914 <= v_23915;
      if (v_16148 == 1) v_23920 <= v_23921;
      if (v_16192 == 1) v_23926 <= v_23927;
      if (v_16155 == 1) v_23934 <= v_23935;
      if (v_16055 == 1) v_23942 <= v_23943;
      if (v_16099 == 1) v_23948 <= v_23949;
      if (v_16062 == 1) v_23956 <= v_23957;
      if (v_15157 == 1) v_23964 <= v_23965;
      if (v_15593 == 1) v_23970 <= v_23971;
      if (v_15805 == 1) v_23976 <= v_23977;
      if (v_15905 == 1) v_23982 <= v_23983;
      if (v_15949 == 1) v_23988 <= v_23989;
      if (v_15912 == 1) v_23996 <= v_23997;
      if (v_15812 == 1) v_24004 <= v_24005;
      if (v_15856 == 1) v_24010 <= v_24011;
      if (v_15819 == 1) v_24018 <= v_24019;
      if (v_15600 == 1) v_24026 <= v_24027;
      if (v_15700 == 1) v_24032 <= v_24033;
      if (v_15744 == 1) v_24038 <= v_24039;
      if (v_15707 == 1) v_24046 <= v_24047;
      if (v_15607 == 1) v_24054 <= v_24055;
      if (v_15651 == 1) v_24060 <= v_24061;
      if (v_15614 == 1) v_24068 <= v_24069;
      if (v_15164 == 1) v_24076 <= v_24077;
      if (v_15376 == 1) v_24082 <= v_24083;
      if (v_15476 == 1) v_24088 <= v_24089;
      if (v_15520 == 1) v_24094 <= v_24095;
      if (v_15483 == 1) v_24102 <= v_24103;
      if (v_15383 == 1) v_24110 <= v_24111;
      if (v_15427 == 1) v_24116 <= v_24117;
      if (v_15390 == 1) v_24124 <= v_24125;
      if (v_15171 == 1) v_24132 <= v_24133;
      if (v_15271 == 1) v_24138 <= v_24139;
      if (v_15315 == 1) v_24144 <= v_24145;
      if (v_15278 == 1) v_24152 <= v_24153;
      if (v_15178 == 1) v_24160 <= v_24161;
      if (v_15222 == 1) v_24166 <= v_24167;
      if (v_15185 == 1) v_24174 <= v_24175;
      if (v_7987 == 1) v_24182 <= v_24183;
      if (v_11559 == 1) v_24188 <= v_24189;
      if (v_13339 == 1) v_24194 <= v_24195;
      if (v_14223 == 1) v_24200 <= v_24201;
      if (v_14659 == 1) v_24206 <= v_24207;
      if (v_14871 == 1) v_24212 <= v_24213;
      if (v_14971 == 1) v_24218 <= v_24219;
      if (v_15015 == 1) v_24224 <= v_24225;
      if (v_14978 == 1) v_24232 <= v_24233;
      if (v_14878 == 1) v_24240 <= v_24241;
      if (v_14922 == 1) v_24246 <= v_24247;
      if (v_14885 == 1) v_24254 <= v_24255;
      if (v_14666 == 1) v_24262 <= v_24263;
      if (v_14766 == 1) v_24268 <= v_24269;
      if (v_14810 == 1) v_24274 <= v_24275;
      if (v_14773 == 1) v_24282 <= v_24283;
      if (v_14673 == 1) v_24290 <= v_24291;
      if (v_14717 == 1) v_24296 <= v_24297;
      if (v_14680 == 1) v_24304 <= v_24305;
      if (v_14230 == 1) v_24312 <= v_24313;
      if (v_14442 == 1) v_24318 <= v_24319;
      if (v_14542 == 1) v_24324 <= v_24325;
      if (v_14586 == 1) v_24330 <= v_24331;
      if (v_14549 == 1) v_24338 <= v_24339;
      if (v_14449 == 1) v_24346 <= v_24347;
      if (v_14493 == 1) v_24352 <= v_24353;
      if (v_14456 == 1) v_24360 <= v_24361;
      if (v_14237 == 1) v_24368 <= v_24369;
      if (v_14337 == 1) v_24374 <= v_24375;
      if (v_14381 == 1) v_24380 <= v_24381;
      if (v_14344 == 1) v_24388 <= v_24389;
      if (v_14244 == 1) v_24396 <= v_24397;
      if (v_14288 == 1) v_24402 <= v_24403;
      if (v_14251 == 1) v_24410 <= v_24411;
      if (v_13346 == 1) v_24418 <= v_24419;
      if (v_13782 == 1) v_24424 <= v_24425;
      if (v_13994 == 1) v_24430 <= v_24431;
      if (v_14094 == 1) v_24436 <= v_24437;
      if (v_14138 == 1) v_24442 <= v_24443;
      if (v_14101 == 1) v_24450 <= v_24451;
      if (v_14001 == 1) v_24458 <= v_24459;
      if (v_14045 == 1) v_24464 <= v_24465;
      if (v_14008 == 1) v_24472 <= v_24473;
      if (v_13789 == 1) v_24480 <= v_24481;
      if (v_13889 == 1) v_24486 <= v_24487;
      if (v_13933 == 1) v_24492 <= v_24493;
      if (v_13896 == 1) v_24500 <= v_24501;
      if (v_13796 == 1) v_24508 <= v_24509;
      if (v_13840 == 1) v_24514 <= v_24515;
      if (v_13803 == 1) v_24522 <= v_24523;
      if (v_13353 == 1) v_24530 <= v_24531;
      if (v_13565 == 1) v_24536 <= v_24537;
      if (v_13665 == 1) v_24542 <= v_24543;
      if (v_13709 == 1) v_24548 <= v_24549;
      if (v_13672 == 1) v_24556 <= v_24557;
      if (v_13572 == 1) v_24564 <= v_24565;
      if (v_13616 == 1) v_24570 <= v_24571;
      if (v_13579 == 1) v_24578 <= v_24579;
      if (v_13360 == 1) v_24586 <= v_24587;
      if (v_13460 == 1) v_24592 <= v_24593;
      if (v_13504 == 1) v_24598 <= v_24599;
      if (v_13467 == 1) v_24606 <= v_24607;
      if (v_13367 == 1) v_24614 <= v_24615;
      if (v_13411 == 1) v_24620 <= v_24621;
      if (v_13374 == 1) v_24628 <= v_24629;
      if (v_11566 == 1) v_24636 <= v_24637;
      if (v_12450 == 1) v_24642 <= v_24643;
      if (v_12886 == 1) v_24648 <= v_24649;
      if (v_13098 == 1) v_24654 <= v_24655;
      if (v_13198 == 1) v_24660 <= v_24661;
      if (v_13242 == 1) v_24666 <= v_24667;
      if (v_13205 == 1) v_24674 <= v_24675;
      if (v_13105 == 1) v_24682 <= v_24683;
      if (v_13149 == 1) v_24688 <= v_24689;
      if (v_13112 == 1) v_24696 <= v_24697;
      if (v_12893 == 1) v_24704 <= v_24705;
      if (v_12993 == 1) v_24710 <= v_24711;
      if (v_13037 == 1) v_24716 <= v_24717;
      if (v_13000 == 1) v_24724 <= v_24725;
      if (v_12900 == 1) v_24732 <= v_24733;
      if (v_12944 == 1) v_24738 <= v_24739;
      if (v_12907 == 1) v_24746 <= v_24747;
      if (v_12457 == 1) v_24754 <= v_24755;
      if (v_12669 == 1) v_24760 <= v_24761;
      if (v_12769 == 1) v_24766 <= v_24767;
      if (v_12813 == 1) v_24772 <= v_24773;
      if (v_12776 == 1) v_24780 <= v_24781;
      if (v_12676 == 1) v_24788 <= v_24789;
      if (v_12720 == 1) v_24794 <= v_24795;
      if (v_12683 == 1) v_24802 <= v_24803;
      if (v_12464 == 1) v_24810 <= v_24811;
      if (v_12564 == 1) v_24816 <= v_24817;
      if (v_12608 == 1) v_24822 <= v_24823;
      if (v_12571 == 1) v_24830 <= v_24831;
      if (v_12471 == 1) v_24838 <= v_24839;
      if (v_12515 == 1) v_24844 <= v_24845;
      if (v_12478 == 1) v_24852 <= v_24853;
      if (v_11573 == 1) v_24860 <= v_24861;
      if (v_12009 == 1) v_24866 <= v_24867;
      if (v_12221 == 1) v_24872 <= v_24873;
      if (v_12321 == 1) v_24878 <= v_24879;
      if (v_12365 == 1) v_24884 <= v_24885;
      if (v_12328 == 1) v_24892 <= v_24893;
      if (v_12228 == 1) v_24900 <= v_24901;
      if (v_12272 == 1) v_24906 <= v_24907;
      if (v_12235 == 1) v_24914 <= v_24915;
      if (v_12016 == 1) v_24922 <= v_24923;
      if (v_12116 == 1) v_24928 <= v_24929;
      if (v_12160 == 1) v_24934 <= v_24935;
      if (v_12123 == 1) v_24942 <= v_24943;
      if (v_12023 == 1) v_24950 <= v_24951;
      if (v_12067 == 1) v_24956 <= v_24957;
      if (v_12030 == 1) v_24964 <= v_24965;
      if (v_11580 == 1) v_24972 <= v_24973;
      if (v_11792 == 1) v_24978 <= v_24979;
      if (v_11892 == 1) v_24984 <= v_24985;
      if (v_11936 == 1) v_24990 <= v_24991;
      if (v_11899 == 1) v_24998 <= v_24999;
      if (v_11799 == 1) v_25006 <= v_25007;
      if (v_11843 == 1) v_25012 <= v_25013;
      if (v_11806 == 1) v_25020 <= v_25021;
      if (v_11587 == 1) v_25028 <= v_25029;
      if (v_11687 == 1) v_25034 <= v_25035;
      if (v_11731 == 1) v_25040 <= v_25041;
      if (v_11694 == 1) v_25048 <= v_25049;
      if (v_11594 == 1) v_25056 <= v_25057;
      if (v_11638 == 1) v_25062 <= v_25063;
      if (v_11601 == 1) v_25070 <= v_25071;
      if (v_7994 == 1) v_25078 <= v_25079;
      if (v_9774 == 1) v_25084 <= v_25085;
      if (v_10658 == 1) v_25090 <= v_25091;
      if (v_11094 == 1) v_25096 <= v_25097;
      if (v_11306 == 1) v_25102 <= v_25103;
      if (v_11406 == 1) v_25108 <= v_25109;
      if (v_11450 == 1) v_25114 <= v_25115;
      if (v_11413 == 1) v_25122 <= v_25123;
      if (v_11313 == 1) v_25130 <= v_25131;
      if (v_11357 == 1) v_25136 <= v_25137;
      if (v_11320 == 1) v_25144 <= v_25145;
      if (v_11101 == 1) v_25152 <= v_25153;
      if (v_11201 == 1) v_25158 <= v_25159;
      if (v_11245 == 1) v_25164 <= v_25165;
      if (v_11208 == 1) v_25172 <= v_25173;
      if (v_11108 == 1) v_25180 <= v_25181;
      if (v_11152 == 1) v_25186 <= v_25187;
      if (v_11115 == 1) v_25194 <= v_25195;
      if (v_10665 == 1) v_25202 <= v_25203;
      if (v_10877 == 1) v_25208 <= v_25209;
      if (v_10977 == 1) v_25214 <= v_25215;
      if (v_11021 == 1) v_25220 <= v_25221;
      if (v_10984 == 1) v_25228 <= v_25229;
      if (v_10884 == 1) v_25236 <= v_25237;
      if (v_10928 == 1) v_25242 <= v_25243;
      if (v_10891 == 1) v_25250 <= v_25251;
      if (v_10672 == 1) v_25258 <= v_25259;
      if (v_10772 == 1) v_25264 <= v_25265;
      if (v_10816 == 1) v_25270 <= v_25271;
      if (v_10779 == 1) v_25278 <= v_25279;
      if (v_10679 == 1) v_25286 <= v_25287;
      if (v_10723 == 1) v_25292 <= v_25293;
      if (v_10686 == 1) v_25300 <= v_25301;
      if (v_9781 == 1) v_25308 <= v_25309;
      if (v_10217 == 1) v_25314 <= v_25315;
      if (v_10429 == 1) v_25320 <= v_25321;
      if (v_10529 == 1) v_25326 <= v_25327;
      if (v_10573 == 1) v_25332 <= v_25333;
      if (v_10536 == 1) v_25340 <= v_25341;
      if (v_10436 == 1) v_25348 <= v_25349;
      if (v_10480 == 1) v_25354 <= v_25355;
      if (v_10443 == 1) v_25362 <= v_25363;
      if (v_10224 == 1) v_25370 <= v_25371;
      if (v_10324 == 1) v_25376 <= v_25377;
      if (v_10368 == 1) v_25382 <= v_25383;
      if (v_10331 == 1) v_25390 <= v_25391;
      if (v_10231 == 1) v_25398 <= v_25399;
      if (v_10275 == 1) v_25404 <= v_25405;
      if (v_10238 == 1) v_25412 <= v_25413;
      if (v_9788 == 1) v_25420 <= v_25421;
      if (v_10000 == 1) v_25426 <= v_25427;
      if (v_10100 == 1) v_25432 <= v_25433;
      if (v_10144 == 1) v_25438 <= v_25439;
      if (v_10107 == 1) v_25446 <= v_25447;
      if (v_10007 == 1) v_25454 <= v_25455;
      if (v_10051 == 1) v_25460 <= v_25461;
      if (v_10014 == 1) v_25468 <= v_25469;
      if (v_9795 == 1) v_25476 <= v_25477;
      if (v_9895 == 1) v_25482 <= v_25483;
      if (v_9939 == 1) v_25488 <= v_25489;
      if (v_9902 == 1) v_25496 <= v_25497;
      if (v_9802 == 1) v_25504 <= v_25505;
      if (v_9846 == 1) v_25510 <= v_25511;
      if (v_9809 == 1) v_25518 <= v_25519;
      if (v_8001 == 1) v_25526 <= v_25527;
      if (v_8885 == 1) v_25532 <= v_25533;
      if (v_9321 == 1) v_25538 <= v_25539;
      if (v_9533 == 1) v_25544 <= v_25545;
      if (v_9633 == 1) v_25550 <= v_25551;
      if (v_9677 == 1) v_25556 <= v_25557;
      if (v_9640 == 1) v_25564 <= v_25565;
      if (v_9540 == 1) v_25572 <= v_25573;
      if (v_9584 == 1) v_25578 <= v_25579;
      if (v_9547 == 1) v_25586 <= v_25587;
      if (v_9328 == 1) v_25594 <= v_25595;
      if (v_9428 == 1) v_25600 <= v_25601;
      if (v_9472 == 1) v_25606 <= v_25607;
      if (v_9435 == 1) v_25614 <= v_25615;
      if (v_9335 == 1) v_25622 <= v_25623;
      if (v_9379 == 1) v_25628 <= v_25629;
      if (v_9342 == 1) v_25636 <= v_25637;
      if (v_8892 == 1) v_25644 <= v_25645;
      if (v_9104 == 1) v_25650 <= v_25651;
      if (v_9204 == 1) v_25656 <= v_25657;
      if (v_9248 == 1) v_25662 <= v_25663;
      if (v_9211 == 1) v_25670 <= v_25671;
      if (v_9111 == 1) v_25678 <= v_25679;
      if (v_9155 == 1) v_25684 <= v_25685;
      if (v_9118 == 1) v_25692 <= v_25693;
      if (v_8899 == 1) v_25700 <= v_25701;
      if (v_8999 == 1) v_25706 <= v_25707;
      if (v_9043 == 1) v_25712 <= v_25713;
      if (v_9006 == 1) v_25720 <= v_25721;
      if (v_8906 == 1) v_25728 <= v_25729;
      if (v_8950 == 1) v_25734 <= v_25735;
      if (v_8913 == 1) v_25742 <= v_25743;
      if (v_8008 == 1) v_25750 <= v_25751;
      if (v_8444 == 1) v_25756 <= v_25757;
      if (v_8656 == 1) v_25762 <= v_25763;
      if (v_8756 == 1) v_25768 <= v_25769;
      if (v_8800 == 1) v_25774 <= v_25775;
      if (v_8763 == 1) v_25782 <= v_25783;
      if (v_8663 == 1) v_25790 <= v_25791;
      if (v_8707 == 1) v_25796 <= v_25797;
      if (v_8670 == 1) v_25804 <= v_25805;
      if (v_8451 == 1) v_25812 <= v_25813;
      if (v_8551 == 1) v_25818 <= v_25819;
      if (v_8595 == 1) v_25824 <= v_25825;
      if (v_8558 == 1) v_25832 <= v_25833;
      if (v_8458 == 1) v_25840 <= v_25841;
      if (v_8502 == 1) v_25846 <= v_25847;
      if (v_8465 == 1) v_25854 <= v_25855;
      if (v_8015 == 1) v_25862 <= v_25863;
      if (v_8227 == 1) v_25868 <= v_25869;
      if (v_8327 == 1) v_25874 <= v_25875;
      if (v_8371 == 1) v_25880 <= v_25881;
      if (v_8334 == 1) v_25888 <= v_25889;
      if (v_8234 == 1) v_25896 <= v_25897;
      if (v_8278 == 1) v_25902 <= v_25903;
      if (v_8241 == 1) v_25910 <= v_25911;
      if (v_8022 == 1) v_25918 <= v_25919;
      if (v_8122 == 1) v_25924 <= v_25925;
      if (v_8166 == 1) v_25930 <= v_25931;
      if (v_8129 == 1) v_25938 <= v_25939;
      if (v_8029 == 1) v_25946 <= v_25947;
      if (v_8073 == 1) v_25952 <= v_25953;
      if (v_8036 == 1) v_25960 <= v_25961;
      if (v_7959 == 1) v_25968 <= v_25969;
      if (v_4387 == 1) v_25974 <= v_25975;
      if (v_2607 == 1) v_25980 <= v_25981;
      if (v_847 == 1) v_25986 <= v_25987;
      if (v_854 == 1) v_25992 <= v_25993;
      if (v_1290 == 1) v_25998 <= v_25999;
      if (v_1502 == 1) v_26004 <= v_26005;
      if (v_1602 == 1) v_26010 <= v_26011;
      if (v_1646 == 1) v_26016 <= v_26017;
      if (v_1609 == 1) v_26024 <= v_26025;
      if (v_1509 == 1) v_26032 <= v_26033;
      if (v_1553 == 1) v_26038 <= v_26039;
      if (v_1516 == 1) v_26046 <= v_26047;
      if (v_1297 == 1) v_26054 <= v_26055;
      if (v_1397 == 1) v_26060 <= v_26061;
      if (v_1441 == 1) v_26066 <= v_26067;
      if (v_1404 == 1) v_26074 <= v_26075;
      if (v_1304 == 1) v_26082 <= v_26083;
      if (v_1348 == 1) v_26088 <= v_26089;
      if (v_1311 == 1) v_26096 <= v_26097;
      if (v_861 == 1) v_26104 <= v_26105;
      if (v_1073 == 1) v_26110 <= v_26111;
      if (v_1173 == 1) v_26116 <= v_26117;
      if (v_1217 == 1) v_26122 <= v_26123;
      if (v_1180 == 1) v_26130 <= v_26131;
      if (v_1080 == 1) v_26138 <= v_26139;
      if (v_1124 == 1) v_26144 <= v_26145;
      if (v_1087 == 1) v_26152 <= v_26153;
      if (v_868 == 1) v_26160 <= v_26161;
      if (v_968 == 1) v_26166 <= v_26167;
      if (v_1012 == 1) v_26172 <= v_26173;
      if (v_975 == 1) v_26180 <= v_26181;
      if (v_875 == 1) v_26188 <= v_26189;
      if (v_919 == 1) v_26194 <= v_26195;
      if (v_882 == 1) v_26202 <= v_26203;
      if (v_405 == 1) v_26210 <= v_26211;
      if (v_412 == 1) v_26216 <= v_26217;
      if (v_624 == 1) v_26222 <= v_26223;
      if (v_724 == 1) v_26228 <= v_26229;
      if (v_768 == 1) v_26234 <= v_26235;
      if (v_731 == 1) v_26242 <= v_26243;
      if (v_631 == 1) v_26250 <= v_26251;
      if (v_675 == 1) v_26256 <= v_26257;
      if (v_638 == 1) v_26264 <= v_26265;
      if (v_419 == 1) v_26272 <= v_26273;
      if (v_519 == 1) v_26278 <= v_26279;
      if (v_563 == 1) v_26284 <= v_26285;
      if (v_526 == 1) v_26292 <= v_26293;
      if (v_426 == 1) v_26300 <= v_26301;
      if (v_470 == 1) v_26306 <= v_26307;
      if (v_433 == 1) v_26314 <= v_26315;
      if (v_187 == 1) v_26322 <= v_26323;
      if (v_194 == 1) v_26328 <= v_26329;
      if (v_294 == 1) v_26334 <= v_26335;
      if (v_338 == 1) v_26340 <= v_26341;
      if (v_301 == 1) v_26348 <= v_26349;
      if (v_201 == 1) v_26356 <= v_26357;
      if (v_245 == 1) v_26362 <= v_26363;
      if (v_208 == 1) v_26370 <= v_26371;
      if (v_81 == 1) v_26378 <= v_26379;
      if (v_88 == 1) v_26384 <= v_26385;
      if (v_132 == 1) v_26390 <= v_26391;
      if (v_95 == 1) v_26398 <= v_26399;
      if (v_31 == 1) v_26406 <= v_26407;
      if (v_38 == 1) v_26412 <= v_26413;
      if (v_9 == 1) v_26420 <= v_26421;
      if (v_1736 == 1) v_26428 <= v_26429;
      if (v_2172 == 1) v_26434 <= v_26435;
      if (v_2384 == 1) v_26440 <= v_26441;
      if (v_2484 == 1) v_26446 <= v_26447;
      if (v_2528 == 1) v_26452 <= v_26453;
      if (v_2491 == 1) v_26460 <= v_26461;
      if (v_2391 == 1) v_26468 <= v_26469;
      if (v_2435 == 1) v_26474 <= v_26475;
      if (v_2398 == 1) v_26482 <= v_26483;
      if (v_2179 == 1) v_26490 <= v_26491;
      if (v_2279 == 1) v_26496 <= v_26497;
      if (v_2323 == 1) v_26502 <= v_26503;
      if (v_2286 == 1) v_26510 <= v_26511;
      if (v_2186 == 1) v_26518 <= v_26519;
      if (v_2230 == 1) v_26524 <= v_26525;
      if (v_2193 == 1) v_26532 <= v_26533;
      if (v_1743 == 1) v_26540 <= v_26541;
      if (v_1955 == 1) v_26546 <= v_26547;
      if (v_2055 == 1) v_26552 <= v_26553;
      if (v_2099 == 1) v_26558 <= v_26559;
      if (v_2062 == 1) v_26566 <= v_26567;
      if (v_1962 == 1) v_26574 <= v_26575;
      if (v_2006 == 1) v_26580 <= v_26581;
      if (v_1969 == 1) v_26588 <= v_26589;
      if (v_1750 == 1) v_26596 <= v_26597;
      if (v_1850 == 1) v_26602 <= v_26603;
      if (v_1894 == 1) v_26608 <= v_26609;
      if (v_1857 == 1) v_26616 <= v_26617;
      if (v_1757 == 1) v_26624 <= v_26625;
      if (v_1801 == 1) v_26630 <= v_26631;
      if (v_1764 == 1) v_26638 <= v_26639;
      if (v_2620 == 1) v_26646 <= v_26647;
      if (v_3504 == 1) v_26652 <= v_26653;
      if (v_3940 == 1) v_26658 <= v_26659;
      if (v_4152 == 1) v_26664 <= v_26665;
      if (v_4252 == 1) v_26670 <= v_26671;
      if (v_4296 == 1) v_26676 <= v_26677;
      if (v_4259 == 1) v_26684 <= v_26685;
      if (v_4159 == 1) v_26692 <= v_26693;
      if (v_4203 == 1) v_26698 <= v_26699;
      if (v_4166 == 1) v_26706 <= v_26707;
      if (v_3947 == 1) v_26714 <= v_26715;
      if (v_4047 == 1) v_26720 <= v_26721;
      if (v_4091 == 1) v_26726 <= v_26727;
      if (v_4054 == 1) v_26734 <= v_26735;
      if (v_3954 == 1) v_26742 <= v_26743;
      if (v_3998 == 1) v_26748 <= v_26749;
      if (v_3961 == 1) v_26756 <= v_26757;
      if (v_3511 == 1) v_26764 <= v_26765;
      if (v_3723 == 1) v_26770 <= v_26771;
      if (v_3823 == 1) v_26776 <= v_26777;
      if (v_3867 == 1) v_26782 <= v_26783;
      if (v_3830 == 1) v_26790 <= v_26791;
      if (v_3730 == 1) v_26798 <= v_26799;
      if (v_3774 == 1) v_26804 <= v_26805;
      if (v_3737 == 1) v_26812 <= v_26813;
      if (v_3518 == 1) v_26820 <= v_26821;
      if (v_3618 == 1) v_26826 <= v_26827;
      if (v_3662 == 1) v_26832 <= v_26833;
      if (v_3625 == 1) v_26840 <= v_26841;
      if (v_3525 == 1) v_26848 <= v_26849;
      if (v_3569 == 1) v_26854 <= v_26855;
      if (v_3532 == 1) v_26862 <= v_26863;
      if (v_2627 == 1) v_26870 <= v_26871;
      if (v_3063 == 1) v_26876 <= v_26877;
      if (v_3275 == 1) v_26882 <= v_26883;
      if (v_3375 == 1) v_26888 <= v_26889;
      if (v_3419 == 1) v_26894 <= v_26895;
      if (v_3382 == 1) v_26902 <= v_26903;
      if (v_3282 == 1) v_26910 <= v_26911;
      if (v_3326 == 1) v_26916 <= v_26917;
      if (v_3289 == 1) v_26924 <= v_26925;
      if (v_3070 == 1) v_26932 <= v_26933;
      if (v_3170 == 1) v_26938 <= v_26939;
      if (v_3214 == 1) v_26944 <= v_26945;
      if (v_3177 == 1) v_26952 <= v_26953;
      if (v_3077 == 1) v_26960 <= v_26961;
      if (v_3121 == 1) v_26966 <= v_26967;
      if (v_3084 == 1) v_26974 <= v_26975;
      if (v_2634 == 1) v_26982 <= v_26983;
      if (v_2846 == 1) v_26988 <= v_26989;
      if (v_2946 == 1) v_26994 <= v_26995;
      if (v_2990 == 1) v_27000 <= v_27001;
      if (v_2953 == 1) v_27008 <= v_27009;
      if (v_2853 == 1) v_27016 <= v_27017;
      if (v_2897 == 1) v_27022 <= v_27023;
      if (v_2860 == 1) v_27030 <= v_27031;
      if (v_2641 == 1) v_27038 <= v_27039;
      if (v_2741 == 1) v_27044 <= v_27045;
      if (v_2785 == 1) v_27050 <= v_27051;
      if (v_2748 == 1) v_27058 <= v_27059;
      if (v_2648 == 1) v_27066 <= v_27067;
      if (v_2692 == 1) v_27072 <= v_27073;
      if (v_2655 == 1) v_27080 <= v_27081;
      if (v_4400 == 1) v_27088 <= v_27089;
      if (v_6180 == 1) v_27094 <= v_27095;
      if (v_7064 == 1) v_27100 <= v_27101;
      if (v_7500 == 1) v_27106 <= v_27107;
      if (v_7712 == 1) v_27112 <= v_27113;
      if (v_7812 == 1) v_27118 <= v_27119;
      if (v_7856 == 1) v_27124 <= v_27125;
      if (v_7819 == 1) v_27132 <= v_27133;
      if (v_7719 == 1) v_27140 <= v_27141;
      if (v_7763 == 1) v_27146 <= v_27147;
      if (v_7726 == 1) v_27154 <= v_27155;
      if (v_7507 == 1) v_27162 <= v_27163;
      if (v_7607 == 1) v_27168 <= v_27169;
      if (v_7651 == 1) v_27174 <= v_27175;
      if (v_7614 == 1) v_27182 <= v_27183;
      if (v_7514 == 1) v_27190 <= v_27191;
      if (v_7558 == 1) v_27196 <= v_27197;
      if (v_7521 == 1) v_27204 <= v_27205;
      if (v_7071 == 1) v_27212 <= v_27213;
      if (v_7283 == 1) v_27218 <= v_27219;
      if (v_7383 == 1) v_27224 <= v_27225;
      if (v_7427 == 1) v_27230 <= v_27231;
      if (v_7390 == 1) v_27238 <= v_27239;
      if (v_7290 == 1) v_27246 <= v_27247;
      if (v_7334 == 1) v_27252 <= v_27253;
      if (v_7297 == 1) v_27260 <= v_27261;
      if (v_7078 == 1) v_27268 <= v_27269;
      if (v_7178 == 1) v_27274 <= v_27275;
      if (v_7222 == 1) v_27280 <= v_27281;
      if (v_7185 == 1) v_27288 <= v_27289;
      if (v_7085 == 1) v_27296 <= v_27297;
      if (v_7129 == 1) v_27302 <= v_27303;
      if (v_7092 == 1) v_27310 <= v_27311;
      if (v_6187 == 1) v_27318 <= v_27319;
      if (v_6623 == 1) v_27324 <= v_27325;
      if (v_6835 == 1) v_27330 <= v_27331;
      if (v_6935 == 1) v_27336 <= v_27337;
      if (v_6979 == 1) v_27342 <= v_27343;
      if (v_6942 == 1) v_27350 <= v_27351;
      if (v_6842 == 1) v_27358 <= v_27359;
      if (v_6886 == 1) v_27364 <= v_27365;
      if (v_6849 == 1) v_27372 <= v_27373;
      if (v_6630 == 1) v_27380 <= v_27381;
      if (v_6730 == 1) v_27386 <= v_27387;
      if (v_6774 == 1) v_27392 <= v_27393;
      if (v_6737 == 1) v_27400 <= v_27401;
      if (v_6637 == 1) v_27408 <= v_27409;
      if (v_6681 == 1) v_27414 <= v_27415;
      if (v_6644 == 1) v_27422 <= v_27423;
      if (v_6194 == 1) v_27430 <= v_27431;
      if (v_6406 == 1) v_27436 <= v_27437;
      if (v_6506 == 1) v_27442 <= v_27443;
      if (v_6550 == 1) v_27448 <= v_27449;
      if (v_6513 == 1) v_27456 <= v_27457;
      if (v_6413 == 1) v_27464 <= v_27465;
      if (v_6457 == 1) v_27470 <= v_27471;
      if (v_6420 == 1) v_27478 <= v_27479;
      if (v_6201 == 1) v_27486 <= v_27487;
      if (v_6301 == 1) v_27492 <= v_27493;
      if (v_6345 == 1) v_27498 <= v_27499;
      if (v_6308 == 1) v_27506 <= v_27507;
      if (v_6208 == 1) v_27514 <= v_27515;
      if (v_6252 == 1) v_27520 <= v_27521;
      if (v_6215 == 1) v_27528 <= v_27529;
      if (v_4407 == 1) v_27536 <= v_27537;
      if (v_5291 == 1) v_27542 <= v_27543;
      if (v_5727 == 1) v_27548 <= v_27549;
      if (v_5939 == 1) v_27554 <= v_27555;
      if (v_6039 == 1) v_27560 <= v_27561;
      if (v_6083 == 1) v_27566 <= v_27567;
      if (v_6046 == 1) v_27574 <= v_27575;
      if (v_5946 == 1) v_27582 <= v_27583;
      if (v_5990 == 1) v_27588 <= v_27589;
      if (v_5953 == 1) v_27596 <= v_27597;
      if (v_5734 == 1) v_27604 <= v_27605;
      if (v_5834 == 1) v_27610 <= v_27611;
      if (v_5878 == 1) v_27616 <= v_27617;
      if (v_5841 == 1) v_27624 <= v_27625;
      if (v_5741 == 1) v_27632 <= v_27633;
      if (v_5785 == 1) v_27638 <= v_27639;
      if (v_5748 == 1) v_27646 <= v_27647;
      if (v_5298 == 1) v_27654 <= v_27655;
      if (v_5510 == 1) v_27660 <= v_27661;
      if (v_5610 == 1) v_27666 <= v_27667;
      if (v_5654 == 1) v_27672 <= v_27673;
      if (v_5617 == 1) v_27680 <= v_27681;
      if (v_5517 == 1) v_27688 <= v_27689;
      if (v_5561 == 1) v_27694 <= v_27695;
      if (v_5524 == 1) v_27702 <= v_27703;
      if (v_5305 == 1) v_27710 <= v_27711;
      if (v_5405 == 1) v_27716 <= v_27717;
      if (v_5449 == 1) v_27722 <= v_27723;
      if (v_5412 == 1) v_27730 <= v_27731;
      if (v_5312 == 1) v_27738 <= v_27739;
      if (v_5356 == 1) v_27744 <= v_27745;
      if (v_5319 == 1) v_27752 <= v_27753;
      if (v_4414 == 1) v_27760 <= v_27761;
      if (v_4850 == 1) v_27766 <= v_27767;
      if (v_5062 == 1) v_27772 <= v_27773;
      if (v_5162 == 1) v_27778 <= v_27779;
      if (v_5206 == 1) v_27784 <= v_27785;
      if (v_5169 == 1) v_27792 <= v_27793;
      if (v_5069 == 1) v_27800 <= v_27801;
      if (v_5113 == 1) v_27806 <= v_27807;
      if (v_5076 == 1) v_27814 <= v_27815;
      if (v_4857 == 1) v_27822 <= v_27823;
      if (v_4957 == 1) v_27828 <= v_27829;
      if (v_5001 == 1) v_27834 <= v_27835;
      if (v_4964 == 1) v_27842 <= v_27843;
      if (v_4864 == 1) v_27850 <= v_27851;
      if (v_4908 == 1) v_27856 <= v_27857;
      if (v_4871 == 1) v_27864 <= v_27865;
      if (v_4421 == 1) v_27872 <= v_27873;
      if (v_4633 == 1) v_27878 <= v_27879;
      if (v_4733 == 1) v_27884 <= v_27885;
      if (v_4777 == 1) v_27890 <= v_27891;
      if (v_4740 == 1) v_27898 <= v_27899;
      if (v_4640 == 1) v_27906 <= v_27907;
      if (v_4684 == 1) v_27912 <= v_27913;
      if (v_4647 == 1) v_27920 <= v_27921;
      if (v_4428 == 1) v_27928 <= v_27929;
      if (v_4528 == 1) v_27934 <= v_27935;
      if (v_4572 == 1) v_27940 <= v_27941;
      if (v_4535 == 1) v_27948 <= v_27949;
      if (v_4435 == 1) v_27956 <= v_27957;
      if (v_4479 == 1) v_27962 <= v_27963;
      if (v_4442 == 1) v_27970 <= v_27971;
    end
  end
endmodule