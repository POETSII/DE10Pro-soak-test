module Pebbles
  (input wire clock,
   input wire reset,
   input wire [0:0] out_consume_en,
   input wire [0:0] in0_canPeek,
   input wire [7:0] in0_peek,
   output wire [0:0] in0_consume_en,
   output wire [0:0] out_canPeek,
   output wire [7:0] out_peek);
  // Declarations
  //////////////////////////////////////////////////////////////////////////////
  wire [0:0] v_0;
  wire [0:0] v_1;
  function [0:0] mux_1(input [0:0] sel);
    case (sel) 0: mux_1 = 1'h0; 1: mux_1 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2;
  wire [0:0] vin0_consume_en_3;
  wire [0:0] vout_canPeek_3;
  wire [7:0] vout_peek_3;
  wire [0:0] v_4;
  function [0:0] mux_4(input [0:0] sel);
    case (sel) 0: mux_4 = 1'h0; 1: mux_4 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5;
  wire [0:0] v_6;
  wire [0:0] v_7;
  function [0:0] mux_7(input [0:0] sel);
    case (sel) 0: mux_7 = 1'h0; 1: mux_7 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8;
  wire [0:0] v_9;
  wire [0:0] v_10;
  wire [0:0] vin0_consume_en_11;
  wire [0:0] vout_canPeek_11;
  wire [7:0] vout_peek_11;
  wire [0:0] v_12;
  function [0:0] mux_12(input [0:0] sel);
    case (sel) 0: mux_12 = 1'h0; 1: mux_12 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_13;
  wire [0:0] v_14;
  wire [0:0] v_15;
  function [0:0] mux_15(input [0:0] sel);
    case (sel) 0: mux_15 = 1'h0; 1: mux_15 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_16;
  wire [0:0] vin0_consume_en_17;
  wire [0:0] vout_canPeek_17;
  wire [7:0] vout_peek_17;
  wire [0:0] v_18;
  function [0:0] mux_18(input [0:0] sel);
    case (sel) 0: mux_18 = 1'h0; 1: mux_18 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_19;
  wire [0:0] v_20;
  wire [0:0] v_21;
  function [0:0] mux_21(input [0:0] sel);
    case (sel) 0: mux_21 = 1'h0; 1: mux_21 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_22;
  wire [0:0] v_23;
  wire [0:0] v_24;
  wire [0:0] vin0_consume_en_25;
  wire [0:0] vout_canPeek_25;
  wire [7:0] vout_peek_25;
  wire [0:0] v_26;
  function [0:0] mux_26(input [0:0] sel);
    case (sel) 0: mux_26 = 1'h0; 1: mux_26 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_27;
  wire [0:0] v_28;
  wire [0:0] v_29;
  function [0:0] mux_29(input [0:0] sel);
    case (sel) 0: mux_29 = 1'h0; 1: mux_29 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_30;
  wire [0:0] vin0_consume_en_31;
  wire [0:0] vout_canPeek_31;
  wire [7:0] vout_peek_31;
  wire [0:0] v_32;
  function [0:0] mux_32(input [0:0] sel);
    case (sel) 0: mux_32 = 1'h0; 1: mux_32 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_33;
  wire [0:0] v_34;
  wire [0:0] v_35;
  function [0:0] mux_35(input [0:0] sel);
    case (sel) 0: mux_35 = 1'h0; 1: mux_35 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_36;
  wire [0:0] v_37;
  wire [0:0] v_38;
  wire [0:0] vin0_consume_en_39;
  wire [0:0] vout_canPeek_39;
  wire [7:0] vout_peek_39;
  wire [0:0] v_40;
  function [0:0] mux_40(input [0:0] sel);
    case (sel) 0: mux_40 = 1'h0; 1: mux_40 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_41;
  wire [0:0] v_42;
  wire [0:0] v_43;
  function [0:0] mux_43(input [0:0] sel);
    case (sel) 0: mux_43 = 1'h0; 1: mux_43 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_44;
  wire [0:0] vin0_consume_en_45;
  wire [0:0] vout_canPeek_45;
  wire [7:0] vout_peek_45;
  wire [0:0] v_46;
  function [0:0] mux_46(input [0:0] sel);
    case (sel) 0: mux_46 = 1'h0; 1: mux_46 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_47;
  wire [0:0] v_48;
  wire [0:0] v_49;
  function [0:0] mux_49(input [0:0] sel);
    case (sel) 0: mux_49 = 1'h0; 1: mux_49 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_50;
  wire [0:0] v_51;
  wire [0:0] v_52;
  wire [0:0] vin0_consume_en_53;
  wire [0:0] vout_canPeek_53;
  wire [7:0] vout_peek_53;
  wire [0:0] v_54;
  function [0:0] mux_54(input [0:0] sel);
    case (sel) 0: mux_54 = 1'h0; 1: mux_54 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_55;
  wire [0:0] v_56;
  wire [0:0] v_57;
  function [0:0] mux_57(input [0:0] sel);
    case (sel) 0: mux_57 = 1'h0; 1: mux_57 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_58;
  wire [0:0] vin0_consume_en_59;
  wire [0:0] vout_canPeek_59;
  wire [7:0] vout_peek_59;
  wire [0:0] v_60;
  function [0:0] mux_60(input [0:0] sel);
    case (sel) 0: mux_60 = 1'h0; 1: mux_60 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_61;
  wire [0:0] v_62;
  wire [0:0] v_63;
  function [0:0] mux_63(input [0:0] sel);
    case (sel) 0: mux_63 = 1'h0; 1: mux_63 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_64;
  wire [0:0] v_65;
  wire [0:0] v_66;
  wire [0:0] vin0_consume_en_67;
  wire [0:0] vout_canPeek_67;
  wire [7:0] vout_peek_67;
  wire [0:0] v_68;
  function [0:0] mux_68(input [0:0] sel);
    case (sel) 0: mux_68 = 1'h0; 1: mux_68 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_69;
  wire [0:0] v_70;
  wire [0:0] v_71;
  function [0:0] mux_71(input [0:0] sel);
    case (sel) 0: mux_71 = 1'h0; 1: mux_71 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_72;
  wire [0:0] vin0_consume_en_73;
  wire [0:0] vout_canPeek_73;
  wire [7:0] vout_peek_73;
  wire [0:0] v_74;
  function [0:0] mux_74(input [0:0] sel);
    case (sel) 0: mux_74 = 1'h0; 1: mux_74 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_75;
  wire [0:0] v_76;
  wire [0:0] v_77;
  function [0:0] mux_77(input [0:0] sel);
    case (sel) 0: mux_77 = 1'h0; 1: mux_77 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_78;
  wire [0:0] v_79;
  wire [0:0] v_80;
  wire [0:0] vin0_consume_en_81;
  wire [0:0] vout_canPeek_81;
  wire [7:0] vout_peek_81;
  wire [0:0] v_82;
  function [0:0] mux_82(input [0:0] sel);
    case (sel) 0: mux_82 = 1'h0; 1: mux_82 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_83;
  wire [0:0] v_84;
  wire [0:0] v_85;
  function [0:0] mux_85(input [0:0] sel);
    case (sel) 0: mux_85 = 1'h0; 1: mux_85 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_86;
  wire [0:0] vin0_consume_en_87;
  wire [0:0] vout_canPeek_87;
  wire [7:0] vout_peek_87;
  wire [0:0] v_88;
  function [0:0] mux_88(input [0:0] sel);
    case (sel) 0: mux_88 = 1'h0; 1: mux_88 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_89;
  wire [0:0] v_90;
  wire [0:0] v_91;
  function [0:0] mux_91(input [0:0] sel);
    case (sel) 0: mux_91 = 1'h0; 1: mux_91 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_92;
  wire [0:0] v_93;
  wire [0:0] v_94;
  wire [0:0] vin0_consume_en_95;
  wire [0:0] vout_canPeek_95;
  wire [7:0] vout_peek_95;
  wire [0:0] v_96;
  function [0:0] mux_96(input [0:0] sel);
    case (sel) 0: mux_96 = 1'h0; 1: mux_96 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_97;
  wire [0:0] v_98;
  wire [0:0] v_99;
  function [0:0] mux_99(input [0:0] sel);
    case (sel) 0: mux_99 = 1'h0; 1: mux_99 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_100;
  wire [0:0] vin0_consume_en_101;
  wire [0:0] vout_canPeek_101;
  wire [7:0] vout_peek_101;
  wire [0:0] v_102;
  function [0:0] mux_102(input [0:0] sel);
    case (sel) 0: mux_102 = 1'h0; 1: mux_102 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_103;
  wire [0:0] v_104;
  wire [0:0] v_105;
  function [0:0] mux_105(input [0:0] sel);
    case (sel) 0: mux_105 = 1'h0; 1: mux_105 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_106;
  wire [0:0] v_107;
  wire [0:0] v_108;
  wire [0:0] vin0_consume_en_109;
  wire [0:0] vout_canPeek_109;
  wire [7:0] vout_peek_109;
  wire [0:0] v_110;
  function [0:0] mux_110(input [0:0] sel);
    case (sel) 0: mux_110 = 1'h0; 1: mux_110 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_111;
  wire [0:0] v_112;
  wire [0:0] v_113;
  function [0:0] mux_113(input [0:0] sel);
    case (sel) 0: mux_113 = 1'h0; 1: mux_113 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_114;
  wire [0:0] vin0_consume_en_115;
  wire [0:0] vout_canPeek_115;
  wire [7:0] vout_peek_115;
  wire [0:0] v_116;
  function [0:0] mux_116(input [0:0] sel);
    case (sel) 0: mux_116 = 1'h0; 1: mux_116 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_117;
  wire [0:0] v_118;
  wire [0:0] v_119;
  function [0:0] mux_119(input [0:0] sel);
    case (sel) 0: mux_119 = 1'h0; 1: mux_119 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_120;
  wire [0:0] v_121;
  wire [0:0] v_122;
  wire [0:0] vin0_consume_en_123;
  wire [0:0] vout_canPeek_123;
  wire [7:0] vout_peek_123;
  wire [0:0] v_124;
  function [0:0] mux_124(input [0:0] sel);
    case (sel) 0: mux_124 = 1'h0; 1: mux_124 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_125;
  wire [0:0] v_126;
  wire [0:0] v_127;
  function [0:0] mux_127(input [0:0] sel);
    case (sel) 0: mux_127 = 1'h0; 1: mux_127 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_128;
  wire [0:0] vin0_consume_en_129;
  wire [0:0] vout_canPeek_129;
  wire [7:0] vout_peek_129;
  wire [0:0] v_130;
  function [0:0] mux_130(input [0:0] sel);
    case (sel) 0: mux_130 = 1'h0; 1: mux_130 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_131;
  wire [0:0] v_132;
  wire [0:0] v_133;
  function [0:0] mux_133(input [0:0] sel);
    case (sel) 0: mux_133 = 1'h0; 1: mux_133 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_134;
  wire [0:0] v_135;
  wire [0:0] v_136;
  wire [0:0] vin0_consume_en_137;
  wire [0:0] vout_canPeek_137;
  wire [7:0] vout_peek_137;
  wire [0:0] v_138;
  function [0:0] mux_138(input [0:0] sel);
    case (sel) 0: mux_138 = 1'h0; 1: mux_138 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_139;
  wire [0:0] v_140;
  wire [0:0] v_141;
  function [0:0] mux_141(input [0:0] sel);
    case (sel) 0: mux_141 = 1'h0; 1: mux_141 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_142;
  wire [0:0] vin0_consume_en_143;
  wire [0:0] vout_canPeek_143;
  wire [7:0] vout_peek_143;
  wire [0:0] v_144;
  function [0:0] mux_144(input [0:0] sel);
    case (sel) 0: mux_144 = 1'h0; 1: mux_144 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_145;
  wire [0:0] v_146;
  wire [0:0] v_147;
  function [0:0] mux_147(input [0:0] sel);
    case (sel) 0: mux_147 = 1'h0; 1: mux_147 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_148;
  wire [0:0] v_149;
  wire [0:0] v_150;
  wire [0:0] vin0_consume_en_151;
  wire [0:0] vout_canPeek_151;
  wire [7:0] vout_peek_151;
  wire [0:0] v_152;
  function [0:0] mux_152(input [0:0] sel);
    case (sel) 0: mux_152 = 1'h0; 1: mux_152 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_153;
  wire [0:0] v_154;
  wire [0:0] v_155;
  function [0:0] mux_155(input [0:0] sel);
    case (sel) 0: mux_155 = 1'h0; 1: mux_155 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_156;
  wire [0:0] vin0_consume_en_157;
  wire [0:0] vout_canPeek_157;
  wire [7:0] vout_peek_157;
  wire [0:0] v_158;
  function [0:0] mux_158(input [0:0] sel);
    case (sel) 0: mux_158 = 1'h0; 1: mux_158 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_159;
  wire [0:0] v_160;
  wire [0:0] v_161;
  function [0:0] mux_161(input [0:0] sel);
    case (sel) 0: mux_161 = 1'h0; 1: mux_161 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_162;
  wire [0:0] v_163;
  wire [0:0] v_164;
  wire [0:0] vin0_consume_en_165;
  wire [0:0] vout_canPeek_165;
  wire [7:0] vout_peek_165;
  wire [0:0] v_166;
  function [0:0] mux_166(input [0:0] sel);
    case (sel) 0: mux_166 = 1'h0; 1: mux_166 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_167;
  wire [0:0] v_168;
  wire [0:0] v_169;
  function [0:0] mux_169(input [0:0] sel);
    case (sel) 0: mux_169 = 1'h0; 1: mux_169 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_170;
  wire [0:0] vin0_consume_en_171;
  wire [0:0] vout_canPeek_171;
  wire [7:0] vout_peek_171;
  wire [0:0] v_172;
  function [0:0] mux_172(input [0:0] sel);
    case (sel) 0: mux_172 = 1'h0; 1: mux_172 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_173;
  wire [0:0] v_174;
  wire [0:0] v_175;
  function [0:0] mux_175(input [0:0] sel);
    case (sel) 0: mux_175 = 1'h0; 1: mux_175 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_176;
  wire [0:0] v_177;
  wire [0:0] v_178;
  wire [0:0] vin0_consume_en_179;
  wire [0:0] vout_canPeek_179;
  wire [7:0] vout_peek_179;
  wire [0:0] v_180;
  function [0:0] mux_180(input [0:0] sel);
    case (sel) 0: mux_180 = 1'h0; 1: mux_180 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_181;
  wire [0:0] v_182;
  wire [0:0] v_183;
  function [0:0] mux_183(input [0:0] sel);
    case (sel) 0: mux_183 = 1'h0; 1: mux_183 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_184;
  wire [0:0] vin0_consume_en_185;
  wire [0:0] vout_canPeek_185;
  wire [7:0] vout_peek_185;
  wire [0:0] v_186;
  function [0:0] mux_186(input [0:0] sel);
    case (sel) 0: mux_186 = 1'h0; 1: mux_186 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_187;
  wire [0:0] v_188;
  wire [0:0] v_189;
  function [0:0] mux_189(input [0:0] sel);
    case (sel) 0: mux_189 = 1'h0; 1: mux_189 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_190;
  wire [0:0] v_191;
  wire [0:0] v_192;
  wire [0:0] vin0_consume_en_193;
  wire [0:0] vout_canPeek_193;
  wire [7:0] vout_peek_193;
  wire [0:0] v_194;
  function [0:0] mux_194(input [0:0] sel);
    case (sel) 0: mux_194 = 1'h0; 1: mux_194 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_195;
  wire [0:0] v_196;
  wire [0:0] v_197;
  function [0:0] mux_197(input [0:0] sel);
    case (sel) 0: mux_197 = 1'h0; 1: mux_197 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_198;
  wire [0:0] vin0_consume_en_199;
  wire [0:0] vout_canPeek_199;
  wire [7:0] vout_peek_199;
  wire [0:0] v_200;
  function [0:0] mux_200(input [0:0] sel);
    case (sel) 0: mux_200 = 1'h0; 1: mux_200 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_201;
  wire [0:0] v_202;
  wire [0:0] v_203;
  function [0:0] mux_203(input [0:0] sel);
    case (sel) 0: mux_203 = 1'h0; 1: mux_203 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_204;
  wire [0:0] v_205;
  wire [0:0] v_206;
  wire [0:0] vin0_consume_en_207;
  wire [0:0] vout_canPeek_207;
  wire [7:0] vout_peek_207;
  wire [0:0] v_208;
  function [0:0] mux_208(input [0:0] sel);
    case (sel) 0: mux_208 = 1'h0; 1: mux_208 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_209;
  wire [0:0] v_210;
  wire [0:0] v_211;
  function [0:0] mux_211(input [0:0] sel);
    case (sel) 0: mux_211 = 1'h0; 1: mux_211 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_212;
  wire [0:0] vin0_consume_en_213;
  wire [0:0] vout_canPeek_213;
  wire [7:0] vout_peek_213;
  wire [0:0] v_214;
  function [0:0] mux_214(input [0:0] sel);
    case (sel) 0: mux_214 = 1'h0; 1: mux_214 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_215;
  wire [0:0] v_216;
  wire [0:0] v_217;
  function [0:0] mux_217(input [0:0] sel);
    case (sel) 0: mux_217 = 1'h0; 1: mux_217 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_218;
  wire [0:0] v_219;
  wire [0:0] v_220;
  wire [0:0] vin0_consume_en_221;
  wire [0:0] vout_canPeek_221;
  wire [7:0] vout_peek_221;
  wire [0:0] v_222;
  function [0:0] mux_222(input [0:0] sel);
    case (sel) 0: mux_222 = 1'h0; 1: mux_222 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_223;
  wire [0:0] v_224;
  wire [0:0] v_225;
  function [0:0] mux_225(input [0:0] sel);
    case (sel) 0: mux_225 = 1'h0; 1: mux_225 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_226;
  wire [0:0] vin0_consume_en_227;
  wire [0:0] vout_canPeek_227;
  wire [7:0] vout_peek_227;
  wire [0:0] v_228;
  function [0:0] mux_228(input [0:0] sel);
    case (sel) 0: mux_228 = 1'h0; 1: mux_228 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_229;
  wire [0:0] v_230;
  wire [0:0] v_231;
  function [0:0] mux_231(input [0:0] sel);
    case (sel) 0: mux_231 = 1'h0; 1: mux_231 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_232;
  wire [0:0] v_233;
  wire [0:0] v_234;
  wire [0:0] vin0_consume_en_235;
  wire [0:0] vout_canPeek_235;
  wire [7:0] vout_peek_235;
  wire [0:0] v_236;
  function [0:0] mux_236(input [0:0] sel);
    case (sel) 0: mux_236 = 1'h0; 1: mux_236 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_237;
  wire [0:0] v_238;
  wire [0:0] v_239;
  function [0:0] mux_239(input [0:0] sel);
    case (sel) 0: mux_239 = 1'h0; 1: mux_239 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_240;
  wire [0:0] vin0_consume_en_241;
  wire [0:0] vout_canPeek_241;
  wire [7:0] vout_peek_241;
  wire [0:0] v_242;
  function [0:0] mux_242(input [0:0] sel);
    case (sel) 0: mux_242 = 1'h0; 1: mux_242 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_243;
  wire [0:0] v_244;
  wire [0:0] v_245;
  function [0:0] mux_245(input [0:0] sel);
    case (sel) 0: mux_245 = 1'h0; 1: mux_245 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_246;
  wire [0:0] v_247;
  wire [0:0] v_248;
  wire [0:0] vin0_consume_en_249;
  wire [0:0] vout_canPeek_249;
  wire [7:0] vout_peek_249;
  wire [0:0] v_250;
  function [0:0] mux_250(input [0:0] sel);
    case (sel) 0: mux_250 = 1'h0; 1: mux_250 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_251;
  wire [0:0] v_252;
  wire [0:0] v_253;
  function [0:0] mux_253(input [0:0] sel);
    case (sel) 0: mux_253 = 1'h0; 1: mux_253 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_254;
  wire [0:0] vin0_consume_en_255;
  wire [0:0] vout_canPeek_255;
  wire [7:0] vout_peek_255;
  wire [0:0] v_256;
  function [0:0] mux_256(input [0:0] sel);
    case (sel) 0: mux_256 = 1'h0; 1: mux_256 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_257;
  wire [0:0] v_258;
  wire [0:0] v_259;
  function [0:0] mux_259(input [0:0] sel);
    case (sel) 0: mux_259 = 1'h0; 1: mux_259 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_260;
  wire [0:0] v_261;
  wire [0:0] v_262;
  wire [0:0] vin0_consume_en_263;
  wire [0:0] vout_canPeek_263;
  wire [7:0] vout_peek_263;
  wire [0:0] v_264;
  function [0:0] mux_264(input [0:0] sel);
    case (sel) 0: mux_264 = 1'h0; 1: mux_264 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_265;
  wire [0:0] v_266;
  wire [0:0] v_267;
  function [0:0] mux_267(input [0:0] sel);
    case (sel) 0: mux_267 = 1'h0; 1: mux_267 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_268;
  wire [0:0] vin0_consume_en_269;
  wire [0:0] vout_canPeek_269;
  wire [7:0] vout_peek_269;
  wire [0:0] v_270;
  function [0:0] mux_270(input [0:0] sel);
    case (sel) 0: mux_270 = 1'h0; 1: mux_270 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_271;
  wire [0:0] v_272;
  wire [0:0] v_273;
  function [0:0] mux_273(input [0:0] sel);
    case (sel) 0: mux_273 = 1'h0; 1: mux_273 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_274;
  wire [0:0] v_275;
  wire [0:0] v_276;
  wire [0:0] vin0_consume_en_277;
  wire [0:0] vout_canPeek_277;
  wire [7:0] vout_peek_277;
  wire [0:0] v_278;
  function [0:0] mux_278(input [0:0] sel);
    case (sel) 0: mux_278 = 1'h0; 1: mux_278 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_279;
  wire [0:0] v_280;
  wire [0:0] v_281;
  function [0:0] mux_281(input [0:0] sel);
    case (sel) 0: mux_281 = 1'h0; 1: mux_281 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_282;
  wire [0:0] vin0_consume_en_283;
  wire [0:0] vout_canPeek_283;
  wire [7:0] vout_peek_283;
  wire [0:0] v_284;
  function [0:0] mux_284(input [0:0] sel);
    case (sel) 0: mux_284 = 1'h0; 1: mux_284 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_285;
  wire [0:0] v_286;
  wire [0:0] v_287;
  function [0:0] mux_287(input [0:0] sel);
    case (sel) 0: mux_287 = 1'h0; 1: mux_287 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_288;
  wire [0:0] v_289;
  wire [0:0] v_290;
  wire [0:0] vin0_consume_en_291;
  wire [0:0] vout_canPeek_291;
  wire [7:0] vout_peek_291;
  wire [0:0] v_292;
  function [0:0] mux_292(input [0:0] sel);
    case (sel) 0: mux_292 = 1'h0; 1: mux_292 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_293;
  wire [0:0] v_294;
  wire [0:0] v_295;
  function [0:0] mux_295(input [0:0] sel);
    case (sel) 0: mux_295 = 1'h0; 1: mux_295 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_296;
  wire [0:0] vin0_consume_en_297;
  wire [0:0] vout_canPeek_297;
  wire [7:0] vout_peek_297;
  wire [0:0] v_298;
  function [0:0] mux_298(input [0:0] sel);
    case (sel) 0: mux_298 = 1'h0; 1: mux_298 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_299;
  wire [0:0] v_300;
  wire [0:0] v_301;
  function [0:0] mux_301(input [0:0] sel);
    case (sel) 0: mux_301 = 1'h0; 1: mux_301 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_302;
  wire [0:0] v_303;
  wire [0:0] v_304;
  wire [0:0] vin0_consume_en_305;
  wire [0:0] vout_canPeek_305;
  wire [7:0] vout_peek_305;
  wire [0:0] v_306;
  function [0:0] mux_306(input [0:0] sel);
    case (sel) 0: mux_306 = 1'h0; 1: mux_306 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_307;
  wire [0:0] v_308;
  wire [0:0] v_309;
  function [0:0] mux_309(input [0:0] sel);
    case (sel) 0: mux_309 = 1'h0; 1: mux_309 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_310;
  wire [0:0] vin0_consume_en_311;
  wire [0:0] vout_canPeek_311;
  wire [7:0] vout_peek_311;
  wire [0:0] v_312;
  function [0:0] mux_312(input [0:0] sel);
    case (sel) 0: mux_312 = 1'h0; 1: mux_312 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_313;
  wire [0:0] v_314;
  wire [0:0] v_315;
  function [0:0] mux_315(input [0:0] sel);
    case (sel) 0: mux_315 = 1'h0; 1: mux_315 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_316;
  wire [0:0] v_317;
  wire [0:0] v_318;
  wire [0:0] vin0_consume_en_319;
  wire [0:0] vout_canPeek_319;
  wire [7:0] vout_peek_319;
  wire [0:0] v_320;
  function [0:0] mux_320(input [0:0] sel);
    case (sel) 0: mux_320 = 1'h0; 1: mux_320 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_321;
  wire [0:0] v_322;
  wire [0:0] v_323;
  function [0:0] mux_323(input [0:0] sel);
    case (sel) 0: mux_323 = 1'h0; 1: mux_323 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_324;
  wire [0:0] vin0_consume_en_325;
  wire [0:0] vout_canPeek_325;
  wire [7:0] vout_peek_325;
  wire [0:0] v_326;
  function [0:0] mux_326(input [0:0] sel);
    case (sel) 0: mux_326 = 1'h0; 1: mux_326 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_327;
  wire [0:0] v_328;
  wire [0:0] v_329;
  function [0:0] mux_329(input [0:0] sel);
    case (sel) 0: mux_329 = 1'h0; 1: mux_329 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_330;
  wire [0:0] v_331;
  wire [0:0] v_332;
  wire [0:0] vin0_consume_en_333;
  wire [0:0] vout_canPeek_333;
  wire [7:0] vout_peek_333;
  wire [0:0] v_334;
  function [0:0] mux_334(input [0:0] sel);
    case (sel) 0: mux_334 = 1'h0; 1: mux_334 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_335;
  wire [0:0] v_336;
  wire [0:0] v_337;
  function [0:0] mux_337(input [0:0] sel);
    case (sel) 0: mux_337 = 1'h0; 1: mux_337 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_338;
  wire [0:0] vin0_consume_en_339;
  wire [0:0] vout_canPeek_339;
  wire [7:0] vout_peek_339;
  wire [0:0] v_340;
  function [0:0] mux_340(input [0:0] sel);
    case (sel) 0: mux_340 = 1'h0; 1: mux_340 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_341;
  wire [0:0] v_342;
  wire [0:0] v_343;
  function [0:0] mux_343(input [0:0] sel);
    case (sel) 0: mux_343 = 1'h0; 1: mux_343 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_344;
  wire [0:0] v_345;
  wire [0:0] v_346;
  wire [0:0] vin0_consume_en_347;
  wire [0:0] vout_canPeek_347;
  wire [7:0] vout_peek_347;
  wire [0:0] v_348;
  function [0:0] mux_348(input [0:0] sel);
    case (sel) 0: mux_348 = 1'h0; 1: mux_348 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_349;
  wire [0:0] v_350;
  wire [0:0] v_351;
  function [0:0] mux_351(input [0:0] sel);
    case (sel) 0: mux_351 = 1'h0; 1: mux_351 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_352;
  wire [0:0] vin0_consume_en_353;
  wire [0:0] vout_canPeek_353;
  wire [7:0] vout_peek_353;
  wire [0:0] v_354;
  function [0:0] mux_354(input [0:0] sel);
    case (sel) 0: mux_354 = 1'h0; 1: mux_354 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_355;
  wire [0:0] v_356;
  wire [0:0] v_357;
  function [0:0] mux_357(input [0:0] sel);
    case (sel) 0: mux_357 = 1'h0; 1: mux_357 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_358;
  wire [0:0] v_359;
  wire [0:0] v_360;
  wire [0:0] vin0_consume_en_361;
  wire [0:0] vout_canPeek_361;
  wire [7:0] vout_peek_361;
  wire [0:0] v_362;
  function [0:0] mux_362(input [0:0] sel);
    case (sel) 0: mux_362 = 1'h0; 1: mux_362 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_363;
  wire [0:0] v_364;
  wire [0:0] v_365;
  function [0:0] mux_365(input [0:0] sel);
    case (sel) 0: mux_365 = 1'h0; 1: mux_365 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_366;
  wire [0:0] vin0_consume_en_367;
  wire [0:0] vout_canPeek_367;
  wire [7:0] vout_peek_367;
  wire [0:0] v_368;
  function [0:0] mux_368(input [0:0] sel);
    case (sel) 0: mux_368 = 1'h0; 1: mux_368 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_369;
  wire [0:0] v_370;
  wire [0:0] v_371;
  function [0:0] mux_371(input [0:0] sel);
    case (sel) 0: mux_371 = 1'h0; 1: mux_371 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_372;
  wire [0:0] v_373;
  wire [0:0] v_374;
  wire [0:0] vin0_consume_en_375;
  wire [0:0] vout_canPeek_375;
  wire [7:0] vout_peek_375;
  wire [0:0] v_376;
  function [0:0] mux_376(input [0:0] sel);
    case (sel) 0: mux_376 = 1'h0; 1: mux_376 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_377;
  wire [0:0] v_378;
  wire [0:0] v_379;
  function [0:0] mux_379(input [0:0] sel);
    case (sel) 0: mux_379 = 1'h0; 1: mux_379 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_380;
  wire [0:0] vin0_consume_en_381;
  wire [0:0] vout_canPeek_381;
  wire [7:0] vout_peek_381;
  wire [0:0] v_382;
  function [0:0] mux_382(input [0:0] sel);
    case (sel) 0: mux_382 = 1'h0; 1: mux_382 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_383;
  wire [0:0] v_384;
  wire [0:0] v_385;
  function [0:0] mux_385(input [0:0] sel);
    case (sel) 0: mux_385 = 1'h0; 1: mux_385 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_386;
  wire [0:0] v_387;
  wire [0:0] v_388;
  wire [0:0] vin0_consume_en_389;
  wire [0:0] vout_canPeek_389;
  wire [7:0] vout_peek_389;
  wire [0:0] v_390;
  function [0:0] mux_390(input [0:0] sel);
    case (sel) 0: mux_390 = 1'h0; 1: mux_390 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_391;
  wire [0:0] v_392;
  wire [0:0] v_393;
  function [0:0] mux_393(input [0:0] sel);
    case (sel) 0: mux_393 = 1'h0; 1: mux_393 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_394;
  wire [0:0] vin0_consume_en_395;
  wire [0:0] vout_canPeek_395;
  wire [7:0] vout_peek_395;
  wire [0:0] v_396;
  function [0:0] mux_396(input [0:0] sel);
    case (sel) 0: mux_396 = 1'h0; 1: mux_396 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_397;
  wire [0:0] v_398;
  wire [0:0] v_399;
  function [0:0] mux_399(input [0:0] sel);
    case (sel) 0: mux_399 = 1'h0; 1: mux_399 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_400;
  wire [0:0] v_401;
  wire [0:0] v_402;
  wire [0:0] vin0_consume_en_403;
  wire [0:0] vout_canPeek_403;
  wire [7:0] vout_peek_403;
  wire [0:0] v_404;
  function [0:0] mux_404(input [0:0] sel);
    case (sel) 0: mux_404 = 1'h0; 1: mux_404 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_405;
  wire [0:0] v_406;
  wire [0:0] v_407;
  function [0:0] mux_407(input [0:0] sel);
    case (sel) 0: mux_407 = 1'h0; 1: mux_407 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_408;
  wire [0:0] vin0_consume_en_409;
  wire [0:0] vout_canPeek_409;
  wire [7:0] vout_peek_409;
  wire [0:0] v_410;
  function [0:0] mux_410(input [0:0] sel);
    case (sel) 0: mux_410 = 1'h0; 1: mux_410 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_411;
  wire [0:0] v_412;
  wire [0:0] v_413;
  function [0:0] mux_413(input [0:0] sel);
    case (sel) 0: mux_413 = 1'h0; 1: mux_413 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_414;
  wire [0:0] v_415;
  wire [0:0] v_416;
  wire [0:0] vin0_consume_en_417;
  wire [0:0] vout_canPeek_417;
  wire [7:0] vout_peek_417;
  wire [0:0] v_418;
  function [0:0] mux_418(input [0:0] sel);
    case (sel) 0: mux_418 = 1'h0; 1: mux_418 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_419;
  wire [0:0] v_420;
  wire [0:0] v_421;
  function [0:0] mux_421(input [0:0] sel);
    case (sel) 0: mux_421 = 1'h0; 1: mux_421 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_422;
  wire [0:0] vin0_consume_en_423;
  wire [0:0] vout_canPeek_423;
  wire [7:0] vout_peek_423;
  wire [0:0] v_424;
  function [0:0] mux_424(input [0:0] sel);
    case (sel) 0: mux_424 = 1'h0; 1: mux_424 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_425;
  wire [0:0] v_426;
  wire [0:0] v_427;
  function [0:0] mux_427(input [0:0] sel);
    case (sel) 0: mux_427 = 1'h0; 1: mux_427 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_428;
  wire [0:0] v_429;
  wire [0:0] v_430;
  wire [0:0] vin0_consume_en_431;
  wire [0:0] vout_canPeek_431;
  wire [7:0] vout_peek_431;
  wire [0:0] v_432;
  function [0:0] mux_432(input [0:0] sel);
    case (sel) 0: mux_432 = 1'h0; 1: mux_432 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_433;
  wire [0:0] v_434;
  wire [0:0] v_435;
  function [0:0] mux_435(input [0:0] sel);
    case (sel) 0: mux_435 = 1'h0; 1: mux_435 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_436;
  wire [0:0] vin0_consume_en_437;
  wire [0:0] vout_canPeek_437;
  wire [7:0] vout_peek_437;
  wire [0:0] v_438;
  function [0:0] mux_438(input [0:0] sel);
    case (sel) 0: mux_438 = 1'h0; 1: mux_438 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_439;
  wire [0:0] v_440;
  wire [0:0] v_441;
  function [0:0] mux_441(input [0:0] sel);
    case (sel) 0: mux_441 = 1'h0; 1: mux_441 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_442;
  wire [0:0] v_443;
  wire [0:0] v_444;
  wire [0:0] vin0_consume_en_445;
  wire [0:0] vout_canPeek_445;
  wire [7:0] vout_peek_445;
  wire [0:0] v_446;
  function [0:0] mux_446(input [0:0] sel);
    case (sel) 0: mux_446 = 1'h0; 1: mux_446 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_447;
  wire [0:0] v_448;
  wire [0:0] v_449;
  function [0:0] mux_449(input [0:0] sel);
    case (sel) 0: mux_449 = 1'h0; 1: mux_449 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_450;
  wire [0:0] vin0_consume_en_451;
  wire [0:0] vout_canPeek_451;
  wire [7:0] vout_peek_451;
  wire [0:0] v_452;
  function [0:0] mux_452(input [0:0] sel);
    case (sel) 0: mux_452 = 1'h0; 1: mux_452 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_453;
  wire [0:0] v_454;
  wire [0:0] v_455;
  function [0:0] mux_455(input [0:0] sel);
    case (sel) 0: mux_455 = 1'h0; 1: mux_455 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_456;
  wire [0:0] v_457;
  wire [0:0] v_458;
  wire [0:0] vin0_consume_en_459;
  wire [0:0] vout_canPeek_459;
  wire [7:0] vout_peek_459;
  wire [0:0] v_460;
  function [0:0] mux_460(input [0:0] sel);
    case (sel) 0: mux_460 = 1'h0; 1: mux_460 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_461;
  wire [0:0] v_462;
  wire [0:0] v_463;
  function [0:0] mux_463(input [0:0] sel);
    case (sel) 0: mux_463 = 1'h0; 1: mux_463 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_464;
  wire [0:0] vin0_consume_en_465;
  wire [0:0] vout_canPeek_465;
  wire [7:0] vout_peek_465;
  wire [0:0] v_466;
  function [0:0] mux_466(input [0:0] sel);
    case (sel) 0: mux_466 = 1'h0; 1: mux_466 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_467;
  wire [0:0] v_468;
  wire [0:0] v_469;
  function [0:0] mux_469(input [0:0] sel);
    case (sel) 0: mux_469 = 1'h0; 1: mux_469 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_470;
  wire [0:0] v_471;
  wire [0:0] v_472;
  wire [0:0] vin0_consume_en_473;
  wire [0:0] vout_canPeek_473;
  wire [7:0] vout_peek_473;
  wire [0:0] v_474;
  function [0:0] mux_474(input [0:0] sel);
    case (sel) 0: mux_474 = 1'h0; 1: mux_474 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_475;
  wire [0:0] v_476;
  wire [0:0] v_477;
  function [0:0] mux_477(input [0:0] sel);
    case (sel) 0: mux_477 = 1'h0; 1: mux_477 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_478;
  wire [0:0] vin0_consume_en_479;
  wire [0:0] vout_canPeek_479;
  wire [7:0] vout_peek_479;
  wire [0:0] v_480;
  function [0:0] mux_480(input [0:0] sel);
    case (sel) 0: mux_480 = 1'h0; 1: mux_480 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_481;
  wire [0:0] v_482;
  wire [0:0] v_483;
  function [0:0] mux_483(input [0:0] sel);
    case (sel) 0: mux_483 = 1'h0; 1: mux_483 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_484;
  wire [0:0] v_485;
  wire [0:0] v_486;
  wire [0:0] vin0_consume_en_487;
  wire [0:0] vout_canPeek_487;
  wire [7:0] vout_peek_487;
  wire [0:0] v_488;
  function [0:0] mux_488(input [0:0] sel);
    case (sel) 0: mux_488 = 1'h0; 1: mux_488 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_489;
  wire [0:0] v_490;
  wire [0:0] v_491;
  function [0:0] mux_491(input [0:0] sel);
    case (sel) 0: mux_491 = 1'h0; 1: mux_491 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_492;
  wire [0:0] vin0_consume_en_493;
  wire [0:0] vout_canPeek_493;
  wire [7:0] vout_peek_493;
  wire [0:0] v_494;
  function [0:0] mux_494(input [0:0] sel);
    case (sel) 0: mux_494 = 1'h0; 1: mux_494 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_495;
  wire [0:0] v_496;
  wire [0:0] v_497;
  function [0:0] mux_497(input [0:0] sel);
    case (sel) 0: mux_497 = 1'h0; 1: mux_497 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_498;
  wire [0:0] v_499;
  wire [0:0] v_500;
  wire [0:0] vin0_consume_en_501;
  wire [0:0] vout_canPeek_501;
  wire [7:0] vout_peek_501;
  wire [0:0] v_502;
  function [0:0] mux_502(input [0:0] sel);
    case (sel) 0: mux_502 = 1'h0; 1: mux_502 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_503;
  wire [0:0] v_504;
  wire [0:0] v_505;
  function [0:0] mux_505(input [0:0] sel);
    case (sel) 0: mux_505 = 1'h0; 1: mux_505 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_506;
  wire [0:0] vin0_consume_en_507;
  wire [0:0] vout_canPeek_507;
  wire [7:0] vout_peek_507;
  wire [0:0] v_508;
  function [0:0] mux_508(input [0:0] sel);
    case (sel) 0: mux_508 = 1'h0; 1: mux_508 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_509;
  wire [0:0] v_510;
  wire [0:0] v_511;
  function [0:0] mux_511(input [0:0] sel);
    case (sel) 0: mux_511 = 1'h0; 1: mux_511 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_512;
  wire [0:0] v_513;
  wire [0:0] v_514;
  wire [0:0] vin0_consume_en_515;
  wire [0:0] vout_canPeek_515;
  wire [7:0] vout_peek_515;
  wire [0:0] v_516;
  function [0:0] mux_516(input [0:0] sel);
    case (sel) 0: mux_516 = 1'h0; 1: mux_516 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_517;
  wire [0:0] v_518;
  wire [0:0] v_519;
  function [0:0] mux_519(input [0:0] sel);
    case (sel) 0: mux_519 = 1'h0; 1: mux_519 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_520;
  wire [0:0] vin0_consume_en_521;
  wire [0:0] vout_canPeek_521;
  wire [7:0] vout_peek_521;
  wire [0:0] v_522;
  function [0:0] mux_522(input [0:0] sel);
    case (sel) 0: mux_522 = 1'h0; 1: mux_522 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_523;
  wire [0:0] v_524;
  wire [0:0] v_525;
  function [0:0] mux_525(input [0:0] sel);
    case (sel) 0: mux_525 = 1'h0; 1: mux_525 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_526;
  wire [0:0] v_527;
  wire [0:0] v_528;
  wire [0:0] vin0_consume_en_529;
  wire [0:0] vout_canPeek_529;
  wire [7:0] vout_peek_529;
  wire [0:0] v_530;
  function [0:0] mux_530(input [0:0] sel);
    case (sel) 0: mux_530 = 1'h0; 1: mux_530 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_531;
  wire [0:0] v_532;
  wire [0:0] v_533;
  function [0:0] mux_533(input [0:0] sel);
    case (sel) 0: mux_533 = 1'h0; 1: mux_533 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_534;
  wire [0:0] vin0_consume_en_535;
  wire [0:0] vout_canPeek_535;
  wire [7:0] vout_peek_535;
  wire [0:0] v_536;
  function [0:0] mux_536(input [0:0] sel);
    case (sel) 0: mux_536 = 1'h0; 1: mux_536 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_537;
  wire [0:0] v_538;
  wire [0:0] v_539;
  function [0:0] mux_539(input [0:0] sel);
    case (sel) 0: mux_539 = 1'h0; 1: mux_539 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_540;
  wire [0:0] v_541;
  wire [0:0] v_542;
  wire [0:0] vin0_consume_en_543;
  wire [0:0] vout_canPeek_543;
  wire [7:0] vout_peek_543;
  wire [0:0] v_544;
  function [0:0] mux_544(input [0:0] sel);
    case (sel) 0: mux_544 = 1'h0; 1: mux_544 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_545;
  wire [0:0] v_546;
  wire [0:0] v_547;
  function [0:0] mux_547(input [0:0] sel);
    case (sel) 0: mux_547 = 1'h0; 1: mux_547 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_548;
  wire [0:0] vin0_consume_en_549;
  wire [0:0] vout_canPeek_549;
  wire [7:0] vout_peek_549;
  wire [0:0] v_550;
  function [0:0] mux_550(input [0:0] sel);
    case (sel) 0: mux_550 = 1'h0; 1: mux_550 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_551;
  wire [0:0] v_552;
  wire [0:0] v_553;
  function [0:0] mux_553(input [0:0] sel);
    case (sel) 0: mux_553 = 1'h0; 1: mux_553 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_554;
  wire [0:0] v_555;
  wire [0:0] v_556;
  wire [0:0] vin0_consume_en_557;
  wire [0:0] vout_canPeek_557;
  wire [7:0] vout_peek_557;
  wire [0:0] v_558;
  function [0:0] mux_558(input [0:0] sel);
    case (sel) 0: mux_558 = 1'h0; 1: mux_558 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_559;
  wire [0:0] v_560;
  wire [0:0] v_561;
  function [0:0] mux_561(input [0:0] sel);
    case (sel) 0: mux_561 = 1'h0; 1: mux_561 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_562;
  wire [0:0] vin0_consume_en_563;
  wire [0:0] vout_canPeek_563;
  wire [7:0] vout_peek_563;
  wire [0:0] v_564;
  function [0:0] mux_564(input [0:0] sel);
    case (sel) 0: mux_564 = 1'h0; 1: mux_564 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_565;
  wire [0:0] v_566;
  wire [0:0] v_567;
  function [0:0] mux_567(input [0:0] sel);
    case (sel) 0: mux_567 = 1'h0; 1: mux_567 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_568;
  wire [0:0] v_569;
  wire [0:0] v_570;
  wire [0:0] vin0_consume_en_571;
  wire [0:0] vout_canPeek_571;
  wire [7:0] vout_peek_571;
  wire [0:0] v_572;
  function [0:0] mux_572(input [0:0] sel);
    case (sel) 0: mux_572 = 1'h0; 1: mux_572 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_573;
  wire [0:0] v_574;
  wire [0:0] v_575;
  function [0:0] mux_575(input [0:0] sel);
    case (sel) 0: mux_575 = 1'h0; 1: mux_575 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_576;
  wire [0:0] vin0_consume_en_577;
  wire [0:0] vout_canPeek_577;
  wire [7:0] vout_peek_577;
  wire [0:0] v_578;
  function [0:0] mux_578(input [0:0] sel);
    case (sel) 0: mux_578 = 1'h0; 1: mux_578 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_579;
  wire [0:0] v_580;
  wire [0:0] v_581;
  function [0:0] mux_581(input [0:0] sel);
    case (sel) 0: mux_581 = 1'h0; 1: mux_581 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_582;
  wire [0:0] v_583;
  wire [0:0] v_584;
  wire [0:0] vin0_consume_en_585;
  wire [0:0] vout_canPeek_585;
  wire [7:0] vout_peek_585;
  wire [0:0] v_586;
  function [0:0] mux_586(input [0:0] sel);
    case (sel) 0: mux_586 = 1'h0; 1: mux_586 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_587;
  wire [0:0] v_588;
  wire [0:0] v_589;
  function [0:0] mux_589(input [0:0] sel);
    case (sel) 0: mux_589 = 1'h0; 1: mux_589 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_590;
  wire [0:0] vin0_consume_en_591;
  wire [0:0] vout_canPeek_591;
  wire [7:0] vout_peek_591;
  wire [0:0] v_592;
  function [0:0] mux_592(input [0:0] sel);
    case (sel) 0: mux_592 = 1'h0; 1: mux_592 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_593;
  wire [0:0] v_594;
  wire [0:0] v_595;
  function [0:0] mux_595(input [0:0] sel);
    case (sel) 0: mux_595 = 1'h0; 1: mux_595 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_596;
  wire [0:0] v_597;
  wire [0:0] v_598;
  wire [0:0] vin0_consume_en_599;
  wire [0:0] vout_canPeek_599;
  wire [7:0] vout_peek_599;
  wire [0:0] v_600;
  function [0:0] mux_600(input [0:0] sel);
    case (sel) 0: mux_600 = 1'h0; 1: mux_600 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_601;
  wire [0:0] v_602;
  wire [0:0] v_603;
  function [0:0] mux_603(input [0:0] sel);
    case (sel) 0: mux_603 = 1'h0; 1: mux_603 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_604;
  wire [0:0] vin0_consume_en_605;
  wire [0:0] vout_canPeek_605;
  wire [7:0] vout_peek_605;
  wire [0:0] v_606;
  function [0:0] mux_606(input [0:0] sel);
    case (sel) 0: mux_606 = 1'h0; 1: mux_606 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_607;
  wire [0:0] v_608;
  wire [0:0] v_609;
  function [0:0] mux_609(input [0:0] sel);
    case (sel) 0: mux_609 = 1'h0; 1: mux_609 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_610;
  wire [0:0] v_611;
  wire [0:0] v_612;
  wire [0:0] vin0_consume_en_613;
  wire [0:0] vout_canPeek_613;
  wire [7:0] vout_peek_613;
  wire [0:0] v_614;
  function [0:0] mux_614(input [0:0] sel);
    case (sel) 0: mux_614 = 1'h0; 1: mux_614 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_615;
  wire [0:0] v_616;
  wire [0:0] v_617;
  function [0:0] mux_617(input [0:0] sel);
    case (sel) 0: mux_617 = 1'h0; 1: mux_617 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_618;
  wire [0:0] vin0_consume_en_619;
  wire [0:0] vout_canPeek_619;
  wire [7:0] vout_peek_619;
  wire [0:0] v_620;
  function [0:0] mux_620(input [0:0] sel);
    case (sel) 0: mux_620 = 1'h0; 1: mux_620 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_621;
  wire [0:0] v_622;
  wire [0:0] v_623;
  function [0:0] mux_623(input [0:0] sel);
    case (sel) 0: mux_623 = 1'h0; 1: mux_623 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_624;
  wire [0:0] v_625;
  wire [0:0] v_626;
  wire [0:0] vin0_consume_en_627;
  wire [0:0] vout_canPeek_627;
  wire [7:0] vout_peek_627;
  wire [0:0] v_628;
  function [0:0] mux_628(input [0:0] sel);
    case (sel) 0: mux_628 = 1'h0; 1: mux_628 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_629;
  wire [0:0] v_630;
  wire [0:0] v_631;
  function [0:0] mux_631(input [0:0] sel);
    case (sel) 0: mux_631 = 1'h0; 1: mux_631 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_632;
  wire [0:0] vin0_consume_en_633;
  wire [0:0] vout_canPeek_633;
  wire [7:0] vout_peek_633;
  wire [0:0] v_634;
  function [0:0] mux_634(input [0:0] sel);
    case (sel) 0: mux_634 = 1'h0; 1: mux_634 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_635;
  wire [0:0] v_636;
  wire [0:0] v_637;
  function [0:0] mux_637(input [0:0] sel);
    case (sel) 0: mux_637 = 1'h0; 1: mux_637 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_638;
  wire [0:0] v_639;
  wire [0:0] v_640;
  wire [0:0] vin0_consume_en_641;
  wire [0:0] vout_canPeek_641;
  wire [7:0] vout_peek_641;
  wire [0:0] v_642;
  function [0:0] mux_642(input [0:0] sel);
    case (sel) 0: mux_642 = 1'h0; 1: mux_642 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_643;
  wire [0:0] v_644;
  wire [0:0] v_645;
  function [0:0] mux_645(input [0:0] sel);
    case (sel) 0: mux_645 = 1'h0; 1: mux_645 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_646;
  wire [0:0] vin0_consume_en_647;
  wire [0:0] vout_canPeek_647;
  wire [7:0] vout_peek_647;
  wire [0:0] v_648;
  function [0:0] mux_648(input [0:0] sel);
    case (sel) 0: mux_648 = 1'h0; 1: mux_648 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_649;
  wire [0:0] v_650;
  wire [0:0] v_651;
  function [0:0] mux_651(input [0:0] sel);
    case (sel) 0: mux_651 = 1'h0; 1: mux_651 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_652;
  wire [0:0] v_653;
  wire [0:0] v_654;
  wire [0:0] vin0_consume_en_655;
  wire [0:0] vout_canPeek_655;
  wire [7:0] vout_peek_655;
  wire [0:0] v_656;
  function [0:0] mux_656(input [0:0] sel);
    case (sel) 0: mux_656 = 1'h0; 1: mux_656 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_657;
  wire [0:0] v_658;
  wire [0:0] v_659;
  function [0:0] mux_659(input [0:0] sel);
    case (sel) 0: mux_659 = 1'h0; 1: mux_659 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_660;
  wire [0:0] vin0_consume_en_661;
  wire [0:0] vout_canPeek_661;
  wire [7:0] vout_peek_661;
  wire [0:0] v_662;
  function [0:0] mux_662(input [0:0] sel);
    case (sel) 0: mux_662 = 1'h0; 1: mux_662 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_663;
  wire [0:0] v_664;
  wire [0:0] v_665;
  function [0:0] mux_665(input [0:0] sel);
    case (sel) 0: mux_665 = 1'h0; 1: mux_665 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_666;
  wire [0:0] v_667;
  wire [0:0] v_668;
  wire [0:0] vin0_consume_en_669;
  wire [0:0] vout_canPeek_669;
  wire [7:0] vout_peek_669;
  wire [0:0] v_670;
  function [0:0] mux_670(input [0:0] sel);
    case (sel) 0: mux_670 = 1'h0; 1: mux_670 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_671;
  wire [0:0] v_672;
  wire [0:0] v_673;
  function [0:0] mux_673(input [0:0] sel);
    case (sel) 0: mux_673 = 1'h0; 1: mux_673 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_674;
  wire [0:0] vin0_consume_en_675;
  wire [0:0] vout_canPeek_675;
  wire [7:0] vout_peek_675;
  wire [0:0] v_676;
  function [0:0] mux_676(input [0:0] sel);
    case (sel) 0: mux_676 = 1'h0; 1: mux_676 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_677;
  wire [0:0] v_678;
  wire [0:0] v_679;
  function [0:0] mux_679(input [0:0] sel);
    case (sel) 0: mux_679 = 1'h0; 1: mux_679 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_680;
  wire [0:0] v_681;
  wire [0:0] v_682;
  wire [0:0] vin0_consume_en_683;
  wire [0:0] vout_canPeek_683;
  wire [7:0] vout_peek_683;
  wire [0:0] v_684;
  function [0:0] mux_684(input [0:0] sel);
    case (sel) 0: mux_684 = 1'h0; 1: mux_684 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_685;
  wire [0:0] v_686;
  wire [0:0] v_687;
  function [0:0] mux_687(input [0:0] sel);
    case (sel) 0: mux_687 = 1'h0; 1: mux_687 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_688;
  wire [0:0] vin0_consume_en_689;
  wire [0:0] vout_canPeek_689;
  wire [7:0] vout_peek_689;
  wire [0:0] v_690;
  function [0:0] mux_690(input [0:0] sel);
    case (sel) 0: mux_690 = 1'h0; 1: mux_690 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_691;
  wire [0:0] v_692;
  wire [0:0] v_693;
  function [0:0] mux_693(input [0:0] sel);
    case (sel) 0: mux_693 = 1'h0; 1: mux_693 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_694;
  wire [0:0] v_695;
  wire [0:0] v_696;
  wire [0:0] vin0_consume_en_697;
  wire [0:0] vout_canPeek_697;
  wire [7:0] vout_peek_697;
  wire [0:0] v_698;
  function [0:0] mux_698(input [0:0] sel);
    case (sel) 0: mux_698 = 1'h0; 1: mux_698 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_699;
  wire [0:0] v_700;
  wire [0:0] v_701;
  function [0:0] mux_701(input [0:0] sel);
    case (sel) 0: mux_701 = 1'h0; 1: mux_701 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_702;
  wire [0:0] vin0_consume_en_703;
  wire [0:0] vout_canPeek_703;
  wire [7:0] vout_peek_703;
  wire [0:0] v_704;
  function [0:0] mux_704(input [0:0] sel);
    case (sel) 0: mux_704 = 1'h0; 1: mux_704 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_705;
  wire [0:0] v_706;
  wire [0:0] v_707;
  function [0:0] mux_707(input [0:0] sel);
    case (sel) 0: mux_707 = 1'h0; 1: mux_707 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_708;
  wire [0:0] v_709;
  wire [0:0] v_710;
  wire [0:0] vin0_consume_en_711;
  wire [0:0] vout_canPeek_711;
  wire [7:0] vout_peek_711;
  wire [0:0] v_712;
  function [0:0] mux_712(input [0:0] sel);
    case (sel) 0: mux_712 = 1'h0; 1: mux_712 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_713;
  wire [0:0] v_714;
  wire [0:0] v_715;
  function [0:0] mux_715(input [0:0] sel);
    case (sel) 0: mux_715 = 1'h0; 1: mux_715 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_716;
  wire [0:0] vin0_consume_en_717;
  wire [0:0] vout_canPeek_717;
  wire [7:0] vout_peek_717;
  wire [0:0] v_718;
  function [0:0] mux_718(input [0:0] sel);
    case (sel) 0: mux_718 = 1'h0; 1: mux_718 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_719;
  wire [0:0] v_720;
  wire [0:0] v_721;
  function [0:0] mux_721(input [0:0] sel);
    case (sel) 0: mux_721 = 1'h0; 1: mux_721 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_722;
  wire [0:0] v_723;
  wire [0:0] v_724;
  wire [0:0] vin0_consume_en_725;
  wire [0:0] vout_canPeek_725;
  wire [7:0] vout_peek_725;
  wire [0:0] v_726;
  function [0:0] mux_726(input [0:0] sel);
    case (sel) 0: mux_726 = 1'h0; 1: mux_726 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_727;
  wire [0:0] v_728;
  wire [0:0] v_729;
  function [0:0] mux_729(input [0:0] sel);
    case (sel) 0: mux_729 = 1'h0; 1: mux_729 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_730;
  wire [0:0] vin0_consume_en_731;
  wire [0:0] vout_canPeek_731;
  wire [7:0] vout_peek_731;
  wire [0:0] v_732;
  function [0:0] mux_732(input [0:0] sel);
    case (sel) 0: mux_732 = 1'h0; 1: mux_732 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_733;
  wire [0:0] v_734;
  wire [0:0] v_735;
  function [0:0] mux_735(input [0:0] sel);
    case (sel) 0: mux_735 = 1'h0; 1: mux_735 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_736;
  wire [0:0] v_737;
  wire [0:0] v_738;
  wire [0:0] vin0_consume_en_739;
  wire [0:0] vout_canPeek_739;
  wire [7:0] vout_peek_739;
  wire [0:0] v_740;
  function [0:0] mux_740(input [0:0] sel);
    case (sel) 0: mux_740 = 1'h0; 1: mux_740 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_741;
  wire [0:0] v_742;
  wire [0:0] v_743;
  function [0:0] mux_743(input [0:0] sel);
    case (sel) 0: mux_743 = 1'h0; 1: mux_743 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_744;
  wire [0:0] vin0_consume_en_745;
  wire [0:0] vout_canPeek_745;
  wire [7:0] vout_peek_745;
  wire [0:0] v_746;
  function [0:0] mux_746(input [0:0] sel);
    case (sel) 0: mux_746 = 1'h0; 1: mux_746 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_747;
  wire [0:0] v_748;
  wire [0:0] v_749;
  function [0:0] mux_749(input [0:0] sel);
    case (sel) 0: mux_749 = 1'h0; 1: mux_749 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_750;
  wire [0:0] v_751;
  wire [0:0] v_752;
  wire [0:0] vin0_consume_en_753;
  wire [0:0] vout_canPeek_753;
  wire [7:0] vout_peek_753;
  wire [0:0] v_754;
  function [0:0] mux_754(input [0:0] sel);
    case (sel) 0: mux_754 = 1'h0; 1: mux_754 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_755;
  wire [0:0] v_756;
  wire [0:0] v_757;
  function [0:0] mux_757(input [0:0] sel);
    case (sel) 0: mux_757 = 1'h0; 1: mux_757 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_758;
  wire [0:0] vin0_consume_en_759;
  wire [0:0] vout_canPeek_759;
  wire [7:0] vout_peek_759;
  wire [0:0] v_760;
  function [0:0] mux_760(input [0:0] sel);
    case (sel) 0: mux_760 = 1'h0; 1: mux_760 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_761;
  wire [0:0] v_762;
  wire [0:0] v_763;
  function [0:0] mux_763(input [0:0] sel);
    case (sel) 0: mux_763 = 1'h0; 1: mux_763 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_764;
  wire [0:0] v_765;
  wire [0:0] v_766;
  wire [0:0] vin0_consume_en_767;
  wire [0:0] vout_canPeek_767;
  wire [7:0] vout_peek_767;
  wire [0:0] v_768;
  function [0:0] mux_768(input [0:0] sel);
    case (sel) 0: mux_768 = 1'h0; 1: mux_768 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_769;
  wire [0:0] v_770;
  wire [0:0] v_771;
  function [0:0] mux_771(input [0:0] sel);
    case (sel) 0: mux_771 = 1'h0; 1: mux_771 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_772;
  wire [0:0] vin0_consume_en_773;
  wire [0:0] vout_canPeek_773;
  wire [7:0] vout_peek_773;
  wire [0:0] v_774;
  function [0:0] mux_774(input [0:0] sel);
    case (sel) 0: mux_774 = 1'h0; 1: mux_774 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_775;
  wire [0:0] v_776;
  wire [0:0] v_777;
  function [0:0] mux_777(input [0:0] sel);
    case (sel) 0: mux_777 = 1'h0; 1: mux_777 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_778;
  wire [0:0] v_779;
  wire [0:0] v_780;
  wire [0:0] vin0_consume_en_781;
  wire [0:0] vout_canPeek_781;
  wire [7:0] vout_peek_781;
  wire [0:0] v_782;
  function [0:0] mux_782(input [0:0] sel);
    case (sel) 0: mux_782 = 1'h0; 1: mux_782 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_783;
  wire [0:0] v_784;
  wire [0:0] v_785;
  function [0:0] mux_785(input [0:0] sel);
    case (sel) 0: mux_785 = 1'h0; 1: mux_785 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_786;
  wire [0:0] vin0_consume_en_787;
  wire [0:0] vout_canPeek_787;
  wire [7:0] vout_peek_787;
  wire [0:0] v_788;
  function [0:0] mux_788(input [0:0] sel);
    case (sel) 0: mux_788 = 1'h0; 1: mux_788 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_789;
  wire [0:0] v_790;
  wire [0:0] v_791;
  function [0:0] mux_791(input [0:0] sel);
    case (sel) 0: mux_791 = 1'h0; 1: mux_791 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_792;
  wire [0:0] v_793;
  wire [0:0] v_794;
  wire [0:0] vin0_consume_en_795;
  wire [0:0] vout_canPeek_795;
  wire [7:0] vout_peek_795;
  wire [0:0] v_796;
  function [0:0] mux_796(input [0:0] sel);
    case (sel) 0: mux_796 = 1'h0; 1: mux_796 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_797;
  wire [0:0] v_798;
  wire [0:0] v_799;
  function [0:0] mux_799(input [0:0] sel);
    case (sel) 0: mux_799 = 1'h0; 1: mux_799 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_800;
  wire [0:0] vin0_consume_en_801;
  wire [0:0] vout_canPeek_801;
  wire [7:0] vout_peek_801;
  wire [0:0] v_802;
  function [0:0] mux_802(input [0:0] sel);
    case (sel) 0: mux_802 = 1'h0; 1: mux_802 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_803;
  wire [0:0] v_804;
  wire [0:0] v_805;
  function [0:0] mux_805(input [0:0] sel);
    case (sel) 0: mux_805 = 1'h0; 1: mux_805 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_806;
  wire [0:0] v_807;
  wire [0:0] v_808;
  wire [0:0] vin0_consume_en_809;
  wire [0:0] vout_canPeek_809;
  wire [7:0] vout_peek_809;
  wire [0:0] v_810;
  function [0:0] mux_810(input [0:0] sel);
    case (sel) 0: mux_810 = 1'h0; 1: mux_810 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_811;
  wire [0:0] v_812;
  wire [0:0] v_813;
  function [0:0] mux_813(input [0:0] sel);
    case (sel) 0: mux_813 = 1'h0; 1: mux_813 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_814;
  wire [0:0] vin0_consume_en_815;
  wire [0:0] vout_canPeek_815;
  wire [7:0] vout_peek_815;
  wire [0:0] v_816;
  function [0:0] mux_816(input [0:0] sel);
    case (sel) 0: mux_816 = 1'h0; 1: mux_816 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_817;
  wire [0:0] v_818;
  wire [0:0] v_819;
  function [0:0] mux_819(input [0:0] sel);
    case (sel) 0: mux_819 = 1'h0; 1: mux_819 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_820;
  wire [0:0] v_821;
  wire [0:0] v_822;
  wire [0:0] vin0_consume_en_823;
  wire [0:0] vout_canPeek_823;
  wire [7:0] vout_peek_823;
  wire [0:0] v_824;
  function [0:0] mux_824(input [0:0] sel);
    case (sel) 0: mux_824 = 1'h0; 1: mux_824 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_825;
  wire [0:0] v_826;
  wire [0:0] v_827;
  function [0:0] mux_827(input [0:0] sel);
    case (sel) 0: mux_827 = 1'h0; 1: mux_827 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_828;
  wire [0:0] vin0_consume_en_829;
  wire [0:0] vout_canPeek_829;
  wire [7:0] vout_peek_829;
  wire [0:0] v_830;
  function [0:0] mux_830(input [0:0] sel);
    case (sel) 0: mux_830 = 1'h0; 1: mux_830 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_831;
  wire [0:0] v_832;
  wire [0:0] v_833;
  function [0:0] mux_833(input [0:0] sel);
    case (sel) 0: mux_833 = 1'h0; 1: mux_833 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_834;
  wire [0:0] v_835;
  wire [0:0] v_836;
  wire [0:0] vin0_consume_en_837;
  wire [0:0] vout_canPeek_837;
  wire [7:0] vout_peek_837;
  wire [0:0] v_838;
  function [0:0] mux_838(input [0:0] sel);
    case (sel) 0: mux_838 = 1'h0; 1: mux_838 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_839;
  wire [0:0] v_840;
  wire [0:0] v_841;
  function [0:0] mux_841(input [0:0] sel);
    case (sel) 0: mux_841 = 1'h0; 1: mux_841 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_842;
  wire [0:0] vin0_consume_en_843;
  wire [0:0] vout_canPeek_843;
  wire [7:0] vout_peek_843;
  wire [0:0] v_844;
  function [0:0] mux_844(input [0:0] sel);
    case (sel) 0: mux_844 = 1'h0; 1: mux_844 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_845;
  wire [0:0] v_846;
  wire [0:0] v_847;
  function [0:0] mux_847(input [0:0] sel);
    case (sel) 0: mux_847 = 1'h0; 1: mux_847 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_848;
  wire [0:0] v_849;
  wire [0:0] v_850;
  wire [0:0] vin0_consume_en_851;
  wire [0:0] vout_canPeek_851;
  wire [7:0] vout_peek_851;
  wire [0:0] v_852;
  function [0:0] mux_852(input [0:0] sel);
    case (sel) 0: mux_852 = 1'h0; 1: mux_852 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_853;
  wire [0:0] v_854;
  wire [0:0] v_855;
  function [0:0] mux_855(input [0:0] sel);
    case (sel) 0: mux_855 = 1'h0; 1: mux_855 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_856;
  wire [0:0] vin0_consume_en_857;
  wire [0:0] vout_canPeek_857;
  wire [7:0] vout_peek_857;
  wire [0:0] v_858;
  function [0:0] mux_858(input [0:0] sel);
    case (sel) 0: mux_858 = 1'h0; 1: mux_858 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_859;
  wire [0:0] v_860;
  wire [0:0] v_861;
  function [0:0] mux_861(input [0:0] sel);
    case (sel) 0: mux_861 = 1'h0; 1: mux_861 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_862;
  wire [0:0] v_863;
  wire [0:0] v_864;
  wire [0:0] vin0_consume_en_865;
  wire [0:0] vout_canPeek_865;
  wire [7:0] vout_peek_865;
  wire [0:0] v_866;
  function [0:0] mux_866(input [0:0] sel);
    case (sel) 0: mux_866 = 1'h0; 1: mux_866 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_867;
  wire [0:0] v_868;
  wire [0:0] v_869;
  function [0:0] mux_869(input [0:0] sel);
    case (sel) 0: mux_869 = 1'h0; 1: mux_869 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_870;
  wire [0:0] vin0_consume_en_871;
  wire [0:0] vout_canPeek_871;
  wire [7:0] vout_peek_871;
  wire [0:0] v_872;
  function [0:0] mux_872(input [0:0] sel);
    case (sel) 0: mux_872 = 1'h0; 1: mux_872 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_873;
  wire [0:0] v_874;
  wire [0:0] v_875;
  function [0:0] mux_875(input [0:0] sel);
    case (sel) 0: mux_875 = 1'h0; 1: mux_875 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_876;
  wire [0:0] v_877;
  wire [0:0] v_878;
  wire [0:0] vin0_consume_en_879;
  wire [0:0] vout_canPeek_879;
  wire [7:0] vout_peek_879;
  wire [0:0] v_880;
  function [0:0] mux_880(input [0:0] sel);
    case (sel) 0: mux_880 = 1'h0; 1: mux_880 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_881;
  wire [0:0] v_882;
  wire [0:0] v_883;
  function [0:0] mux_883(input [0:0] sel);
    case (sel) 0: mux_883 = 1'h0; 1: mux_883 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_884;
  wire [0:0] vin0_consume_en_885;
  wire [0:0] vout_canPeek_885;
  wire [7:0] vout_peek_885;
  wire [0:0] v_886;
  function [0:0] mux_886(input [0:0] sel);
    case (sel) 0: mux_886 = 1'h0; 1: mux_886 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_887;
  wire [0:0] v_888;
  wire [0:0] v_889;
  function [0:0] mux_889(input [0:0] sel);
    case (sel) 0: mux_889 = 1'h0; 1: mux_889 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_890;
  wire [0:0] v_891;
  wire [0:0] v_892;
  wire [0:0] vin0_consume_en_893;
  wire [0:0] vout_canPeek_893;
  wire [7:0] vout_peek_893;
  wire [0:0] v_894;
  function [0:0] mux_894(input [0:0] sel);
    case (sel) 0: mux_894 = 1'h0; 1: mux_894 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_895;
  wire [0:0] v_896;
  wire [0:0] v_897;
  function [0:0] mux_897(input [0:0] sel);
    case (sel) 0: mux_897 = 1'h0; 1: mux_897 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_898;
  wire [0:0] vin0_consume_en_899;
  wire [0:0] vout_canPeek_899;
  wire [7:0] vout_peek_899;
  wire [0:0] v_900;
  function [0:0] mux_900(input [0:0] sel);
    case (sel) 0: mux_900 = 1'h0; 1: mux_900 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_901;
  wire [0:0] v_902;
  wire [0:0] v_903;
  function [0:0] mux_903(input [0:0] sel);
    case (sel) 0: mux_903 = 1'h0; 1: mux_903 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_904;
  wire [0:0] v_905;
  wire [0:0] v_906;
  wire [0:0] vin0_consume_en_907;
  wire [0:0] vout_canPeek_907;
  wire [7:0] vout_peek_907;
  wire [0:0] v_908;
  function [0:0] mux_908(input [0:0] sel);
    case (sel) 0: mux_908 = 1'h0; 1: mux_908 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_909;
  wire [0:0] v_910;
  wire [0:0] v_911;
  function [0:0] mux_911(input [0:0] sel);
    case (sel) 0: mux_911 = 1'h0; 1: mux_911 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_912;
  wire [0:0] vin0_consume_en_913;
  wire [0:0] vout_canPeek_913;
  wire [7:0] vout_peek_913;
  wire [0:0] v_914;
  function [0:0] mux_914(input [0:0] sel);
    case (sel) 0: mux_914 = 1'h0; 1: mux_914 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_915;
  wire [0:0] v_916;
  wire [0:0] v_917;
  function [0:0] mux_917(input [0:0] sel);
    case (sel) 0: mux_917 = 1'h0; 1: mux_917 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_918;
  wire [0:0] v_919;
  wire [0:0] v_920;
  wire [0:0] vin0_consume_en_921;
  wire [0:0] vout_canPeek_921;
  wire [7:0] vout_peek_921;
  wire [0:0] v_922;
  function [0:0] mux_922(input [0:0] sel);
    case (sel) 0: mux_922 = 1'h0; 1: mux_922 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_923;
  wire [0:0] v_924;
  wire [0:0] v_925;
  function [0:0] mux_925(input [0:0] sel);
    case (sel) 0: mux_925 = 1'h0; 1: mux_925 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_926;
  wire [0:0] vin0_consume_en_927;
  wire [0:0] vout_canPeek_927;
  wire [7:0] vout_peek_927;
  wire [0:0] v_928;
  function [0:0] mux_928(input [0:0] sel);
    case (sel) 0: mux_928 = 1'h0; 1: mux_928 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_929;
  wire [0:0] v_930;
  wire [0:0] v_931;
  function [0:0] mux_931(input [0:0] sel);
    case (sel) 0: mux_931 = 1'h0; 1: mux_931 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_932;
  wire [0:0] v_933;
  wire [0:0] v_934;
  wire [0:0] vin0_consume_en_935;
  wire [0:0] vout_canPeek_935;
  wire [7:0] vout_peek_935;
  wire [0:0] v_936;
  function [0:0] mux_936(input [0:0] sel);
    case (sel) 0: mux_936 = 1'h0; 1: mux_936 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_937;
  wire [0:0] v_938;
  wire [0:0] v_939;
  function [0:0] mux_939(input [0:0] sel);
    case (sel) 0: mux_939 = 1'h0; 1: mux_939 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_940;
  wire [0:0] vin0_consume_en_941;
  wire [0:0] vout_canPeek_941;
  wire [7:0] vout_peek_941;
  wire [0:0] v_942;
  function [0:0] mux_942(input [0:0] sel);
    case (sel) 0: mux_942 = 1'h0; 1: mux_942 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_943;
  wire [0:0] v_944;
  wire [0:0] v_945;
  function [0:0] mux_945(input [0:0] sel);
    case (sel) 0: mux_945 = 1'h0; 1: mux_945 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_946;
  wire [0:0] v_947;
  wire [0:0] v_948;
  wire [0:0] vin0_consume_en_949;
  wire [0:0] vout_canPeek_949;
  wire [7:0] vout_peek_949;
  wire [0:0] v_950;
  function [0:0] mux_950(input [0:0] sel);
    case (sel) 0: mux_950 = 1'h0; 1: mux_950 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_951;
  wire [0:0] v_952;
  wire [0:0] v_953;
  function [0:0] mux_953(input [0:0] sel);
    case (sel) 0: mux_953 = 1'h0; 1: mux_953 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_954;
  wire [0:0] vin0_consume_en_955;
  wire [0:0] vout_canPeek_955;
  wire [7:0] vout_peek_955;
  wire [0:0] v_956;
  function [0:0] mux_956(input [0:0] sel);
    case (sel) 0: mux_956 = 1'h0; 1: mux_956 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_957;
  wire [0:0] v_958;
  wire [0:0] v_959;
  function [0:0] mux_959(input [0:0] sel);
    case (sel) 0: mux_959 = 1'h0; 1: mux_959 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_960;
  wire [0:0] v_961;
  wire [0:0] v_962;
  wire [0:0] vin0_consume_en_963;
  wire [0:0] vout_canPeek_963;
  wire [7:0] vout_peek_963;
  wire [0:0] v_964;
  function [0:0] mux_964(input [0:0] sel);
    case (sel) 0: mux_964 = 1'h0; 1: mux_964 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_965;
  wire [0:0] v_966;
  wire [0:0] v_967;
  function [0:0] mux_967(input [0:0] sel);
    case (sel) 0: mux_967 = 1'h0; 1: mux_967 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_968;
  wire [0:0] vin0_consume_en_969;
  wire [0:0] vout_canPeek_969;
  wire [7:0] vout_peek_969;
  wire [0:0] v_970;
  function [0:0] mux_970(input [0:0] sel);
    case (sel) 0: mux_970 = 1'h0; 1: mux_970 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_971;
  wire [0:0] v_972;
  wire [0:0] v_973;
  function [0:0] mux_973(input [0:0] sel);
    case (sel) 0: mux_973 = 1'h0; 1: mux_973 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_974;
  wire [0:0] v_975;
  wire [0:0] v_976;
  wire [0:0] vin0_consume_en_977;
  wire [0:0] vout_canPeek_977;
  wire [7:0] vout_peek_977;
  wire [0:0] v_978;
  function [0:0] mux_978(input [0:0] sel);
    case (sel) 0: mux_978 = 1'h0; 1: mux_978 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_979;
  wire [0:0] v_980;
  wire [0:0] v_981;
  function [0:0] mux_981(input [0:0] sel);
    case (sel) 0: mux_981 = 1'h0; 1: mux_981 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_982;
  wire [0:0] vin0_consume_en_983;
  wire [0:0] vout_canPeek_983;
  wire [7:0] vout_peek_983;
  wire [0:0] v_984;
  function [0:0] mux_984(input [0:0] sel);
    case (sel) 0: mux_984 = 1'h0; 1: mux_984 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_985;
  wire [0:0] v_986;
  wire [0:0] v_987;
  function [0:0] mux_987(input [0:0] sel);
    case (sel) 0: mux_987 = 1'h0; 1: mux_987 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_988;
  wire [0:0] v_989;
  wire [0:0] v_990;
  wire [0:0] vin0_consume_en_991;
  wire [0:0] vout_canPeek_991;
  wire [7:0] vout_peek_991;
  wire [0:0] v_992;
  function [0:0] mux_992(input [0:0] sel);
    case (sel) 0: mux_992 = 1'h0; 1: mux_992 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_993;
  wire [0:0] v_994;
  wire [0:0] v_995;
  function [0:0] mux_995(input [0:0] sel);
    case (sel) 0: mux_995 = 1'h0; 1: mux_995 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_996;
  wire [0:0] vin0_consume_en_997;
  wire [0:0] vout_canPeek_997;
  wire [7:0] vout_peek_997;
  wire [0:0] v_998;
  function [0:0] mux_998(input [0:0] sel);
    case (sel) 0: mux_998 = 1'h0; 1: mux_998 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_999;
  wire [0:0] v_1000;
  wire [0:0] v_1001;
  function [0:0] mux_1001(input [0:0] sel);
    case (sel) 0: mux_1001 = 1'h0; 1: mux_1001 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1002;
  wire [0:0] v_1003;
  wire [0:0] v_1004;
  wire [0:0] vin0_consume_en_1005;
  wire [0:0] vout_canPeek_1005;
  wire [7:0] vout_peek_1005;
  wire [0:0] v_1006;
  function [0:0] mux_1006(input [0:0] sel);
    case (sel) 0: mux_1006 = 1'h0; 1: mux_1006 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1007;
  wire [0:0] v_1008;
  wire [0:0] v_1009;
  function [0:0] mux_1009(input [0:0] sel);
    case (sel) 0: mux_1009 = 1'h0; 1: mux_1009 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1010;
  wire [0:0] vin0_consume_en_1011;
  wire [0:0] vout_canPeek_1011;
  wire [7:0] vout_peek_1011;
  wire [0:0] v_1012;
  function [0:0] mux_1012(input [0:0] sel);
    case (sel) 0: mux_1012 = 1'h0; 1: mux_1012 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1013;
  wire [0:0] v_1014;
  wire [0:0] v_1015;
  function [0:0] mux_1015(input [0:0] sel);
    case (sel) 0: mux_1015 = 1'h0; 1: mux_1015 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1016;
  wire [0:0] v_1017;
  wire [0:0] v_1018;
  wire [0:0] vin0_consume_en_1019;
  wire [0:0] vout_canPeek_1019;
  wire [7:0] vout_peek_1019;
  wire [0:0] v_1020;
  function [0:0] mux_1020(input [0:0] sel);
    case (sel) 0: mux_1020 = 1'h0; 1: mux_1020 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1021;
  wire [0:0] v_1022;
  wire [0:0] v_1023;
  function [0:0] mux_1023(input [0:0] sel);
    case (sel) 0: mux_1023 = 1'h0; 1: mux_1023 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1024;
  wire [0:0] vin0_consume_en_1025;
  wire [0:0] vout_canPeek_1025;
  wire [7:0] vout_peek_1025;
  wire [0:0] v_1026;
  function [0:0] mux_1026(input [0:0] sel);
    case (sel) 0: mux_1026 = 1'h0; 1: mux_1026 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1027;
  wire [0:0] v_1028;
  wire [0:0] v_1029;
  function [0:0] mux_1029(input [0:0] sel);
    case (sel) 0: mux_1029 = 1'h0; 1: mux_1029 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1030;
  wire [0:0] v_1031;
  wire [0:0] v_1032;
  wire [0:0] vin0_consume_en_1033;
  wire [0:0] vout_canPeek_1033;
  wire [7:0] vout_peek_1033;
  wire [0:0] v_1034;
  function [0:0] mux_1034(input [0:0] sel);
    case (sel) 0: mux_1034 = 1'h0; 1: mux_1034 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1035;
  wire [0:0] v_1036;
  wire [0:0] v_1037;
  function [0:0] mux_1037(input [0:0] sel);
    case (sel) 0: mux_1037 = 1'h0; 1: mux_1037 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1038;
  wire [0:0] vin0_consume_en_1039;
  wire [0:0] vout_canPeek_1039;
  wire [7:0] vout_peek_1039;
  wire [0:0] v_1040;
  function [0:0] mux_1040(input [0:0] sel);
    case (sel) 0: mux_1040 = 1'h0; 1: mux_1040 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1041;
  wire [0:0] v_1042;
  wire [0:0] v_1043;
  function [0:0] mux_1043(input [0:0] sel);
    case (sel) 0: mux_1043 = 1'h0; 1: mux_1043 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1044;
  wire [0:0] v_1045;
  wire [0:0] v_1046;
  wire [0:0] vin0_consume_en_1047;
  wire [0:0] vout_canPeek_1047;
  wire [7:0] vout_peek_1047;
  wire [0:0] v_1048;
  function [0:0] mux_1048(input [0:0] sel);
    case (sel) 0: mux_1048 = 1'h0; 1: mux_1048 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1049;
  wire [0:0] v_1050;
  wire [0:0] v_1051;
  function [0:0] mux_1051(input [0:0] sel);
    case (sel) 0: mux_1051 = 1'h0; 1: mux_1051 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1052;
  wire [0:0] vin0_consume_en_1053;
  wire [0:0] vout_canPeek_1053;
  wire [7:0] vout_peek_1053;
  wire [0:0] v_1054;
  function [0:0] mux_1054(input [0:0] sel);
    case (sel) 0: mux_1054 = 1'h0; 1: mux_1054 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1055;
  wire [0:0] v_1056;
  wire [0:0] v_1057;
  function [0:0] mux_1057(input [0:0] sel);
    case (sel) 0: mux_1057 = 1'h0; 1: mux_1057 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1058;
  wire [0:0] v_1059;
  wire [0:0] v_1060;
  wire [0:0] vin0_consume_en_1061;
  wire [0:0] vout_canPeek_1061;
  wire [7:0] vout_peek_1061;
  wire [0:0] v_1062;
  function [0:0] mux_1062(input [0:0] sel);
    case (sel) 0: mux_1062 = 1'h0; 1: mux_1062 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1063;
  wire [0:0] v_1064;
  wire [0:0] v_1065;
  function [0:0] mux_1065(input [0:0] sel);
    case (sel) 0: mux_1065 = 1'h0; 1: mux_1065 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1066;
  wire [0:0] vin0_consume_en_1067;
  wire [0:0] vout_canPeek_1067;
  wire [7:0] vout_peek_1067;
  wire [0:0] v_1068;
  function [0:0] mux_1068(input [0:0] sel);
    case (sel) 0: mux_1068 = 1'h0; 1: mux_1068 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1069;
  wire [0:0] v_1070;
  wire [0:0] v_1071;
  function [0:0] mux_1071(input [0:0] sel);
    case (sel) 0: mux_1071 = 1'h0; 1: mux_1071 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1072;
  wire [0:0] v_1073;
  wire [0:0] v_1074;
  wire [0:0] vin0_consume_en_1075;
  wire [0:0] vout_canPeek_1075;
  wire [7:0] vout_peek_1075;
  wire [0:0] v_1076;
  function [0:0] mux_1076(input [0:0] sel);
    case (sel) 0: mux_1076 = 1'h0; 1: mux_1076 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1077;
  wire [0:0] v_1078;
  wire [0:0] v_1079;
  function [0:0] mux_1079(input [0:0] sel);
    case (sel) 0: mux_1079 = 1'h0; 1: mux_1079 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1080;
  wire [0:0] vin0_consume_en_1081;
  wire [0:0] vout_canPeek_1081;
  wire [7:0] vout_peek_1081;
  wire [0:0] v_1082;
  function [0:0] mux_1082(input [0:0] sel);
    case (sel) 0: mux_1082 = 1'h0; 1: mux_1082 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1083;
  wire [0:0] v_1084;
  wire [0:0] v_1085;
  function [0:0] mux_1085(input [0:0] sel);
    case (sel) 0: mux_1085 = 1'h0; 1: mux_1085 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1086;
  wire [0:0] v_1087;
  wire [0:0] v_1088;
  wire [0:0] vin0_consume_en_1089;
  wire [0:0] vout_canPeek_1089;
  wire [7:0] vout_peek_1089;
  wire [0:0] v_1090;
  function [0:0] mux_1090(input [0:0] sel);
    case (sel) 0: mux_1090 = 1'h0; 1: mux_1090 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1091;
  wire [0:0] v_1092;
  wire [0:0] v_1093;
  function [0:0] mux_1093(input [0:0] sel);
    case (sel) 0: mux_1093 = 1'h0; 1: mux_1093 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1094;
  wire [0:0] vin0_consume_en_1095;
  wire [0:0] vout_canPeek_1095;
  wire [7:0] vout_peek_1095;
  wire [0:0] v_1096;
  function [0:0] mux_1096(input [0:0] sel);
    case (sel) 0: mux_1096 = 1'h0; 1: mux_1096 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1097;
  wire [0:0] v_1098;
  wire [0:0] v_1099;
  function [0:0] mux_1099(input [0:0] sel);
    case (sel) 0: mux_1099 = 1'h0; 1: mux_1099 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1100;
  wire [0:0] v_1101;
  wire [0:0] v_1102;
  wire [0:0] vin0_consume_en_1103;
  wire [0:0] vout_canPeek_1103;
  wire [7:0] vout_peek_1103;
  wire [0:0] v_1104;
  function [0:0] mux_1104(input [0:0] sel);
    case (sel) 0: mux_1104 = 1'h0; 1: mux_1104 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1105;
  wire [0:0] v_1106;
  wire [0:0] v_1107;
  function [0:0] mux_1107(input [0:0] sel);
    case (sel) 0: mux_1107 = 1'h0; 1: mux_1107 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1108;
  wire [0:0] vin0_consume_en_1109;
  wire [0:0] vout_canPeek_1109;
  wire [7:0] vout_peek_1109;
  wire [0:0] v_1110;
  function [0:0] mux_1110(input [0:0] sel);
    case (sel) 0: mux_1110 = 1'h0; 1: mux_1110 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1111;
  wire [0:0] v_1112;
  wire [0:0] v_1113;
  function [0:0] mux_1113(input [0:0] sel);
    case (sel) 0: mux_1113 = 1'h0; 1: mux_1113 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1114;
  wire [0:0] v_1115;
  wire [0:0] v_1116;
  wire [0:0] vin0_consume_en_1117;
  wire [0:0] vout_canPeek_1117;
  wire [7:0] vout_peek_1117;
  wire [0:0] v_1118;
  function [0:0] mux_1118(input [0:0] sel);
    case (sel) 0: mux_1118 = 1'h0; 1: mux_1118 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1119;
  wire [0:0] v_1120;
  wire [0:0] v_1121;
  function [0:0] mux_1121(input [0:0] sel);
    case (sel) 0: mux_1121 = 1'h0; 1: mux_1121 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1122;
  wire [0:0] vin0_consume_en_1123;
  wire [0:0] vout_canPeek_1123;
  wire [7:0] vout_peek_1123;
  wire [0:0] v_1124;
  function [0:0] mux_1124(input [0:0] sel);
    case (sel) 0: mux_1124 = 1'h0; 1: mux_1124 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1125;
  wire [0:0] v_1126;
  wire [0:0] v_1127;
  function [0:0] mux_1127(input [0:0] sel);
    case (sel) 0: mux_1127 = 1'h0; 1: mux_1127 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1128;
  wire [0:0] v_1129;
  wire [0:0] v_1130;
  wire [0:0] vin0_consume_en_1131;
  wire [0:0] vout_canPeek_1131;
  wire [7:0] vout_peek_1131;
  wire [0:0] v_1132;
  function [0:0] mux_1132(input [0:0] sel);
    case (sel) 0: mux_1132 = 1'h0; 1: mux_1132 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1133;
  wire [0:0] v_1134;
  wire [0:0] v_1135;
  function [0:0] mux_1135(input [0:0] sel);
    case (sel) 0: mux_1135 = 1'h0; 1: mux_1135 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1136;
  wire [0:0] vin0_consume_en_1137;
  wire [0:0] vout_canPeek_1137;
  wire [7:0] vout_peek_1137;
  wire [0:0] v_1138;
  function [0:0] mux_1138(input [0:0] sel);
    case (sel) 0: mux_1138 = 1'h0; 1: mux_1138 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1139;
  wire [0:0] v_1140;
  wire [0:0] v_1141;
  function [0:0] mux_1141(input [0:0] sel);
    case (sel) 0: mux_1141 = 1'h0; 1: mux_1141 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1142;
  wire [0:0] v_1143;
  wire [0:0] v_1144;
  wire [0:0] vin0_consume_en_1145;
  wire [0:0] vout_canPeek_1145;
  wire [7:0] vout_peek_1145;
  wire [0:0] v_1146;
  function [0:0] mux_1146(input [0:0] sel);
    case (sel) 0: mux_1146 = 1'h0; 1: mux_1146 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1147;
  wire [0:0] v_1148;
  wire [0:0] v_1149;
  function [0:0] mux_1149(input [0:0] sel);
    case (sel) 0: mux_1149 = 1'h0; 1: mux_1149 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1150;
  wire [0:0] vin0_consume_en_1151;
  wire [0:0] vout_canPeek_1151;
  wire [7:0] vout_peek_1151;
  wire [0:0] v_1152;
  function [0:0] mux_1152(input [0:0] sel);
    case (sel) 0: mux_1152 = 1'h0; 1: mux_1152 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1153;
  wire [0:0] v_1154;
  wire [0:0] v_1155;
  function [0:0] mux_1155(input [0:0] sel);
    case (sel) 0: mux_1155 = 1'h0; 1: mux_1155 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1156;
  wire [0:0] v_1157;
  wire [0:0] v_1158;
  wire [0:0] vin0_consume_en_1159;
  wire [0:0] vout_canPeek_1159;
  wire [7:0] vout_peek_1159;
  wire [0:0] v_1160;
  function [0:0] mux_1160(input [0:0] sel);
    case (sel) 0: mux_1160 = 1'h0; 1: mux_1160 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1161;
  wire [0:0] v_1162;
  wire [0:0] v_1163;
  function [0:0] mux_1163(input [0:0] sel);
    case (sel) 0: mux_1163 = 1'h0; 1: mux_1163 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1164;
  wire [0:0] vin0_consume_en_1165;
  wire [0:0] vout_canPeek_1165;
  wire [7:0] vout_peek_1165;
  wire [0:0] v_1166;
  function [0:0] mux_1166(input [0:0] sel);
    case (sel) 0: mux_1166 = 1'h0; 1: mux_1166 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1167;
  wire [0:0] v_1168;
  wire [0:0] v_1169;
  function [0:0] mux_1169(input [0:0] sel);
    case (sel) 0: mux_1169 = 1'h0; 1: mux_1169 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1170;
  wire [0:0] v_1171;
  wire [0:0] v_1172;
  wire [0:0] vin0_consume_en_1173;
  wire [0:0] vout_canPeek_1173;
  wire [7:0] vout_peek_1173;
  wire [0:0] v_1174;
  function [0:0] mux_1174(input [0:0] sel);
    case (sel) 0: mux_1174 = 1'h0; 1: mux_1174 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1175;
  wire [0:0] v_1176;
  wire [0:0] v_1177;
  function [0:0] mux_1177(input [0:0] sel);
    case (sel) 0: mux_1177 = 1'h0; 1: mux_1177 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1178;
  wire [0:0] vin0_consume_en_1179;
  wire [0:0] vout_canPeek_1179;
  wire [7:0] vout_peek_1179;
  wire [0:0] v_1180;
  function [0:0] mux_1180(input [0:0] sel);
    case (sel) 0: mux_1180 = 1'h0; 1: mux_1180 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1181;
  wire [0:0] v_1182;
  wire [0:0] v_1183;
  function [0:0] mux_1183(input [0:0] sel);
    case (sel) 0: mux_1183 = 1'h0; 1: mux_1183 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1184;
  wire [0:0] v_1185;
  wire [0:0] v_1186;
  wire [0:0] vin0_consume_en_1187;
  wire [0:0] vout_canPeek_1187;
  wire [7:0] vout_peek_1187;
  wire [0:0] v_1188;
  function [0:0] mux_1188(input [0:0] sel);
    case (sel) 0: mux_1188 = 1'h0; 1: mux_1188 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1189;
  wire [0:0] v_1190;
  wire [0:0] v_1191;
  function [0:0] mux_1191(input [0:0] sel);
    case (sel) 0: mux_1191 = 1'h0; 1: mux_1191 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1192;
  wire [0:0] vin0_consume_en_1193;
  wire [0:0] vout_canPeek_1193;
  wire [7:0] vout_peek_1193;
  wire [0:0] v_1194;
  function [0:0] mux_1194(input [0:0] sel);
    case (sel) 0: mux_1194 = 1'h0; 1: mux_1194 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1195;
  wire [0:0] v_1196;
  wire [0:0] v_1197;
  function [0:0] mux_1197(input [0:0] sel);
    case (sel) 0: mux_1197 = 1'h0; 1: mux_1197 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1198;
  wire [0:0] v_1199;
  wire [0:0] v_1200;
  wire [0:0] vin0_consume_en_1201;
  wire [0:0] vout_canPeek_1201;
  wire [7:0] vout_peek_1201;
  wire [0:0] v_1202;
  function [0:0] mux_1202(input [0:0] sel);
    case (sel) 0: mux_1202 = 1'h0; 1: mux_1202 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1203;
  wire [0:0] v_1204;
  wire [0:0] v_1205;
  function [0:0] mux_1205(input [0:0] sel);
    case (sel) 0: mux_1205 = 1'h0; 1: mux_1205 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1206;
  wire [0:0] vin0_consume_en_1207;
  wire [0:0] vout_canPeek_1207;
  wire [7:0] vout_peek_1207;
  wire [0:0] v_1208;
  function [0:0] mux_1208(input [0:0] sel);
    case (sel) 0: mux_1208 = 1'h0; 1: mux_1208 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1209;
  wire [0:0] v_1210;
  wire [0:0] v_1211;
  function [0:0] mux_1211(input [0:0] sel);
    case (sel) 0: mux_1211 = 1'h0; 1: mux_1211 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1212;
  wire [0:0] v_1213;
  wire [0:0] v_1214;
  wire [0:0] vin0_consume_en_1215;
  wire [0:0] vout_canPeek_1215;
  wire [7:0] vout_peek_1215;
  wire [0:0] v_1216;
  function [0:0] mux_1216(input [0:0] sel);
    case (sel) 0: mux_1216 = 1'h0; 1: mux_1216 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1217;
  wire [0:0] v_1218;
  wire [0:0] v_1219;
  function [0:0] mux_1219(input [0:0] sel);
    case (sel) 0: mux_1219 = 1'h0; 1: mux_1219 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1220;
  wire [0:0] vin0_consume_en_1221;
  wire [0:0] vout_canPeek_1221;
  wire [7:0] vout_peek_1221;
  wire [0:0] v_1222;
  function [0:0] mux_1222(input [0:0] sel);
    case (sel) 0: mux_1222 = 1'h0; 1: mux_1222 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1223;
  wire [0:0] v_1224;
  wire [0:0] v_1225;
  function [0:0] mux_1225(input [0:0] sel);
    case (sel) 0: mux_1225 = 1'h0; 1: mux_1225 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1226;
  wire [0:0] v_1227;
  wire [0:0] v_1228;
  wire [0:0] vin0_consume_en_1229;
  wire [0:0] vout_canPeek_1229;
  wire [7:0] vout_peek_1229;
  wire [0:0] v_1230;
  function [0:0] mux_1230(input [0:0] sel);
    case (sel) 0: mux_1230 = 1'h0; 1: mux_1230 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1231;
  wire [0:0] v_1232;
  wire [0:0] v_1233;
  function [0:0] mux_1233(input [0:0] sel);
    case (sel) 0: mux_1233 = 1'h0; 1: mux_1233 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1234;
  wire [0:0] vin0_consume_en_1235;
  wire [0:0] vout_canPeek_1235;
  wire [7:0] vout_peek_1235;
  wire [0:0] v_1236;
  function [0:0] mux_1236(input [0:0] sel);
    case (sel) 0: mux_1236 = 1'h0; 1: mux_1236 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1237;
  wire [0:0] v_1238;
  wire [0:0] v_1239;
  function [0:0] mux_1239(input [0:0] sel);
    case (sel) 0: mux_1239 = 1'h0; 1: mux_1239 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1240;
  wire [0:0] v_1241;
  wire [0:0] v_1242;
  wire [0:0] vin0_consume_en_1243;
  wire [0:0] vout_canPeek_1243;
  wire [7:0] vout_peek_1243;
  wire [0:0] v_1244;
  function [0:0] mux_1244(input [0:0] sel);
    case (sel) 0: mux_1244 = 1'h0; 1: mux_1244 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1245;
  wire [0:0] v_1246;
  wire [0:0] v_1247;
  function [0:0] mux_1247(input [0:0] sel);
    case (sel) 0: mux_1247 = 1'h0; 1: mux_1247 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1248;
  wire [0:0] vin0_consume_en_1249;
  wire [0:0] vout_canPeek_1249;
  wire [7:0] vout_peek_1249;
  wire [0:0] v_1250;
  function [0:0] mux_1250(input [0:0] sel);
    case (sel) 0: mux_1250 = 1'h0; 1: mux_1250 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1251;
  wire [0:0] v_1252;
  wire [0:0] v_1253;
  function [0:0] mux_1253(input [0:0] sel);
    case (sel) 0: mux_1253 = 1'h0; 1: mux_1253 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1254;
  wire [0:0] v_1255;
  wire [0:0] v_1256;
  wire [0:0] vin0_consume_en_1257;
  wire [0:0] vout_canPeek_1257;
  wire [7:0] vout_peek_1257;
  wire [0:0] v_1258;
  function [0:0] mux_1258(input [0:0] sel);
    case (sel) 0: mux_1258 = 1'h0; 1: mux_1258 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1259;
  wire [0:0] v_1260;
  wire [0:0] v_1261;
  function [0:0] mux_1261(input [0:0] sel);
    case (sel) 0: mux_1261 = 1'h0; 1: mux_1261 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1262;
  wire [0:0] vin0_consume_en_1263;
  wire [0:0] vout_canPeek_1263;
  wire [7:0] vout_peek_1263;
  wire [0:0] v_1264;
  function [0:0] mux_1264(input [0:0] sel);
    case (sel) 0: mux_1264 = 1'h0; 1: mux_1264 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1265;
  wire [0:0] v_1266;
  wire [0:0] v_1267;
  function [0:0] mux_1267(input [0:0] sel);
    case (sel) 0: mux_1267 = 1'h0; 1: mux_1267 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1268;
  wire [0:0] v_1269;
  wire [0:0] v_1270;
  wire [0:0] vin0_consume_en_1271;
  wire [0:0] vout_canPeek_1271;
  wire [7:0] vout_peek_1271;
  wire [0:0] v_1272;
  function [0:0] mux_1272(input [0:0] sel);
    case (sel) 0: mux_1272 = 1'h0; 1: mux_1272 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1273;
  wire [0:0] v_1274;
  wire [0:0] v_1275;
  function [0:0] mux_1275(input [0:0] sel);
    case (sel) 0: mux_1275 = 1'h0; 1: mux_1275 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1276;
  wire [0:0] vin0_consume_en_1277;
  wire [0:0] vout_canPeek_1277;
  wire [7:0] vout_peek_1277;
  wire [0:0] v_1278;
  function [0:0] mux_1278(input [0:0] sel);
    case (sel) 0: mux_1278 = 1'h0; 1: mux_1278 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1279;
  wire [0:0] v_1280;
  wire [0:0] v_1281;
  function [0:0] mux_1281(input [0:0] sel);
    case (sel) 0: mux_1281 = 1'h0; 1: mux_1281 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1282;
  wire [0:0] v_1283;
  wire [0:0] v_1284;
  wire [0:0] vin0_consume_en_1285;
  wire [0:0] vout_canPeek_1285;
  wire [7:0] vout_peek_1285;
  wire [0:0] v_1286;
  function [0:0] mux_1286(input [0:0] sel);
    case (sel) 0: mux_1286 = 1'h0; 1: mux_1286 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1287;
  wire [0:0] v_1288;
  wire [0:0] v_1289;
  function [0:0] mux_1289(input [0:0] sel);
    case (sel) 0: mux_1289 = 1'h0; 1: mux_1289 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1290;
  wire [0:0] vin0_consume_en_1291;
  wire [0:0] vout_canPeek_1291;
  wire [7:0] vout_peek_1291;
  wire [0:0] v_1292;
  function [0:0] mux_1292(input [0:0] sel);
    case (sel) 0: mux_1292 = 1'h0; 1: mux_1292 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1293;
  wire [0:0] v_1294;
  wire [0:0] v_1295;
  function [0:0] mux_1295(input [0:0] sel);
    case (sel) 0: mux_1295 = 1'h0; 1: mux_1295 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1296;
  wire [0:0] v_1297;
  wire [0:0] v_1298;
  wire [0:0] vin0_consume_en_1299;
  wire [0:0] vout_canPeek_1299;
  wire [7:0] vout_peek_1299;
  wire [0:0] v_1300;
  function [0:0] mux_1300(input [0:0] sel);
    case (sel) 0: mux_1300 = 1'h0; 1: mux_1300 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1301;
  wire [0:0] v_1302;
  wire [0:0] v_1303;
  function [0:0] mux_1303(input [0:0] sel);
    case (sel) 0: mux_1303 = 1'h0; 1: mux_1303 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1304;
  wire [0:0] vin0_consume_en_1305;
  wire [0:0] vout_canPeek_1305;
  wire [7:0] vout_peek_1305;
  wire [0:0] v_1306;
  function [0:0] mux_1306(input [0:0] sel);
    case (sel) 0: mux_1306 = 1'h0; 1: mux_1306 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1307;
  wire [0:0] v_1308;
  wire [0:0] v_1309;
  function [0:0] mux_1309(input [0:0] sel);
    case (sel) 0: mux_1309 = 1'h0; 1: mux_1309 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1310;
  wire [0:0] v_1311;
  wire [0:0] v_1312;
  wire [0:0] vin0_consume_en_1313;
  wire [0:0] vout_canPeek_1313;
  wire [7:0] vout_peek_1313;
  wire [0:0] v_1314;
  function [0:0] mux_1314(input [0:0] sel);
    case (sel) 0: mux_1314 = 1'h0; 1: mux_1314 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1315;
  wire [0:0] v_1316;
  wire [0:0] v_1317;
  function [0:0] mux_1317(input [0:0] sel);
    case (sel) 0: mux_1317 = 1'h0; 1: mux_1317 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1318;
  wire [0:0] vin0_consume_en_1319;
  wire [0:0] vout_canPeek_1319;
  wire [7:0] vout_peek_1319;
  wire [0:0] v_1320;
  function [0:0] mux_1320(input [0:0] sel);
    case (sel) 0: mux_1320 = 1'h0; 1: mux_1320 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1321;
  wire [0:0] v_1322;
  wire [0:0] v_1323;
  function [0:0] mux_1323(input [0:0] sel);
    case (sel) 0: mux_1323 = 1'h0; 1: mux_1323 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1324;
  wire [0:0] v_1325;
  wire [0:0] v_1326;
  wire [0:0] vin0_consume_en_1327;
  wire [0:0] vout_canPeek_1327;
  wire [7:0] vout_peek_1327;
  wire [0:0] v_1328;
  function [0:0] mux_1328(input [0:0] sel);
    case (sel) 0: mux_1328 = 1'h0; 1: mux_1328 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1329;
  wire [0:0] v_1330;
  wire [0:0] v_1331;
  function [0:0] mux_1331(input [0:0] sel);
    case (sel) 0: mux_1331 = 1'h0; 1: mux_1331 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1332;
  wire [0:0] vin0_consume_en_1333;
  wire [0:0] vout_canPeek_1333;
  wire [7:0] vout_peek_1333;
  wire [0:0] v_1334;
  function [0:0] mux_1334(input [0:0] sel);
    case (sel) 0: mux_1334 = 1'h0; 1: mux_1334 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1335;
  wire [0:0] v_1336;
  wire [0:0] v_1337;
  function [0:0] mux_1337(input [0:0] sel);
    case (sel) 0: mux_1337 = 1'h0; 1: mux_1337 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1338;
  wire [0:0] v_1339;
  wire [0:0] v_1340;
  wire [0:0] vin0_consume_en_1341;
  wire [0:0] vout_canPeek_1341;
  wire [7:0] vout_peek_1341;
  wire [0:0] v_1342;
  function [0:0] mux_1342(input [0:0] sel);
    case (sel) 0: mux_1342 = 1'h0; 1: mux_1342 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1343;
  wire [0:0] v_1344;
  wire [0:0] v_1345;
  function [0:0] mux_1345(input [0:0] sel);
    case (sel) 0: mux_1345 = 1'h0; 1: mux_1345 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1346;
  wire [0:0] vin0_consume_en_1347;
  wire [0:0] vout_canPeek_1347;
  wire [7:0] vout_peek_1347;
  wire [0:0] v_1348;
  function [0:0] mux_1348(input [0:0] sel);
    case (sel) 0: mux_1348 = 1'h0; 1: mux_1348 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1349;
  wire [0:0] v_1350;
  wire [0:0] v_1351;
  function [0:0] mux_1351(input [0:0] sel);
    case (sel) 0: mux_1351 = 1'h0; 1: mux_1351 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1352;
  wire [0:0] v_1353;
  wire [0:0] v_1354;
  wire [0:0] vin0_consume_en_1355;
  wire [0:0] vout_canPeek_1355;
  wire [7:0] vout_peek_1355;
  wire [0:0] v_1356;
  function [0:0] mux_1356(input [0:0] sel);
    case (sel) 0: mux_1356 = 1'h0; 1: mux_1356 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1357;
  wire [0:0] v_1358;
  wire [0:0] v_1359;
  function [0:0] mux_1359(input [0:0] sel);
    case (sel) 0: mux_1359 = 1'h0; 1: mux_1359 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1360;
  wire [0:0] vin0_consume_en_1361;
  wire [0:0] vout_canPeek_1361;
  wire [7:0] vout_peek_1361;
  wire [0:0] v_1362;
  function [0:0] mux_1362(input [0:0] sel);
    case (sel) 0: mux_1362 = 1'h0; 1: mux_1362 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1363;
  wire [0:0] v_1364;
  wire [0:0] v_1365;
  function [0:0] mux_1365(input [0:0] sel);
    case (sel) 0: mux_1365 = 1'h0; 1: mux_1365 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1366;
  wire [0:0] v_1367;
  wire [0:0] v_1368;
  wire [0:0] vin0_consume_en_1369;
  wire [0:0] vout_canPeek_1369;
  wire [7:0] vout_peek_1369;
  wire [0:0] v_1370;
  function [0:0] mux_1370(input [0:0] sel);
    case (sel) 0: mux_1370 = 1'h0; 1: mux_1370 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1371;
  wire [0:0] v_1372;
  wire [0:0] v_1373;
  function [0:0] mux_1373(input [0:0] sel);
    case (sel) 0: mux_1373 = 1'h0; 1: mux_1373 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1374;
  wire [0:0] vin0_consume_en_1375;
  wire [0:0] vout_canPeek_1375;
  wire [7:0] vout_peek_1375;
  wire [0:0] v_1376;
  function [0:0] mux_1376(input [0:0] sel);
    case (sel) 0: mux_1376 = 1'h0; 1: mux_1376 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1377;
  wire [0:0] v_1378;
  wire [0:0] v_1379;
  function [0:0] mux_1379(input [0:0] sel);
    case (sel) 0: mux_1379 = 1'h0; 1: mux_1379 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1380;
  wire [0:0] v_1381;
  wire [0:0] v_1382;
  wire [0:0] vin0_consume_en_1383;
  wire [0:0] vout_canPeek_1383;
  wire [7:0] vout_peek_1383;
  wire [0:0] v_1384;
  function [0:0] mux_1384(input [0:0] sel);
    case (sel) 0: mux_1384 = 1'h0; 1: mux_1384 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1385;
  wire [0:0] v_1386;
  wire [0:0] v_1387;
  function [0:0] mux_1387(input [0:0] sel);
    case (sel) 0: mux_1387 = 1'h0; 1: mux_1387 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1388;
  wire [0:0] vin0_consume_en_1389;
  wire [0:0] vout_canPeek_1389;
  wire [7:0] vout_peek_1389;
  wire [0:0] v_1390;
  function [0:0] mux_1390(input [0:0] sel);
    case (sel) 0: mux_1390 = 1'h0; 1: mux_1390 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1391;
  wire [0:0] v_1392;
  wire [0:0] v_1393;
  function [0:0] mux_1393(input [0:0] sel);
    case (sel) 0: mux_1393 = 1'h0; 1: mux_1393 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1394;
  wire [0:0] v_1395;
  wire [0:0] v_1396;
  wire [0:0] vin0_consume_en_1397;
  wire [0:0] vout_canPeek_1397;
  wire [7:0] vout_peek_1397;
  wire [0:0] v_1398;
  function [0:0] mux_1398(input [0:0] sel);
    case (sel) 0: mux_1398 = 1'h0; 1: mux_1398 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1399;
  wire [0:0] v_1400;
  wire [0:0] v_1401;
  function [0:0] mux_1401(input [0:0] sel);
    case (sel) 0: mux_1401 = 1'h0; 1: mux_1401 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1402;
  wire [0:0] vin0_consume_en_1403;
  wire [0:0] vout_canPeek_1403;
  wire [7:0] vout_peek_1403;
  wire [0:0] v_1404;
  function [0:0] mux_1404(input [0:0] sel);
    case (sel) 0: mux_1404 = 1'h0; 1: mux_1404 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1405;
  wire [0:0] v_1406;
  wire [0:0] v_1407;
  function [0:0] mux_1407(input [0:0] sel);
    case (sel) 0: mux_1407 = 1'h0; 1: mux_1407 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1408;
  wire [0:0] v_1409;
  wire [0:0] v_1410;
  wire [0:0] vin0_consume_en_1411;
  wire [0:0] vout_canPeek_1411;
  wire [7:0] vout_peek_1411;
  wire [0:0] v_1412;
  function [0:0] mux_1412(input [0:0] sel);
    case (sel) 0: mux_1412 = 1'h0; 1: mux_1412 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1413;
  wire [0:0] v_1414;
  wire [0:0] v_1415;
  function [0:0] mux_1415(input [0:0] sel);
    case (sel) 0: mux_1415 = 1'h0; 1: mux_1415 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1416;
  wire [0:0] vin0_consume_en_1417;
  wire [0:0] vout_canPeek_1417;
  wire [7:0] vout_peek_1417;
  wire [0:0] v_1418;
  function [0:0] mux_1418(input [0:0] sel);
    case (sel) 0: mux_1418 = 1'h0; 1: mux_1418 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1419;
  wire [0:0] v_1420;
  wire [0:0] v_1421;
  function [0:0] mux_1421(input [0:0] sel);
    case (sel) 0: mux_1421 = 1'h0; 1: mux_1421 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1422;
  wire [0:0] v_1423;
  wire [0:0] v_1424;
  wire [0:0] vin0_consume_en_1425;
  wire [0:0] vout_canPeek_1425;
  wire [7:0] vout_peek_1425;
  wire [0:0] v_1426;
  function [0:0] mux_1426(input [0:0] sel);
    case (sel) 0: mux_1426 = 1'h0; 1: mux_1426 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1427;
  wire [0:0] v_1428;
  wire [0:0] v_1429;
  function [0:0] mux_1429(input [0:0] sel);
    case (sel) 0: mux_1429 = 1'h0; 1: mux_1429 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1430;
  wire [0:0] vin0_consume_en_1431;
  wire [0:0] vout_canPeek_1431;
  wire [7:0] vout_peek_1431;
  wire [0:0] v_1432;
  function [0:0] mux_1432(input [0:0] sel);
    case (sel) 0: mux_1432 = 1'h0; 1: mux_1432 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1433;
  wire [0:0] v_1434;
  wire [0:0] v_1435;
  function [0:0] mux_1435(input [0:0] sel);
    case (sel) 0: mux_1435 = 1'h0; 1: mux_1435 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1436;
  wire [0:0] v_1437;
  wire [0:0] v_1438;
  wire [0:0] vin0_consume_en_1439;
  wire [0:0] vout_canPeek_1439;
  wire [7:0] vout_peek_1439;
  wire [0:0] v_1440;
  function [0:0] mux_1440(input [0:0] sel);
    case (sel) 0: mux_1440 = 1'h0; 1: mux_1440 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1441;
  wire [0:0] v_1442;
  wire [0:0] v_1443;
  function [0:0] mux_1443(input [0:0] sel);
    case (sel) 0: mux_1443 = 1'h0; 1: mux_1443 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1444;
  wire [0:0] vin0_consume_en_1445;
  wire [0:0] vout_canPeek_1445;
  wire [7:0] vout_peek_1445;
  wire [0:0] v_1446;
  function [0:0] mux_1446(input [0:0] sel);
    case (sel) 0: mux_1446 = 1'h0; 1: mux_1446 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1447;
  wire [0:0] v_1448;
  wire [0:0] v_1449;
  function [0:0] mux_1449(input [0:0] sel);
    case (sel) 0: mux_1449 = 1'h0; 1: mux_1449 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1450;
  wire [0:0] v_1451;
  wire [0:0] v_1452;
  wire [0:0] vin0_consume_en_1453;
  wire [0:0] vout_canPeek_1453;
  wire [7:0] vout_peek_1453;
  wire [0:0] v_1454;
  function [0:0] mux_1454(input [0:0] sel);
    case (sel) 0: mux_1454 = 1'h0; 1: mux_1454 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1455;
  wire [0:0] v_1456;
  wire [0:0] v_1457;
  function [0:0] mux_1457(input [0:0] sel);
    case (sel) 0: mux_1457 = 1'h0; 1: mux_1457 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1458;
  wire [0:0] vin0_consume_en_1459;
  wire [0:0] vout_canPeek_1459;
  wire [7:0] vout_peek_1459;
  wire [0:0] v_1460;
  function [0:0] mux_1460(input [0:0] sel);
    case (sel) 0: mux_1460 = 1'h0; 1: mux_1460 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1461;
  wire [0:0] v_1462;
  wire [0:0] v_1463;
  function [0:0] mux_1463(input [0:0] sel);
    case (sel) 0: mux_1463 = 1'h0; 1: mux_1463 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1464;
  wire [0:0] v_1465;
  wire [0:0] v_1466;
  wire [0:0] vin0_consume_en_1467;
  wire [0:0] vout_canPeek_1467;
  wire [7:0] vout_peek_1467;
  wire [0:0] v_1468;
  function [0:0] mux_1468(input [0:0] sel);
    case (sel) 0: mux_1468 = 1'h0; 1: mux_1468 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1469;
  wire [0:0] v_1470;
  wire [0:0] v_1471;
  function [0:0] mux_1471(input [0:0] sel);
    case (sel) 0: mux_1471 = 1'h0; 1: mux_1471 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1472;
  wire [0:0] vin0_consume_en_1473;
  wire [0:0] vout_canPeek_1473;
  wire [7:0] vout_peek_1473;
  wire [0:0] v_1474;
  function [0:0] mux_1474(input [0:0] sel);
    case (sel) 0: mux_1474 = 1'h0; 1: mux_1474 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1475;
  wire [0:0] v_1476;
  wire [0:0] v_1477;
  function [0:0] mux_1477(input [0:0] sel);
    case (sel) 0: mux_1477 = 1'h0; 1: mux_1477 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1478;
  wire [0:0] v_1479;
  wire [0:0] v_1480;
  wire [0:0] vin0_consume_en_1481;
  wire [0:0] vout_canPeek_1481;
  wire [7:0] vout_peek_1481;
  wire [0:0] v_1482;
  function [0:0] mux_1482(input [0:0] sel);
    case (sel) 0: mux_1482 = 1'h0; 1: mux_1482 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1483;
  wire [0:0] v_1484;
  wire [0:0] v_1485;
  function [0:0] mux_1485(input [0:0] sel);
    case (sel) 0: mux_1485 = 1'h0; 1: mux_1485 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1486;
  wire [0:0] vin0_consume_en_1487;
  wire [0:0] vout_canPeek_1487;
  wire [7:0] vout_peek_1487;
  wire [0:0] v_1488;
  function [0:0] mux_1488(input [0:0] sel);
    case (sel) 0: mux_1488 = 1'h0; 1: mux_1488 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1489;
  wire [0:0] v_1490;
  wire [0:0] v_1491;
  function [0:0] mux_1491(input [0:0] sel);
    case (sel) 0: mux_1491 = 1'h0; 1: mux_1491 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1492;
  wire [0:0] v_1493;
  wire [0:0] v_1494;
  wire [0:0] vin0_consume_en_1495;
  wire [0:0] vout_canPeek_1495;
  wire [7:0] vout_peek_1495;
  wire [0:0] v_1496;
  function [0:0] mux_1496(input [0:0] sel);
    case (sel) 0: mux_1496 = 1'h0; 1: mux_1496 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1497;
  wire [0:0] v_1498;
  wire [0:0] v_1499;
  function [0:0] mux_1499(input [0:0] sel);
    case (sel) 0: mux_1499 = 1'h0; 1: mux_1499 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1500;
  wire [0:0] vin0_consume_en_1501;
  wire [0:0] vout_canPeek_1501;
  wire [7:0] vout_peek_1501;
  wire [0:0] v_1502;
  function [0:0] mux_1502(input [0:0] sel);
    case (sel) 0: mux_1502 = 1'h0; 1: mux_1502 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1503;
  wire [0:0] v_1504;
  wire [0:0] v_1505;
  function [0:0] mux_1505(input [0:0] sel);
    case (sel) 0: mux_1505 = 1'h0; 1: mux_1505 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1506;
  wire [0:0] v_1507;
  wire [0:0] v_1508;
  wire [0:0] vin0_consume_en_1509;
  wire [0:0] vout_canPeek_1509;
  wire [7:0] vout_peek_1509;
  wire [0:0] v_1510;
  function [0:0] mux_1510(input [0:0] sel);
    case (sel) 0: mux_1510 = 1'h0; 1: mux_1510 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1511;
  wire [0:0] v_1512;
  wire [0:0] v_1513;
  function [0:0] mux_1513(input [0:0] sel);
    case (sel) 0: mux_1513 = 1'h0; 1: mux_1513 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1514;
  wire [0:0] vin0_consume_en_1515;
  wire [0:0] vout_canPeek_1515;
  wire [7:0] vout_peek_1515;
  wire [0:0] v_1516;
  function [0:0] mux_1516(input [0:0] sel);
    case (sel) 0: mux_1516 = 1'h0; 1: mux_1516 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1517;
  wire [0:0] v_1518;
  wire [0:0] v_1519;
  function [0:0] mux_1519(input [0:0] sel);
    case (sel) 0: mux_1519 = 1'h0; 1: mux_1519 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1520;
  wire [0:0] v_1521;
  wire [0:0] v_1522;
  wire [0:0] vin0_consume_en_1523;
  wire [0:0] vout_canPeek_1523;
  wire [7:0] vout_peek_1523;
  wire [0:0] v_1524;
  function [0:0] mux_1524(input [0:0] sel);
    case (sel) 0: mux_1524 = 1'h0; 1: mux_1524 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1525;
  wire [0:0] v_1526;
  wire [0:0] v_1527;
  function [0:0] mux_1527(input [0:0] sel);
    case (sel) 0: mux_1527 = 1'h0; 1: mux_1527 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1528;
  wire [0:0] vin0_consume_en_1529;
  wire [0:0] vout_canPeek_1529;
  wire [7:0] vout_peek_1529;
  wire [0:0] v_1530;
  function [0:0] mux_1530(input [0:0] sel);
    case (sel) 0: mux_1530 = 1'h0; 1: mux_1530 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1531;
  wire [0:0] v_1532;
  wire [0:0] v_1533;
  function [0:0] mux_1533(input [0:0] sel);
    case (sel) 0: mux_1533 = 1'h0; 1: mux_1533 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1534;
  wire [0:0] v_1535;
  wire [0:0] v_1536;
  wire [0:0] vin0_consume_en_1537;
  wire [0:0] vout_canPeek_1537;
  wire [7:0] vout_peek_1537;
  wire [0:0] v_1538;
  function [0:0] mux_1538(input [0:0] sel);
    case (sel) 0: mux_1538 = 1'h0; 1: mux_1538 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1539;
  wire [0:0] v_1540;
  wire [0:0] v_1541;
  function [0:0] mux_1541(input [0:0] sel);
    case (sel) 0: mux_1541 = 1'h0; 1: mux_1541 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1542;
  wire [0:0] vin0_consume_en_1543;
  wire [0:0] vout_canPeek_1543;
  wire [7:0] vout_peek_1543;
  wire [0:0] v_1544;
  function [0:0] mux_1544(input [0:0] sel);
    case (sel) 0: mux_1544 = 1'h0; 1: mux_1544 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1545;
  wire [0:0] v_1546;
  wire [0:0] v_1547;
  function [0:0] mux_1547(input [0:0] sel);
    case (sel) 0: mux_1547 = 1'h0; 1: mux_1547 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1548;
  wire [0:0] v_1549;
  wire [0:0] v_1550;
  wire [0:0] vin0_consume_en_1551;
  wire [0:0] vout_canPeek_1551;
  wire [7:0] vout_peek_1551;
  wire [0:0] v_1552;
  function [0:0] mux_1552(input [0:0] sel);
    case (sel) 0: mux_1552 = 1'h0; 1: mux_1552 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1553;
  wire [0:0] v_1554;
  wire [0:0] v_1555;
  function [0:0] mux_1555(input [0:0] sel);
    case (sel) 0: mux_1555 = 1'h0; 1: mux_1555 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1556;
  wire [0:0] vin0_consume_en_1557;
  wire [0:0] vout_canPeek_1557;
  wire [7:0] vout_peek_1557;
  wire [0:0] v_1558;
  function [0:0] mux_1558(input [0:0] sel);
    case (sel) 0: mux_1558 = 1'h0; 1: mux_1558 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1559;
  wire [0:0] v_1560;
  wire [0:0] v_1561;
  function [0:0] mux_1561(input [0:0] sel);
    case (sel) 0: mux_1561 = 1'h0; 1: mux_1561 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1562;
  wire [0:0] v_1563;
  wire [0:0] v_1564;
  wire [0:0] vin0_consume_en_1565;
  wire [0:0] vout_canPeek_1565;
  wire [7:0] vout_peek_1565;
  wire [0:0] v_1566;
  function [0:0] mux_1566(input [0:0] sel);
    case (sel) 0: mux_1566 = 1'h0; 1: mux_1566 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1567;
  wire [0:0] v_1568;
  wire [0:0] v_1569;
  function [0:0] mux_1569(input [0:0] sel);
    case (sel) 0: mux_1569 = 1'h0; 1: mux_1569 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1570;
  wire [0:0] vin0_consume_en_1571;
  wire [0:0] vout_canPeek_1571;
  wire [7:0] vout_peek_1571;
  wire [0:0] v_1572;
  function [0:0] mux_1572(input [0:0] sel);
    case (sel) 0: mux_1572 = 1'h0; 1: mux_1572 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1573;
  wire [0:0] v_1574;
  wire [0:0] v_1575;
  function [0:0] mux_1575(input [0:0] sel);
    case (sel) 0: mux_1575 = 1'h0; 1: mux_1575 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1576;
  wire [0:0] v_1577;
  wire [0:0] v_1578;
  wire [0:0] vin0_consume_en_1579;
  wire [0:0] vout_canPeek_1579;
  wire [7:0] vout_peek_1579;
  wire [0:0] v_1580;
  function [0:0] mux_1580(input [0:0] sel);
    case (sel) 0: mux_1580 = 1'h0; 1: mux_1580 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1581;
  wire [0:0] v_1582;
  wire [0:0] v_1583;
  function [0:0] mux_1583(input [0:0] sel);
    case (sel) 0: mux_1583 = 1'h0; 1: mux_1583 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1584;
  wire [0:0] vin0_consume_en_1585;
  wire [0:0] vout_canPeek_1585;
  wire [7:0] vout_peek_1585;
  wire [0:0] v_1586;
  function [0:0] mux_1586(input [0:0] sel);
    case (sel) 0: mux_1586 = 1'h0; 1: mux_1586 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1587;
  wire [0:0] v_1588;
  wire [0:0] v_1589;
  function [0:0] mux_1589(input [0:0] sel);
    case (sel) 0: mux_1589 = 1'h0; 1: mux_1589 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1590;
  wire [0:0] v_1591;
  wire [0:0] v_1592;
  wire [0:0] vin0_consume_en_1593;
  wire [0:0] vout_canPeek_1593;
  wire [7:0] vout_peek_1593;
  wire [0:0] v_1594;
  function [0:0] mux_1594(input [0:0] sel);
    case (sel) 0: mux_1594 = 1'h0; 1: mux_1594 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1595;
  wire [0:0] v_1596;
  wire [0:0] v_1597;
  function [0:0] mux_1597(input [0:0] sel);
    case (sel) 0: mux_1597 = 1'h0; 1: mux_1597 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1598;
  wire [0:0] vin0_consume_en_1599;
  wire [0:0] vout_canPeek_1599;
  wire [7:0] vout_peek_1599;
  wire [0:0] v_1600;
  function [0:0] mux_1600(input [0:0] sel);
    case (sel) 0: mux_1600 = 1'h0; 1: mux_1600 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1601;
  wire [0:0] v_1602;
  wire [0:0] v_1603;
  function [0:0] mux_1603(input [0:0] sel);
    case (sel) 0: mux_1603 = 1'h0; 1: mux_1603 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1604;
  wire [0:0] v_1605;
  wire [0:0] v_1606;
  wire [0:0] vin0_consume_en_1607;
  wire [0:0] vout_canPeek_1607;
  wire [7:0] vout_peek_1607;
  wire [0:0] v_1608;
  function [0:0] mux_1608(input [0:0] sel);
    case (sel) 0: mux_1608 = 1'h0; 1: mux_1608 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1609;
  wire [0:0] v_1610;
  wire [0:0] v_1611;
  function [0:0] mux_1611(input [0:0] sel);
    case (sel) 0: mux_1611 = 1'h0; 1: mux_1611 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1612;
  wire [0:0] vin0_consume_en_1613;
  wire [0:0] vout_canPeek_1613;
  wire [7:0] vout_peek_1613;
  wire [0:0] v_1614;
  function [0:0] mux_1614(input [0:0] sel);
    case (sel) 0: mux_1614 = 1'h0; 1: mux_1614 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1615;
  wire [0:0] v_1616;
  wire [0:0] v_1617;
  function [0:0] mux_1617(input [0:0] sel);
    case (sel) 0: mux_1617 = 1'h0; 1: mux_1617 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1618;
  wire [0:0] v_1619;
  wire [0:0] v_1620;
  wire [0:0] vin0_consume_en_1621;
  wire [0:0] vout_canPeek_1621;
  wire [7:0] vout_peek_1621;
  wire [0:0] v_1622;
  function [0:0] mux_1622(input [0:0] sel);
    case (sel) 0: mux_1622 = 1'h0; 1: mux_1622 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1623;
  wire [0:0] v_1624;
  wire [0:0] v_1625;
  function [0:0] mux_1625(input [0:0] sel);
    case (sel) 0: mux_1625 = 1'h0; 1: mux_1625 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1626;
  wire [0:0] vin0_consume_en_1627;
  wire [0:0] vout_canPeek_1627;
  wire [7:0] vout_peek_1627;
  wire [0:0] v_1628;
  function [0:0] mux_1628(input [0:0] sel);
    case (sel) 0: mux_1628 = 1'h0; 1: mux_1628 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1629;
  wire [0:0] v_1630;
  wire [0:0] v_1631;
  function [0:0] mux_1631(input [0:0] sel);
    case (sel) 0: mux_1631 = 1'h0; 1: mux_1631 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1632;
  wire [0:0] v_1633;
  wire [0:0] v_1634;
  wire [0:0] vin0_consume_en_1635;
  wire [0:0] vout_canPeek_1635;
  wire [7:0] vout_peek_1635;
  wire [0:0] v_1636;
  function [0:0] mux_1636(input [0:0] sel);
    case (sel) 0: mux_1636 = 1'h0; 1: mux_1636 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1637;
  wire [0:0] v_1638;
  wire [0:0] v_1639;
  function [0:0] mux_1639(input [0:0] sel);
    case (sel) 0: mux_1639 = 1'h0; 1: mux_1639 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1640;
  wire [0:0] vin0_consume_en_1641;
  wire [0:0] vout_canPeek_1641;
  wire [7:0] vout_peek_1641;
  wire [0:0] v_1642;
  function [0:0] mux_1642(input [0:0] sel);
    case (sel) 0: mux_1642 = 1'h0; 1: mux_1642 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1643;
  wire [0:0] v_1644;
  wire [0:0] v_1645;
  function [0:0] mux_1645(input [0:0] sel);
    case (sel) 0: mux_1645 = 1'h0; 1: mux_1645 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1646;
  wire [0:0] v_1647;
  wire [0:0] v_1648;
  wire [0:0] vin0_consume_en_1649;
  wire [0:0] vout_canPeek_1649;
  wire [7:0] vout_peek_1649;
  wire [0:0] v_1650;
  function [0:0] mux_1650(input [0:0] sel);
    case (sel) 0: mux_1650 = 1'h0; 1: mux_1650 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1651;
  wire [0:0] v_1652;
  wire [0:0] v_1653;
  function [0:0] mux_1653(input [0:0] sel);
    case (sel) 0: mux_1653 = 1'h0; 1: mux_1653 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1654;
  wire [0:0] vin0_consume_en_1655;
  wire [0:0] vout_canPeek_1655;
  wire [7:0] vout_peek_1655;
  wire [0:0] v_1656;
  function [0:0] mux_1656(input [0:0] sel);
    case (sel) 0: mux_1656 = 1'h0; 1: mux_1656 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1657;
  wire [0:0] v_1658;
  wire [0:0] v_1659;
  function [0:0] mux_1659(input [0:0] sel);
    case (sel) 0: mux_1659 = 1'h0; 1: mux_1659 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1660;
  wire [0:0] v_1661;
  wire [0:0] v_1662;
  wire [0:0] vin0_consume_en_1663;
  wire [0:0] vout_canPeek_1663;
  wire [7:0] vout_peek_1663;
  wire [0:0] v_1664;
  function [0:0] mux_1664(input [0:0] sel);
    case (sel) 0: mux_1664 = 1'h0; 1: mux_1664 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1665;
  wire [0:0] v_1666;
  wire [0:0] v_1667;
  function [0:0] mux_1667(input [0:0] sel);
    case (sel) 0: mux_1667 = 1'h0; 1: mux_1667 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1668;
  wire [0:0] vin0_consume_en_1669;
  wire [0:0] vout_canPeek_1669;
  wire [7:0] vout_peek_1669;
  wire [0:0] v_1670;
  function [0:0] mux_1670(input [0:0] sel);
    case (sel) 0: mux_1670 = 1'h0; 1: mux_1670 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1671;
  wire [0:0] v_1672;
  wire [0:0] v_1673;
  function [0:0] mux_1673(input [0:0] sel);
    case (sel) 0: mux_1673 = 1'h0; 1: mux_1673 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1674;
  wire [0:0] v_1675;
  wire [0:0] v_1676;
  wire [0:0] vin0_consume_en_1677;
  wire [0:0] vout_canPeek_1677;
  wire [7:0] vout_peek_1677;
  wire [0:0] v_1678;
  function [0:0] mux_1678(input [0:0] sel);
    case (sel) 0: mux_1678 = 1'h0; 1: mux_1678 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1679;
  wire [0:0] v_1680;
  wire [0:0] v_1681;
  function [0:0] mux_1681(input [0:0] sel);
    case (sel) 0: mux_1681 = 1'h0; 1: mux_1681 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1682;
  wire [0:0] vin0_consume_en_1683;
  wire [0:0] vout_canPeek_1683;
  wire [7:0] vout_peek_1683;
  wire [0:0] v_1684;
  function [0:0] mux_1684(input [0:0] sel);
    case (sel) 0: mux_1684 = 1'h0; 1: mux_1684 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1685;
  wire [0:0] v_1686;
  wire [0:0] v_1687;
  function [0:0] mux_1687(input [0:0] sel);
    case (sel) 0: mux_1687 = 1'h0; 1: mux_1687 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1688;
  wire [0:0] v_1689;
  wire [0:0] v_1690;
  wire [0:0] vin0_consume_en_1691;
  wire [0:0] vout_canPeek_1691;
  wire [7:0] vout_peek_1691;
  wire [0:0] v_1692;
  function [0:0] mux_1692(input [0:0] sel);
    case (sel) 0: mux_1692 = 1'h0; 1: mux_1692 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1693;
  wire [0:0] v_1694;
  wire [0:0] v_1695;
  function [0:0] mux_1695(input [0:0] sel);
    case (sel) 0: mux_1695 = 1'h0; 1: mux_1695 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1696;
  wire [0:0] vin0_consume_en_1697;
  wire [0:0] vout_canPeek_1697;
  wire [7:0] vout_peek_1697;
  wire [0:0] v_1698;
  function [0:0] mux_1698(input [0:0] sel);
    case (sel) 0: mux_1698 = 1'h0; 1: mux_1698 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1699;
  wire [0:0] v_1700;
  wire [0:0] v_1701;
  function [0:0] mux_1701(input [0:0] sel);
    case (sel) 0: mux_1701 = 1'h0; 1: mux_1701 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1702;
  wire [0:0] v_1703;
  wire [0:0] v_1704;
  wire [0:0] vin0_consume_en_1705;
  wire [0:0] vout_canPeek_1705;
  wire [7:0] vout_peek_1705;
  wire [0:0] v_1706;
  function [0:0] mux_1706(input [0:0] sel);
    case (sel) 0: mux_1706 = 1'h0; 1: mux_1706 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1707;
  wire [0:0] v_1708;
  wire [0:0] v_1709;
  function [0:0] mux_1709(input [0:0] sel);
    case (sel) 0: mux_1709 = 1'h0; 1: mux_1709 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1710;
  wire [0:0] vin0_consume_en_1711;
  wire [0:0] vout_canPeek_1711;
  wire [7:0] vout_peek_1711;
  wire [0:0] v_1712;
  function [0:0] mux_1712(input [0:0] sel);
    case (sel) 0: mux_1712 = 1'h0; 1: mux_1712 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1713;
  wire [0:0] v_1714;
  wire [0:0] v_1715;
  function [0:0] mux_1715(input [0:0] sel);
    case (sel) 0: mux_1715 = 1'h0; 1: mux_1715 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1716;
  wire [0:0] v_1717;
  wire [0:0] v_1718;
  wire [0:0] vin0_consume_en_1719;
  wire [0:0] vout_canPeek_1719;
  wire [7:0] vout_peek_1719;
  wire [0:0] v_1720;
  function [0:0] mux_1720(input [0:0] sel);
    case (sel) 0: mux_1720 = 1'h0; 1: mux_1720 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1721;
  wire [0:0] v_1722;
  wire [0:0] v_1723;
  function [0:0] mux_1723(input [0:0] sel);
    case (sel) 0: mux_1723 = 1'h0; 1: mux_1723 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1724;
  wire [0:0] vin0_consume_en_1725;
  wire [0:0] vout_canPeek_1725;
  wire [7:0] vout_peek_1725;
  wire [0:0] v_1726;
  function [0:0] mux_1726(input [0:0] sel);
    case (sel) 0: mux_1726 = 1'h0; 1: mux_1726 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1727;
  wire [0:0] v_1728;
  wire [0:0] v_1729;
  function [0:0] mux_1729(input [0:0] sel);
    case (sel) 0: mux_1729 = 1'h0; 1: mux_1729 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1730;
  wire [0:0] v_1731;
  wire [0:0] v_1732;
  wire [0:0] vin0_consume_en_1733;
  wire [0:0] vout_canPeek_1733;
  wire [7:0] vout_peek_1733;
  wire [0:0] v_1734;
  function [0:0] mux_1734(input [0:0] sel);
    case (sel) 0: mux_1734 = 1'h0; 1: mux_1734 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1735;
  wire [0:0] v_1736;
  wire [0:0] v_1737;
  function [0:0] mux_1737(input [0:0] sel);
    case (sel) 0: mux_1737 = 1'h0; 1: mux_1737 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1738;
  wire [0:0] vin0_consume_en_1739;
  wire [0:0] vout_canPeek_1739;
  wire [7:0] vout_peek_1739;
  wire [0:0] v_1740;
  function [0:0] mux_1740(input [0:0] sel);
    case (sel) 0: mux_1740 = 1'h0; 1: mux_1740 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1741;
  wire [0:0] v_1742;
  wire [0:0] v_1743;
  function [0:0] mux_1743(input [0:0] sel);
    case (sel) 0: mux_1743 = 1'h0; 1: mux_1743 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1744;
  wire [0:0] v_1745;
  wire [0:0] v_1746;
  wire [0:0] vin0_consume_en_1747;
  wire [0:0] vout_canPeek_1747;
  wire [7:0] vout_peek_1747;
  wire [0:0] v_1748;
  function [0:0] mux_1748(input [0:0] sel);
    case (sel) 0: mux_1748 = 1'h0; 1: mux_1748 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1749;
  wire [0:0] v_1750;
  wire [0:0] v_1751;
  function [0:0] mux_1751(input [0:0] sel);
    case (sel) 0: mux_1751 = 1'h0; 1: mux_1751 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1752;
  wire [0:0] vin0_consume_en_1753;
  wire [0:0] vout_canPeek_1753;
  wire [7:0] vout_peek_1753;
  wire [0:0] v_1754;
  function [0:0] mux_1754(input [0:0] sel);
    case (sel) 0: mux_1754 = 1'h0; 1: mux_1754 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1755;
  wire [0:0] v_1756;
  wire [0:0] v_1757;
  function [0:0] mux_1757(input [0:0] sel);
    case (sel) 0: mux_1757 = 1'h0; 1: mux_1757 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1758;
  wire [0:0] v_1759;
  wire [0:0] v_1760;
  wire [0:0] vin0_consume_en_1761;
  wire [0:0] vout_canPeek_1761;
  wire [7:0] vout_peek_1761;
  wire [0:0] v_1762;
  function [0:0] mux_1762(input [0:0] sel);
    case (sel) 0: mux_1762 = 1'h0; 1: mux_1762 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1763;
  wire [0:0] v_1764;
  wire [0:0] v_1765;
  function [0:0] mux_1765(input [0:0] sel);
    case (sel) 0: mux_1765 = 1'h0; 1: mux_1765 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1766;
  wire [0:0] vin0_consume_en_1767;
  wire [0:0] vout_canPeek_1767;
  wire [7:0] vout_peek_1767;
  wire [0:0] v_1768;
  function [0:0] mux_1768(input [0:0] sel);
    case (sel) 0: mux_1768 = 1'h0; 1: mux_1768 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1769;
  wire [0:0] v_1770;
  wire [0:0] v_1771;
  function [0:0] mux_1771(input [0:0] sel);
    case (sel) 0: mux_1771 = 1'h0; 1: mux_1771 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1772;
  wire [0:0] v_1773;
  wire [0:0] v_1774;
  wire [0:0] vin0_consume_en_1775;
  wire [0:0] vout_canPeek_1775;
  wire [7:0] vout_peek_1775;
  wire [0:0] v_1776;
  function [0:0] mux_1776(input [0:0] sel);
    case (sel) 0: mux_1776 = 1'h0; 1: mux_1776 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1777;
  wire [0:0] v_1778;
  wire [0:0] v_1779;
  function [0:0] mux_1779(input [0:0] sel);
    case (sel) 0: mux_1779 = 1'h0; 1: mux_1779 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1780;
  wire [0:0] vin0_consume_en_1781;
  wire [0:0] vout_canPeek_1781;
  wire [7:0] vout_peek_1781;
  wire [0:0] v_1782;
  function [0:0] mux_1782(input [0:0] sel);
    case (sel) 0: mux_1782 = 1'h0; 1: mux_1782 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1783;
  wire [0:0] v_1784;
  wire [0:0] v_1785;
  function [0:0] mux_1785(input [0:0] sel);
    case (sel) 0: mux_1785 = 1'h0; 1: mux_1785 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1786;
  wire [0:0] v_1787;
  wire [0:0] v_1788;
  wire [0:0] vin0_consume_en_1789;
  wire [0:0] vout_canPeek_1789;
  wire [7:0] vout_peek_1789;
  wire [0:0] v_1790;
  function [0:0] mux_1790(input [0:0] sel);
    case (sel) 0: mux_1790 = 1'h0; 1: mux_1790 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1791;
  wire [0:0] v_1792;
  wire [0:0] v_1793;
  function [0:0] mux_1793(input [0:0] sel);
    case (sel) 0: mux_1793 = 1'h0; 1: mux_1793 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1794;
  wire [0:0] vin0_consume_en_1795;
  wire [0:0] vout_canPeek_1795;
  wire [7:0] vout_peek_1795;
  wire [0:0] v_1796;
  function [0:0] mux_1796(input [0:0] sel);
    case (sel) 0: mux_1796 = 1'h0; 1: mux_1796 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1797;
  wire [0:0] v_1798;
  wire [0:0] v_1799;
  function [0:0] mux_1799(input [0:0] sel);
    case (sel) 0: mux_1799 = 1'h0; 1: mux_1799 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1800;
  wire [0:0] v_1801;
  wire [0:0] v_1802;
  wire [0:0] vin0_consume_en_1803;
  wire [0:0] vout_canPeek_1803;
  wire [7:0] vout_peek_1803;
  wire [0:0] v_1804;
  function [0:0] mux_1804(input [0:0] sel);
    case (sel) 0: mux_1804 = 1'h0; 1: mux_1804 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1805;
  wire [0:0] v_1806;
  wire [0:0] v_1807;
  function [0:0] mux_1807(input [0:0] sel);
    case (sel) 0: mux_1807 = 1'h0; 1: mux_1807 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1808;
  wire [0:0] vin0_consume_en_1809;
  wire [0:0] vout_canPeek_1809;
  wire [7:0] vout_peek_1809;
  wire [0:0] v_1810;
  function [0:0] mux_1810(input [0:0] sel);
    case (sel) 0: mux_1810 = 1'h0; 1: mux_1810 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1811;
  wire [0:0] v_1812;
  wire [0:0] v_1813;
  function [0:0] mux_1813(input [0:0] sel);
    case (sel) 0: mux_1813 = 1'h0; 1: mux_1813 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1814;
  wire [0:0] v_1815;
  wire [0:0] v_1816;
  wire [0:0] vin0_consume_en_1817;
  wire [0:0] vout_canPeek_1817;
  wire [7:0] vout_peek_1817;
  wire [0:0] v_1818;
  function [0:0] mux_1818(input [0:0] sel);
    case (sel) 0: mux_1818 = 1'h0; 1: mux_1818 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1819;
  wire [0:0] v_1820;
  wire [0:0] v_1821;
  function [0:0] mux_1821(input [0:0] sel);
    case (sel) 0: mux_1821 = 1'h0; 1: mux_1821 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1822;
  wire [0:0] vin0_consume_en_1823;
  wire [0:0] vout_canPeek_1823;
  wire [7:0] vout_peek_1823;
  wire [0:0] v_1824;
  function [0:0] mux_1824(input [0:0] sel);
    case (sel) 0: mux_1824 = 1'h0; 1: mux_1824 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1825;
  wire [0:0] v_1826;
  wire [0:0] v_1827;
  function [0:0] mux_1827(input [0:0] sel);
    case (sel) 0: mux_1827 = 1'h0; 1: mux_1827 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1828;
  wire [0:0] v_1829;
  wire [0:0] v_1830;
  wire [0:0] vin0_consume_en_1831;
  wire [0:0] vout_canPeek_1831;
  wire [7:0] vout_peek_1831;
  wire [0:0] v_1832;
  function [0:0] mux_1832(input [0:0] sel);
    case (sel) 0: mux_1832 = 1'h0; 1: mux_1832 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1833;
  wire [0:0] v_1834;
  wire [0:0] v_1835;
  function [0:0] mux_1835(input [0:0] sel);
    case (sel) 0: mux_1835 = 1'h0; 1: mux_1835 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1836;
  wire [0:0] vin0_consume_en_1837;
  wire [0:0] vout_canPeek_1837;
  wire [7:0] vout_peek_1837;
  wire [0:0] v_1838;
  function [0:0] mux_1838(input [0:0] sel);
    case (sel) 0: mux_1838 = 1'h0; 1: mux_1838 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1839;
  wire [0:0] v_1840;
  wire [0:0] v_1841;
  function [0:0] mux_1841(input [0:0] sel);
    case (sel) 0: mux_1841 = 1'h0; 1: mux_1841 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1842;
  wire [0:0] v_1843;
  wire [0:0] v_1844;
  wire [0:0] vin0_consume_en_1845;
  wire [0:0] vout_canPeek_1845;
  wire [7:0] vout_peek_1845;
  wire [0:0] v_1846;
  function [0:0] mux_1846(input [0:0] sel);
    case (sel) 0: mux_1846 = 1'h0; 1: mux_1846 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1847;
  wire [0:0] v_1848;
  wire [0:0] v_1849;
  function [0:0] mux_1849(input [0:0] sel);
    case (sel) 0: mux_1849 = 1'h0; 1: mux_1849 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1850;
  wire [0:0] vin0_consume_en_1851;
  wire [0:0] vout_canPeek_1851;
  wire [7:0] vout_peek_1851;
  wire [0:0] v_1852;
  function [0:0] mux_1852(input [0:0] sel);
    case (sel) 0: mux_1852 = 1'h0; 1: mux_1852 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1853;
  wire [0:0] v_1854;
  wire [0:0] v_1855;
  function [0:0] mux_1855(input [0:0] sel);
    case (sel) 0: mux_1855 = 1'h0; 1: mux_1855 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1856;
  wire [0:0] v_1857;
  wire [0:0] v_1858;
  wire [0:0] vin0_consume_en_1859;
  wire [0:0] vout_canPeek_1859;
  wire [7:0] vout_peek_1859;
  wire [0:0] v_1860;
  function [0:0] mux_1860(input [0:0] sel);
    case (sel) 0: mux_1860 = 1'h0; 1: mux_1860 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1861;
  wire [0:0] v_1862;
  wire [0:0] v_1863;
  function [0:0] mux_1863(input [0:0] sel);
    case (sel) 0: mux_1863 = 1'h0; 1: mux_1863 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1864;
  wire [0:0] vin0_consume_en_1865;
  wire [0:0] vout_canPeek_1865;
  wire [7:0] vout_peek_1865;
  wire [0:0] v_1866;
  function [0:0] mux_1866(input [0:0] sel);
    case (sel) 0: mux_1866 = 1'h0; 1: mux_1866 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1867;
  wire [0:0] v_1868;
  wire [0:0] v_1869;
  function [0:0] mux_1869(input [0:0] sel);
    case (sel) 0: mux_1869 = 1'h0; 1: mux_1869 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1870;
  wire [0:0] v_1871;
  wire [0:0] v_1872;
  wire [0:0] vin0_consume_en_1873;
  wire [0:0] vout_canPeek_1873;
  wire [7:0] vout_peek_1873;
  wire [0:0] v_1874;
  function [0:0] mux_1874(input [0:0] sel);
    case (sel) 0: mux_1874 = 1'h0; 1: mux_1874 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1875;
  wire [0:0] v_1876;
  wire [0:0] v_1877;
  function [0:0] mux_1877(input [0:0] sel);
    case (sel) 0: mux_1877 = 1'h0; 1: mux_1877 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1878;
  wire [0:0] vin0_consume_en_1879;
  wire [0:0] vout_canPeek_1879;
  wire [7:0] vout_peek_1879;
  wire [0:0] v_1880;
  function [0:0] mux_1880(input [0:0] sel);
    case (sel) 0: mux_1880 = 1'h0; 1: mux_1880 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1881;
  wire [0:0] v_1882;
  wire [0:0] v_1883;
  function [0:0] mux_1883(input [0:0] sel);
    case (sel) 0: mux_1883 = 1'h0; 1: mux_1883 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1884;
  wire [0:0] v_1885;
  wire [0:0] v_1886;
  wire [0:0] vin0_consume_en_1887;
  wire [0:0] vout_canPeek_1887;
  wire [7:0] vout_peek_1887;
  wire [0:0] v_1888;
  function [0:0] mux_1888(input [0:0] sel);
    case (sel) 0: mux_1888 = 1'h0; 1: mux_1888 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1889;
  wire [0:0] v_1890;
  wire [0:0] v_1891;
  function [0:0] mux_1891(input [0:0] sel);
    case (sel) 0: mux_1891 = 1'h0; 1: mux_1891 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1892;
  wire [0:0] vin0_consume_en_1893;
  wire [0:0] vout_canPeek_1893;
  wire [7:0] vout_peek_1893;
  wire [0:0] v_1894;
  function [0:0] mux_1894(input [0:0] sel);
    case (sel) 0: mux_1894 = 1'h0; 1: mux_1894 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1895;
  wire [0:0] v_1896;
  wire [0:0] v_1897;
  function [0:0] mux_1897(input [0:0] sel);
    case (sel) 0: mux_1897 = 1'h0; 1: mux_1897 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1898;
  wire [0:0] v_1899;
  wire [0:0] v_1900;
  wire [0:0] vin0_consume_en_1901;
  wire [0:0] vout_canPeek_1901;
  wire [7:0] vout_peek_1901;
  wire [0:0] v_1902;
  function [0:0] mux_1902(input [0:0] sel);
    case (sel) 0: mux_1902 = 1'h0; 1: mux_1902 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1903;
  wire [0:0] v_1904;
  wire [0:0] v_1905;
  function [0:0] mux_1905(input [0:0] sel);
    case (sel) 0: mux_1905 = 1'h0; 1: mux_1905 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1906;
  wire [0:0] vin0_consume_en_1907;
  wire [0:0] vout_canPeek_1907;
  wire [7:0] vout_peek_1907;
  wire [0:0] v_1908;
  function [0:0] mux_1908(input [0:0] sel);
    case (sel) 0: mux_1908 = 1'h0; 1: mux_1908 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1909;
  wire [0:0] v_1910;
  wire [0:0] v_1911;
  function [0:0] mux_1911(input [0:0] sel);
    case (sel) 0: mux_1911 = 1'h0; 1: mux_1911 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1912;
  wire [0:0] v_1913;
  wire [0:0] v_1914;
  wire [0:0] vin0_consume_en_1915;
  wire [0:0] vout_canPeek_1915;
  wire [7:0] vout_peek_1915;
  wire [0:0] v_1916;
  function [0:0] mux_1916(input [0:0] sel);
    case (sel) 0: mux_1916 = 1'h0; 1: mux_1916 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1917;
  wire [0:0] v_1918;
  wire [0:0] v_1919;
  function [0:0] mux_1919(input [0:0] sel);
    case (sel) 0: mux_1919 = 1'h0; 1: mux_1919 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1920;
  wire [0:0] vin0_consume_en_1921;
  wire [0:0] vout_canPeek_1921;
  wire [7:0] vout_peek_1921;
  wire [0:0] v_1922;
  function [0:0] mux_1922(input [0:0] sel);
    case (sel) 0: mux_1922 = 1'h0; 1: mux_1922 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1923;
  wire [0:0] v_1924;
  wire [0:0] v_1925;
  function [0:0] mux_1925(input [0:0] sel);
    case (sel) 0: mux_1925 = 1'h0; 1: mux_1925 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1926;
  wire [0:0] v_1927;
  wire [0:0] v_1928;
  wire [0:0] vin0_consume_en_1929;
  wire [0:0] vout_canPeek_1929;
  wire [7:0] vout_peek_1929;
  wire [0:0] v_1930;
  function [0:0] mux_1930(input [0:0] sel);
    case (sel) 0: mux_1930 = 1'h0; 1: mux_1930 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1931;
  wire [0:0] v_1932;
  wire [0:0] v_1933;
  function [0:0] mux_1933(input [0:0] sel);
    case (sel) 0: mux_1933 = 1'h0; 1: mux_1933 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1934;
  wire [0:0] vin0_consume_en_1935;
  wire [0:0] vout_canPeek_1935;
  wire [7:0] vout_peek_1935;
  wire [0:0] v_1936;
  function [0:0] mux_1936(input [0:0] sel);
    case (sel) 0: mux_1936 = 1'h0; 1: mux_1936 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1937;
  wire [0:0] v_1938;
  wire [0:0] v_1939;
  function [0:0] mux_1939(input [0:0] sel);
    case (sel) 0: mux_1939 = 1'h0; 1: mux_1939 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1940;
  wire [0:0] v_1941;
  wire [0:0] v_1942;
  wire [0:0] vin0_consume_en_1943;
  wire [0:0] vout_canPeek_1943;
  wire [7:0] vout_peek_1943;
  wire [0:0] v_1944;
  function [0:0] mux_1944(input [0:0] sel);
    case (sel) 0: mux_1944 = 1'h0; 1: mux_1944 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1945;
  wire [0:0] v_1946;
  wire [0:0] v_1947;
  function [0:0] mux_1947(input [0:0] sel);
    case (sel) 0: mux_1947 = 1'h0; 1: mux_1947 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1948;
  wire [0:0] vin0_consume_en_1949;
  wire [0:0] vout_canPeek_1949;
  wire [7:0] vout_peek_1949;
  wire [0:0] v_1950;
  function [0:0] mux_1950(input [0:0] sel);
    case (sel) 0: mux_1950 = 1'h0; 1: mux_1950 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1951;
  wire [0:0] v_1952;
  wire [0:0] v_1953;
  function [0:0] mux_1953(input [0:0] sel);
    case (sel) 0: mux_1953 = 1'h0; 1: mux_1953 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1954;
  wire [0:0] v_1955;
  wire [0:0] v_1956;
  wire [0:0] vin0_consume_en_1957;
  wire [0:0] vout_canPeek_1957;
  wire [7:0] vout_peek_1957;
  wire [0:0] v_1958;
  function [0:0] mux_1958(input [0:0] sel);
    case (sel) 0: mux_1958 = 1'h0; 1: mux_1958 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1959;
  wire [0:0] v_1960;
  wire [0:0] v_1961;
  function [0:0] mux_1961(input [0:0] sel);
    case (sel) 0: mux_1961 = 1'h0; 1: mux_1961 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1962;
  wire [0:0] vin0_consume_en_1963;
  wire [0:0] vout_canPeek_1963;
  wire [7:0] vout_peek_1963;
  wire [0:0] v_1964;
  function [0:0] mux_1964(input [0:0] sel);
    case (sel) 0: mux_1964 = 1'h0; 1: mux_1964 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1965;
  wire [0:0] v_1966;
  wire [0:0] v_1967;
  function [0:0] mux_1967(input [0:0] sel);
    case (sel) 0: mux_1967 = 1'h0; 1: mux_1967 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1968;
  wire [0:0] v_1969;
  wire [0:0] v_1970;
  wire [0:0] vin0_consume_en_1971;
  wire [0:0] vout_canPeek_1971;
  wire [7:0] vout_peek_1971;
  wire [0:0] v_1972;
  function [0:0] mux_1972(input [0:0] sel);
    case (sel) 0: mux_1972 = 1'h0; 1: mux_1972 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1973;
  wire [0:0] v_1974;
  wire [0:0] v_1975;
  function [0:0] mux_1975(input [0:0] sel);
    case (sel) 0: mux_1975 = 1'h0; 1: mux_1975 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1976;
  wire [0:0] vin0_consume_en_1977;
  wire [0:0] vout_canPeek_1977;
  wire [7:0] vout_peek_1977;
  wire [0:0] v_1978;
  function [0:0] mux_1978(input [0:0] sel);
    case (sel) 0: mux_1978 = 1'h0; 1: mux_1978 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1979;
  wire [0:0] v_1980;
  wire [0:0] v_1981;
  function [0:0] mux_1981(input [0:0] sel);
    case (sel) 0: mux_1981 = 1'h0; 1: mux_1981 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1982;
  wire [0:0] v_1983;
  wire [0:0] v_1984;
  wire [0:0] vin0_consume_en_1985;
  wire [0:0] vout_canPeek_1985;
  wire [7:0] vout_peek_1985;
  wire [0:0] v_1986;
  function [0:0] mux_1986(input [0:0] sel);
    case (sel) 0: mux_1986 = 1'h0; 1: mux_1986 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1987;
  wire [0:0] v_1988;
  wire [0:0] v_1989;
  function [0:0] mux_1989(input [0:0] sel);
    case (sel) 0: mux_1989 = 1'h0; 1: mux_1989 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1990;
  wire [0:0] vin0_consume_en_1991;
  wire [0:0] vout_canPeek_1991;
  wire [7:0] vout_peek_1991;
  wire [0:0] v_1992;
  function [0:0] mux_1992(input [0:0] sel);
    case (sel) 0: mux_1992 = 1'h0; 1: mux_1992 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_1993;
  wire [0:0] v_1994;
  wire [0:0] v_1995;
  function [0:0] mux_1995(input [0:0] sel);
    case (sel) 0: mux_1995 = 1'h0; 1: mux_1995 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_1996;
  wire [0:0] v_1997;
  wire [0:0] v_1998;
  wire [0:0] vin0_consume_en_1999;
  wire [0:0] vout_canPeek_1999;
  wire [7:0] vout_peek_1999;
  wire [0:0] v_2000;
  function [0:0] mux_2000(input [0:0] sel);
    case (sel) 0: mux_2000 = 1'h0; 1: mux_2000 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2001;
  wire [0:0] v_2002;
  wire [0:0] v_2003;
  function [0:0] mux_2003(input [0:0] sel);
    case (sel) 0: mux_2003 = 1'h0; 1: mux_2003 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2004;
  wire [0:0] vin0_consume_en_2005;
  wire [0:0] vout_canPeek_2005;
  wire [7:0] vout_peek_2005;
  wire [0:0] v_2006;
  function [0:0] mux_2006(input [0:0] sel);
    case (sel) 0: mux_2006 = 1'h0; 1: mux_2006 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2007;
  wire [0:0] v_2008;
  wire [0:0] v_2009;
  function [0:0] mux_2009(input [0:0] sel);
    case (sel) 0: mux_2009 = 1'h0; 1: mux_2009 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2010;
  wire [0:0] v_2011;
  wire [0:0] v_2012;
  wire [0:0] vin0_consume_en_2013;
  wire [0:0] vout_canPeek_2013;
  wire [7:0] vout_peek_2013;
  wire [0:0] v_2014;
  function [0:0] mux_2014(input [0:0] sel);
    case (sel) 0: mux_2014 = 1'h0; 1: mux_2014 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2015;
  wire [0:0] v_2016;
  wire [0:0] v_2017;
  function [0:0] mux_2017(input [0:0] sel);
    case (sel) 0: mux_2017 = 1'h0; 1: mux_2017 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2018;
  wire [0:0] vin0_consume_en_2019;
  wire [0:0] vout_canPeek_2019;
  wire [7:0] vout_peek_2019;
  wire [0:0] v_2020;
  function [0:0] mux_2020(input [0:0] sel);
    case (sel) 0: mux_2020 = 1'h0; 1: mux_2020 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2021;
  wire [0:0] v_2022;
  wire [0:0] v_2023;
  function [0:0] mux_2023(input [0:0] sel);
    case (sel) 0: mux_2023 = 1'h0; 1: mux_2023 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2024;
  wire [0:0] v_2025;
  wire [0:0] v_2026;
  wire [0:0] vin0_consume_en_2027;
  wire [0:0] vout_canPeek_2027;
  wire [7:0] vout_peek_2027;
  wire [0:0] v_2028;
  function [0:0] mux_2028(input [0:0] sel);
    case (sel) 0: mux_2028 = 1'h0; 1: mux_2028 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2029;
  wire [0:0] v_2030;
  wire [0:0] v_2031;
  function [0:0] mux_2031(input [0:0] sel);
    case (sel) 0: mux_2031 = 1'h0; 1: mux_2031 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2032;
  wire [0:0] vin0_consume_en_2033;
  wire [0:0] vout_canPeek_2033;
  wire [7:0] vout_peek_2033;
  wire [0:0] v_2034;
  function [0:0] mux_2034(input [0:0] sel);
    case (sel) 0: mux_2034 = 1'h0; 1: mux_2034 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2035;
  wire [0:0] v_2036;
  wire [0:0] v_2037;
  function [0:0] mux_2037(input [0:0] sel);
    case (sel) 0: mux_2037 = 1'h0; 1: mux_2037 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2038;
  wire [0:0] v_2039;
  wire [0:0] v_2040;
  wire [0:0] vin0_consume_en_2041;
  wire [0:0] vout_canPeek_2041;
  wire [7:0] vout_peek_2041;
  wire [0:0] v_2042;
  function [0:0] mux_2042(input [0:0] sel);
    case (sel) 0: mux_2042 = 1'h0; 1: mux_2042 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2043;
  wire [0:0] v_2044;
  wire [0:0] v_2045;
  function [0:0] mux_2045(input [0:0] sel);
    case (sel) 0: mux_2045 = 1'h0; 1: mux_2045 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2046;
  wire [0:0] vin0_consume_en_2047;
  wire [0:0] vout_canPeek_2047;
  wire [7:0] vout_peek_2047;
  wire [0:0] v_2048;
  function [0:0] mux_2048(input [0:0] sel);
    case (sel) 0: mux_2048 = 1'h0; 1: mux_2048 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2049;
  wire [0:0] v_2050;
  wire [0:0] v_2051;
  function [0:0] mux_2051(input [0:0] sel);
    case (sel) 0: mux_2051 = 1'h0; 1: mux_2051 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2052;
  wire [0:0] v_2053;
  wire [0:0] v_2054;
  wire [0:0] vin0_consume_en_2055;
  wire [0:0] vout_canPeek_2055;
  wire [7:0] vout_peek_2055;
  wire [0:0] v_2056;
  function [0:0] mux_2056(input [0:0] sel);
    case (sel) 0: mux_2056 = 1'h0; 1: mux_2056 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2057;
  wire [0:0] v_2058;
  wire [0:0] v_2059;
  function [0:0] mux_2059(input [0:0] sel);
    case (sel) 0: mux_2059 = 1'h0; 1: mux_2059 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2060;
  wire [0:0] vin0_consume_en_2061;
  wire [0:0] vout_canPeek_2061;
  wire [7:0] vout_peek_2061;
  wire [0:0] v_2062;
  function [0:0] mux_2062(input [0:0] sel);
    case (sel) 0: mux_2062 = 1'h0; 1: mux_2062 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2063;
  wire [0:0] v_2064;
  wire [0:0] v_2065;
  function [0:0] mux_2065(input [0:0] sel);
    case (sel) 0: mux_2065 = 1'h0; 1: mux_2065 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2066;
  wire [0:0] v_2067;
  wire [0:0] v_2068;
  wire [0:0] vin0_consume_en_2069;
  wire [0:0] vout_canPeek_2069;
  wire [7:0] vout_peek_2069;
  wire [0:0] v_2070;
  function [0:0] mux_2070(input [0:0] sel);
    case (sel) 0: mux_2070 = 1'h0; 1: mux_2070 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2071;
  wire [0:0] v_2072;
  wire [0:0] v_2073;
  function [0:0] mux_2073(input [0:0] sel);
    case (sel) 0: mux_2073 = 1'h0; 1: mux_2073 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2074;
  wire [0:0] vin0_consume_en_2075;
  wire [0:0] vout_canPeek_2075;
  wire [7:0] vout_peek_2075;
  wire [0:0] v_2076;
  function [0:0] mux_2076(input [0:0] sel);
    case (sel) 0: mux_2076 = 1'h0; 1: mux_2076 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2077;
  wire [0:0] v_2078;
  wire [0:0] v_2079;
  function [0:0] mux_2079(input [0:0] sel);
    case (sel) 0: mux_2079 = 1'h0; 1: mux_2079 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2080;
  wire [0:0] v_2081;
  wire [0:0] v_2082;
  wire [0:0] vin0_consume_en_2083;
  wire [0:0] vout_canPeek_2083;
  wire [7:0] vout_peek_2083;
  wire [0:0] v_2084;
  function [0:0] mux_2084(input [0:0] sel);
    case (sel) 0: mux_2084 = 1'h0; 1: mux_2084 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2085;
  wire [0:0] v_2086;
  wire [0:0] v_2087;
  function [0:0] mux_2087(input [0:0] sel);
    case (sel) 0: mux_2087 = 1'h0; 1: mux_2087 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2088;
  wire [0:0] vin0_consume_en_2089;
  wire [0:0] vout_canPeek_2089;
  wire [7:0] vout_peek_2089;
  wire [0:0] v_2090;
  function [0:0] mux_2090(input [0:0] sel);
    case (sel) 0: mux_2090 = 1'h0; 1: mux_2090 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2091;
  wire [0:0] v_2092;
  wire [0:0] v_2093;
  function [0:0] mux_2093(input [0:0] sel);
    case (sel) 0: mux_2093 = 1'h0; 1: mux_2093 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2094;
  wire [0:0] v_2095;
  wire [0:0] v_2096;
  wire [0:0] vin0_consume_en_2097;
  wire [0:0] vout_canPeek_2097;
  wire [7:0] vout_peek_2097;
  wire [0:0] v_2098;
  function [0:0] mux_2098(input [0:0] sel);
    case (sel) 0: mux_2098 = 1'h0; 1: mux_2098 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2099;
  wire [0:0] v_2100;
  wire [0:0] v_2101;
  function [0:0] mux_2101(input [0:0] sel);
    case (sel) 0: mux_2101 = 1'h0; 1: mux_2101 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2102;
  wire [0:0] vin0_consume_en_2103;
  wire [0:0] vout_canPeek_2103;
  wire [7:0] vout_peek_2103;
  wire [0:0] v_2104;
  function [0:0] mux_2104(input [0:0] sel);
    case (sel) 0: mux_2104 = 1'h0; 1: mux_2104 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2105;
  wire [0:0] v_2106;
  wire [0:0] v_2107;
  function [0:0] mux_2107(input [0:0] sel);
    case (sel) 0: mux_2107 = 1'h0; 1: mux_2107 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2108;
  wire [0:0] v_2109;
  wire [0:0] v_2110;
  wire [0:0] vin0_consume_en_2111;
  wire [0:0] vout_canPeek_2111;
  wire [7:0] vout_peek_2111;
  wire [0:0] v_2112;
  function [0:0] mux_2112(input [0:0] sel);
    case (sel) 0: mux_2112 = 1'h0; 1: mux_2112 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2113;
  wire [0:0] v_2114;
  wire [0:0] v_2115;
  function [0:0] mux_2115(input [0:0] sel);
    case (sel) 0: mux_2115 = 1'h0; 1: mux_2115 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2116;
  wire [0:0] vin0_consume_en_2117;
  wire [0:0] vout_canPeek_2117;
  wire [7:0] vout_peek_2117;
  wire [0:0] v_2118;
  function [0:0] mux_2118(input [0:0] sel);
    case (sel) 0: mux_2118 = 1'h0; 1: mux_2118 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2119;
  wire [0:0] v_2120;
  wire [0:0] v_2121;
  function [0:0] mux_2121(input [0:0] sel);
    case (sel) 0: mux_2121 = 1'h0; 1: mux_2121 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2122;
  wire [0:0] v_2123;
  wire [0:0] v_2124;
  wire [0:0] vin0_consume_en_2125;
  wire [0:0] vout_canPeek_2125;
  wire [7:0] vout_peek_2125;
  wire [0:0] v_2126;
  function [0:0] mux_2126(input [0:0] sel);
    case (sel) 0: mux_2126 = 1'h0; 1: mux_2126 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2127;
  wire [0:0] v_2128;
  wire [0:0] v_2129;
  function [0:0] mux_2129(input [0:0] sel);
    case (sel) 0: mux_2129 = 1'h0; 1: mux_2129 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2130;
  wire [0:0] vin0_consume_en_2131;
  wire [0:0] vout_canPeek_2131;
  wire [7:0] vout_peek_2131;
  wire [0:0] v_2132;
  function [0:0] mux_2132(input [0:0] sel);
    case (sel) 0: mux_2132 = 1'h0; 1: mux_2132 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2133;
  wire [0:0] v_2134;
  wire [0:0] v_2135;
  function [0:0] mux_2135(input [0:0] sel);
    case (sel) 0: mux_2135 = 1'h0; 1: mux_2135 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2136;
  wire [0:0] v_2137;
  wire [0:0] v_2138;
  wire [0:0] vin0_consume_en_2139;
  wire [0:0] vout_canPeek_2139;
  wire [7:0] vout_peek_2139;
  wire [0:0] v_2140;
  function [0:0] mux_2140(input [0:0] sel);
    case (sel) 0: mux_2140 = 1'h0; 1: mux_2140 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2141;
  wire [0:0] v_2142;
  wire [0:0] v_2143;
  function [0:0] mux_2143(input [0:0] sel);
    case (sel) 0: mux_2143 = 1'h0; 1: mux_2143 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2144;
  wire [0:0] vin0_consume_en_2145;
  wire [0:0] vout_canPeek_2145;
  wire [7:0] vout_peek_2145;
  wire [0:0] v_2146;
  function [0:0] mux_2146(input [0:0] sel);
    case (sel) 0: mux_2146 = 1'h0; 1: mux_2146 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2147;
  wire [0:0] v_2148;
  wire [0:0] v_2149;
  function [0:0] mux_2149(input [0:0] sel);
    case (sel) 0: mux_2149 = 1'h0; 1: mux_2149 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2150;
  wire [0:0] v_2151;
  wire [0:0] v_2152;
  wire [0:0] vin0_consume_en_2153;
  wire [0:0] vout_canPeek_2153;
  wire [7:0] vout_peek_2153;
  wire [0:0] v_2154;
  function [0:0] mux_2154(input [0:0] sel);
    case (sel) 0: mux_2154 = 1'h0; 1: mux_2154 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2155;
  wire [0:0] v_2156;
  wire [0:0] v_2157;
  function [0:0] mux_2157(input [0:0] sel);
    case (sel) 0: mux_2157 = 1'h0; 1: mux_2157 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2158;
  wire [0:0] vin0_consume_en_2159;
  wire [0:0] vout_canPeek_2159;
  wire [7:0] vout_peek_2159;
  wire [0:0] v_2160;
  function [0:0] mux_2160(input [0:0] sel);
    case (sel) 0: mux_2160 = 1'h0; 1: mux_2160 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2161;
  wire [0:0] v_2162;
  wire [0:0] v_2163;
  function [0:0] mux_2163(input [0:0] sel);
    case (sel) 0: mux_2163 = 1'h0; 1: mux_2163 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2164;
  wire [0:0] v_2165;
  wire [0:0] v_2166;
  wire [0:0] vin0_consume_en_2167;
  wire [0:0] vout_canPeek_2167;
  wire [7:0] vout_peek_2167;
  wire [0:0] v_2168;
  function [0:0] mux_2168(input [0:0] sel);
    case (sel) 0: mux_2168 = 1'h0; 1: mux_2168 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2169;
  wire [0:0] v_2170;
  wire [0:0] v_2171;
  function [0:0] mux_2171(input [0:0] sel);
    case (sel) 0: mux_2171 = 1'h0; 1: mux_2171 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2172;
  wire [0:0] vin0_consume_en_2173;
  wire [0:0] vout_canPeek_2173;
  wire [7:0] vout_peek_2173;
  wire [0:0] v_2174;
  function [0:0] mux_2174(input [0:0] sel);
    case (sel) 0: mux_2174 = 1'h0; 1: mux_2174 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2175;
  wire [0:0] v_2176;
  wire [0:0] v_2177;
  function [0:0] mux_2177(input [0:0] sel);
    case (sel) 0: mux_2177 = 1'h0; 1: mux_2177 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2178;
  wire [0:0] v_2179;
  wire [0:0] v_2180;
  wire [0:0] vin0_consume_en_2181;
  wire [0:0] vout_canPeek_2181;
  wire [7:0] vout_peek_2181;
  wire [0:0] v_2182;
  function [0:0] mux_2182(input [0:0] sel);
    case (sel) 0: mux_2182 = 1'h0; 1: mux_2182 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2183;
  wire [0:0] v_2184;
  wire [0:0] v_2185;
  function [0:0] mux_2185(input [0:0] sel);
    case (sel) 0: mux_2185 = 1'h0; 1: mux_2185 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2186;
  wire [0:0] vin0_consume_en_2187;
  wire [0:0] vout_canPeek_2187;
  wire [7:0] vout_peek_2187;
  wire [0:0] v_2188;
  function [0:0] mux_2188(input [0:0] sel);
    case (sel) 0: mux_2188 = 1'h0; 1: mux_2188 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2189;
  wire [0:0] v_2190;
  wire [0:0] v_2191;
  function [0:0] mux_2191(input [0:0] sel);
    case (sel) 0: mux_2191 = 1'h0; 1: mux_2191 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2192;
  wire [0:0] v_2193;
  wire [0:0] v_2194;
  wire [0:0] vin0_consume_en_2195;
  wire [0:0] vout_canPeek_2195;
  wire [7:0] vout_peek_2195;
  wire [0:0] v_2196;
  function [0:0] mux_2196(input [0:0] sel);
    case (sel) 0: mux_2196 = 1'h0; 1: mux_2196 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2197;
  wire [0:0] v_2198;
  wire [0:0] v_2199;
  function [0:0] mux_2199(input [0:0] sel);
    case (sel) 0: mux_2199 = 1'h0; 1: mux_2199 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2200;
  wire [0:0] vin0_consume_en_2201;
  wire [0:0] vout_canPeek_2201;
  wire [7:0] vout_peek_2201;
  wire [0:0] v_2202;
  function [0:0] mux_2202(input [0:0] sel);
    case (sel) 0: mux_2202 = 1'h0; 1: mux_2202 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2203;
  wire [0:0] v_2204;
  wire [0:0] v_2205;
  function [0:0] mux_2205(input [0:0] sel);
    case (sel) 0: mux_2205 = 1'h0; 1: mux_2205 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2206;
  wire [0:0] v_2207;
  wire [0:0] v_2208;
  wire [0:0] vin0_consume_en_2209;
  wire [0:0] vout_canPeek_2209;
  wire [7:0] vout_peek_2209;
  wire [0:0] v_2210;
  function [0:0] mux_2210(input [0:0] sel);
    case (sel) 0: mux_2210 = 1'h0; 1: mux_2210 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2211;
  wire [0:0] v_2212;
  wire [0:0] v_2213;
  function [0:0] mux_2213(input [0:0] sel);
    case (sel) 0: mux_2213 = 1'h0; 1: mux_2213 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2214;
  wire [0:0] vin0_consume_en_2215;
  wire [0:0] vout_canPeek_2215;
  wire [7:0] vout_peek_2215;
  wire [0:0] v_2216;
  function [0:0] mux_2216(input [0:0] sel);
    case (sel) 0: mux_2216 = 1'h0; 1: mux_2216 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2217;
  wire [0:0] v_2218;
  wire [0:0] v_2219;
  function [0:0] mux_2219(input [0:0] sel);
    case (sel) 0: mux_2219 = 1'h0; 1: mux_2219 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2220;
  wire [0:0] v_2221;
  wire [0:0] v_2222;
  wire [0:0] vin0_consume_en_2223;
  wire [0:0] vout_canPeek_2223;
  wire [7:0] vout_peek_2223;
  wire [0:0] v_2224;
  function [0:0] mux_2224(input [0:0] sel);
    case (sel) 0: mux_2224 = 1'h0; 1: mux_2224 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2225;
  wire [0:0] v_2226;
  wire [0:0] v_2227;
  function [0:0] mux_2227(input [0:0] sel);
    case (sel) 0: mux_2227 = 1'h0; 1: mux_2227 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2228;
  wire [0:0] vin0_consume_en_2229;
  wire [0:0] vout_canPeek_2229;
  wire [7:0] vout_peek_2229;
  wire [0:0] v_2230;
  function [0:0] mux_2230(input [0:0] sel);
    case (sel) 0: mux_2230 = 1'h0; 1: mux_2230 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2231;
  wire [0:0] v_2232;
  wire [0:0] v_2233;
  function [0:0] mux_2233(input [0:0] sel);
    case (sel) 0: mux_2233 = 1'h0; 1: mux_2233 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2234;
  wire [0:0] v_2235;
  wire [0:0] v_2236;
  wire [0:0] vin0_consume_en_2237;
  wire [0:0] vout_canPeek_2237;
  wire [7:0] vout_peek_2237;
  wire [0:0] v_2238;
  function [0:0] mux_2238(input [0:0] sel);
    case (sel) 0: mux_2238 = 1'h0; 1: mux_2238 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2239;
  wire [0:0] v_2240;
  wire [0:0] v_2241;
  function [0:0] mux_2241(input [0:0] sel);
    case (sel) 0: mux_2241 = 1'h0; 1: mux_2241 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2242;
  wire [0:0] vin0_consume_en_2243;
  wire [0:0] vout_canPeek_2243;
  wire [7:0] vout_peek_2243;
  wire [0:0] v_2244;
  function [0:0] mux_2244(input [0:0] sel);
    case (sel) 0: mux_2244 = 1'h0; 1: mux_2244 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2245;
  wire [0:0] v_2246;
  wire [0:0] v_2247;
  function [0:0] mux_2247(input [0:0] sel);
    case (sel) 0: mux_2247 = 1'h0; 1: mux_2247 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2248;
  wire [0:0] v_2249;
  wire [0:0] v_2250;
  wire [0:0] vin0_consume_en_2251;
  wire [0:0] vout_canPeek_2251;
  wire [7:0] vout_peek_2251;
  wire [0:0] v_2252;
  function [0:0] mux_2252(input [0:0] sel);
    case (sel) 0: mux_2252 = 1'h0; 1: mux_2252 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2253;
  wire [0:0] v_2254;
  wire [0:0] v_2255;
  function [0:0] mux_2255(input [0:0] sel);
    case (sel) 0: mux_2255 = 1'h0; 1: mux_2255 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2256;
  wire [0:0] vin0_consume_en_2257;
  wire [0:0] vout_canPeek_2257;
  wire [7:0] vout_peek_2257;
  wire [0:0] v_2258;
  function [0:0] mux_2258(input [0:0] sel);
    case (sel) 0: mux_2258 = 1'h0; 1: mux_2258 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2259;
  wire [0:0] v_2260;
  wire [0:0] v_2261;
  function [0:0] mux_2261(input [0:0] sel);
    case (sel) 0: mux_2261 = 1'h0; 1: mux_2261 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2262;
  wire [0:0] v_2263;
  wire [0:0] v_2264;
  wire [0:0] vin0_consume_en_2265;
  wire [0:0] vout_canPeek_2265;
  wire [7:0] vout_peek_2265;
  wire [0:0] v_2266;
  function [0:0] mux_2266(input [0:0] sel);
    case (sel) 0: mux_2266 = 1'h0; 1: mux_2266 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2267;
  wire [0:0] v_2268;
  wire [0:0] v_2269;
  function [0:0] mux_2269(input [0:0] sel);
    case (sel) 0: mux_2269 = 1'h0; 1: mux_2269 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2270;
  wire [0:0] vin0_consume_en_2271;
  wire [0:0] vout_canPeek_2271;
  wire [7:0] vout_peek_2271;
  wire [0:0] v_2272;
  function [0:0] mux_2272(input [0:0] sel);
    case (sel) 0: mux_2272 = 1'h0; 1: mux_2272 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2273;
  wire [0:0] v_2274;
  wire [0:0] v_2275;
  function [0:0] mux_2275(input [0:0] sel);
    case (sel) 0: mux_2275 = 1'h0; 1: mux_2275 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2276;
  wire [0:0] v_2277;
  wire [0:0] v_2278;
  wire [0:0] vin0_consume_en_2279;
  wire [0:0] vout_canPeek_2279;
  wire [7:0] vout_peek_2279;
  wire [0:0] v_2280;
  function [0:0] mux_2280(input [0:0] sel);
    case (sel) 0: mux_2280 = 1'h0; 1: mux_2280 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2281;
  wire [0:0] v_2282;
  wire [0:0] v_2283;
  function [0:0] mux_2283(input [0:0] sel);
    case (sel) 0: mux_2283 = 1'h0; 1: mux_2283 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2284;
  wire [0:0] vin0_consume_en_2285;
  wire [0:0] vout_canPeek_2285;
  wire [7:0] vout_peek_2285;
  wire [0:0] v_2286;
  function [0:0] mux_2286(input [0:0] sel);
    case (sel) 0: mux_2286 = 1'h0; 1: mux_2286 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2287;
  wire [0:0] v_2288;
  wire [0:0] v_2289;
  function [0:0] mux_2289(input [0:0] sel);
    case (sel) 0: mux_2289 = 1'h0; 1: mux_2289 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2290;
  wire [0:0] v_2291;
  wire [0:0] v_2292;
  wire [0:0] vin0_consume_en_2293;
  wire [0:0] vout_canPeek_2293;
  wire [7:0] vout_peek_2293;
  wire [0:0] v_2294;
  function [0:0] mux_2294(input [0:0] sel);
    case (sel) 0: mux_2294 = 1'h0; 1: mux_2294 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2295;
  wire [0:0] v_2296;
  wire [0:0] v_2297;
  function [0:0] mux_2297(input [0:0] sel);
    case (sel) 0: mux_2297 = 1'h0; 1: mux_2297 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2298;
  wire [0:0] vin0_consume_en_2299;
  wire [0:0] vout_canPeek_2299;
  wire [7:0] vout_peek_2299;
  wire [0:0] v_2300;
  function [0:0] mux_2300(input [0:0] sel);
    case (sel) 0: mux_2300 = 1'h0; 1: mux_2300 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2301;
  wire [0:0] v_2302;
  wire [0:0] v_2303;
  function [0:0] mux_2303(input [0:0] sel);
    case (sel) 0: mux_2303 = 1'h0; 1: mux_2303 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2304;
  wire [0:0] v_2305;
  wire [0:0] v_2306;
  wire [0:0] vin0_consume_en_2307;
  wire [0:0] vout_canPeek_2307;
  wire [7:0] vout_peek_2307;
  wire [0:0] v_2308;
  function [0:0] mux_2308(input [0:0] sel);
    case (sel) 0: mux_2308 = 1'h0; 1: mux_2308 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2309;
  wire [0:0] v_2310;
  wire [0:0] v_2311;
  function [0:0] mux_2311(input [0:0] sel);
    case (sel) 0: mux_2311 = 1'h0; 1: mux_2311 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2312;
  wire [0:0] vin0_consume_en_2313;
  wire [0:0] vout_canPeek_2313;
  wire [7:0] vout_peek_2313;
  wire [0:0] v_2314;
  function [0:0] mux_2314(input [0:0] sel);
    case (sel) 0: mux_2314 = 1'h0; 1: mux_2314 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2315;
  wire [0:0] v_2316;
  wire [0:0] v_2317;
  function [0:0] mux_2317(input [0:0] sel);
    case (sel) 0: mux_2317 = 1'h0; 1: mux_2317 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2318;
  wire [0:0] v_2319;
  wire [0:0] v_2320;
  wire [0:0] vin0_consume_en_2321;
  wire [0:0] vout_canPeek_2321;
  wire [7:0] vout_peek_2321;
  wire [0:0] v_2322;
  function [0:0] mux_2322(input [0:0] sel);
    case (sel) 0: mux_2322 = 1'h0; 1: mux_2322 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2323;
  wire [0:0] v_2324;
  wire [0:0] v_2325;
  function [0:0] mux_2325(input [0:0] sel);
    case (sel) 0: mux_2325 = 1'h0; 1: mux_2325 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2326;
  wire [0:0] vin0_consume_en_2327;
  wire [0:0] vout_canPeek_2327;
  wire [7:0] vout_peek_2327;
  wire [0:0] v_2328;
  function [0:0] mux_2328(input [0:0] sel);
    case (sel) 0: mux_2328 = 1'h0; 1: mux_2328 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2329;
  wire [0:0] v_2330;
  wire [0:0] v_2331;
  function [0:0] mux_2331(input [0:0] sel);
    case (sel) 0: mux_2331 = 1'h0; 1: mux_2331 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2332;
  wire [0:0] v_2333;
  wire [0:0] v_2334;
  wire [0:0] vin0_consume_en_2335;
  wire [0:0] vout_canPeek_2335;
  wire [7:0] vout_peek_2335;
  wire [0:0] v_2336;
  function [0:0] mux_2336(input [0:0] sel);
    case (sel) 0: mux_2336 = 1'h0; 1: mux_2336 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2337;
  wire [0:0] v_2338;
  wire [0:0] v_2339;
  function [0:0] mux_2339(input [0:0] sel);
    case (sel) 0: mux_2339 = 1'h0; 1: mux_2339 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2340;
  wire [0:0] vin0_consume_en_2341;
  wire [0:0] vout_canPeek_2341;
  wire [7:0] vout_peek_2341;
  wire [0:0] v_2342;
  function [0:0] mux_2342(input [0:0] sel);
    case (sel) 0: mux_2342 = 1'h0; 1: mux_2342 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2343;
  wire [0:0] v_2344;
  wire [0:0] v_2345;
  function [0:0] mux_2345(input [0:0] sel);
    case (sel) 0: mux_2345 = 1'h0; 1: mux_2345 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2346;
  wire [0:0] v_2347;
  wire [0:0] v_2348;
  wire [0:0] vin0_consume_en_2349;
  wire [0:0] vout_canPeek_2349;
  wire [7:0] vout_peek_2349;
  wire [0:0] v_2350;
  function [0:0] mux_2350(input [0:0] sel);
    case (sel) 0: mux_2350 = 1'h0; 1: mux_2350 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2351;
  wire [0:0] v_2352;
  wire [0:0] v_2353;
  function [0:0] mux_2353(input [0:0] sel);
    case (sel) 0: mux_2353 = 1'h0; 1: mux_2353 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2354;
  wire [0:0] vin0_consume_en_2355;
  wire [0:0] vout_canPeek_2355;
  wire [7:0] vout_peek_2355;
  wire [0:0] v_2356;
  function [0:0] mux_2356(input [0:0] sel);
    case (sel) 0: mux_2356 = 1'h0; 1: mux_2356 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2357;
  wire [0:0] v_2358;
  wire [0:0] v_2359;
  function [0:0] mux_2359(input [0:0] sel);
    case (sel) 0: mux_2359 = 1'h0; 1: mux_2359 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2360;
  wire [0:0] v_2361;
  wire [0:0] v_2362;
  wire [0:0] vin0_consume_en_2363;
  wire [0:0] vout_canPeek_2363;
  wire [7:0] vout_peek_2363;
  wire [0:0] v_2364;
  function [0:0] mux_2364(input [0:0] sel);
    case (sel) 0: mux_2364 = 1'h0; 1: mux_2364 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2365;
  wire [0:0] v_2366;
  wire [0:0] v_2367;
  function [0:0] mux_2367(input [0:0] sel);
    case (sel) 0: mux_2367 = 1'h0; 1: mux_2367 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2368;
  wire [0:0] vin0_consume_en_2369;
  wire [0:0] vout_canPeek_2369;
  wire [7:0] vout_peek_2369;
  wire [0:0] v_2370;
  function [0:0] mux_2370(input [0:0] sel);
    case (sel) 0: mux_2370 = 1'h0; 1: mux_2370 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2371;
  wire [0:0] v_2372;
  wire [0:0] v_2373;
  function [0:0] mux_2373(input [0:0] sel);
    case (sel) 0: mux_2373 = 1'h0; 1: mux_2373 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2374;
  wire [0:0] v_2375;
  wire [0:0] v_2376;
  wire [0:0] vin0_consume_en_2377;
  wire [0:0] vout_canPeek_2377;
  wire [7:0] vout_peek_2377;
  wire [0:0] v_2378;
  function [0:0] mux_2378(input [0:0] sel);
    case (sel) 0: mux_2378 = 1'h0; 1: mux_2378 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2379;
  wire [0:0] v_2380;
  wire [0:0] v_2381;
  function [0:0] mux_2381(input [0:0] sel);
    case (sel) 0: mux_2381 = 1'h0; 1: mux_2381 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2382;
  wire [0:0] vin0_consume_en_2383;
  wire [0:0] vout_canPeek_2383;
  wire [7:0] vout_peek_2383;
  wire [0:0] v_2384;
  function [0:0] mux_2384(input [0:0] sel);
    case (sel) 0: mux_2384 = 1'h0; 1: mux_2384 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2385;
  wire [0:0] v_2386;
  wire [0:0] v_2387;
  function [0:0] mux_2387(input [0:0] sel);
    case (sel) 0: mux_2387 = 1'h0; 1: mux_2387 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2388;
  wire [0:0] v_2389;
  wire [0:0] v_2390;
  wire [0:0] vin0_consume_en_2391;
  wire [0:0] vout_canPeek_2391;
  wire [7:0] vout_peek_2391;
  wire [0:0] v_2392;
  function [0:0] mux_2392(input [0:0] sel);
    case (sel) 0: mux_2392 = 1'h0; 1: mux_2392 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2393;
  wire [0:0] v_2394;
  wire [0:0] v_2395;
  function [0:0] mux_2395(input [0:0] sel);
    case (sel) 0: mux_2395 = 1'h0; 1: mux_2395 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2396;
  wire [0:0] vin0_consume_en_2397;
  wire [0:0] vout_canPeek_2397;
  wire [7:0] vout_peek_2397;
  wire [0:0] v_2398;
  function [0:0] mux_2398(input [0:0] sel);
    case (sel) 0: mux_2398 = 1'h0; 1: mux_2398 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2399;
  wire [0:0] v_2400;
  wire [0:0] v_2401;
  function [0:0] mux_2401(input [0:0] sel);
    case (sel) 0: mux_2401 = 1'h0; 1: mux_2401 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2402;
  wire [0:0] v_2403;
  wire [0:0] v_2404;
  wire [0:0] vin0_consume_en_2405;
  wire [0:0] vout_canPeek_2405;
  wire [7:0] vout_peek_2405;
  wire [0:0] v_2406;
  function [0:0] mux_2406(input [0:0] sel);
    case (sel) 0: mux_2406 = 1'h0; 1: mux_2406 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2407;
  wire [0:0] v_2408;
  wire [0:0] v_2409;
  function [0:0] mux_2409(input [0:0] sel);
    case (sel) 0: mux_2409 = 1'h0; 1: mux_2409 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2410;
  wire [0:0] vin0_consume_en_2411;
  wire [0:0] vout_canPeek_2411;
  wire [7:0] vout_peek_2411;
  wire [0:0] v_2412;
  function [0:0] mux_2412(input [0:0] sel);
    case (sel) 0: mux_2412 = 1'h0; 1: mux_2412 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2413;
  wire [0:0] v_2414;
  wire [0:0] v_2415;
  function [0:0] mux_2415(input [0:0] sel);
    case (sel) 0: mux_2415 = 1'h0; 1: mux_2415 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2416;
  wire [0:0] v_2417;
  wire [0:0] v_2418;
  wire [0:0] vin0_consume_en_2419;
  wire [0:0] vout_canPeek_2419;
  wire [7:0] vout_peek_2419;
  wire [0:0] v_2420;
  function [0:0] mux_2420(input [0:0] sel);
    case (sel) 0: mux_2420 = 1'h0; 1: mux_2420 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2421;
  wire [0:0] v_2422;
  wire [0:0] v_2423;
  function [0:0] mux_2423(input [0:0] sel);
    case (sel) 0: mux_2423 = 1'h0; 1: mux_2423 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2424;
  wire [0:0] vin0_consume_en_2425;
  wire [0:0] vout_canPeek_2425;
  wire [7:0] vout_peek_2425;
  wire [0:0] v_2426;
  function [0:0] mux_2426(input [0:0] sel);
    case (sel) 0: mux_2426 = 1'h0; 1: mux_2426 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2427;
  wire [0:0] v_2428;
  wire [0:0] v_2429;
  function [0:0] mux_2429(input [0:0] sel);
    case (sel) 0: mux_2429 = 1'h0; 1: mux_2429 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2430;
  wire [0:0] v_2431;
  wire [0:0] v_2432;
  wire [0:0] vin0_consume_en_2433;
  wire [0:0] vout_canPeek_2433;
  wire [7:0] vout_peek_2433;
  wire [0:0] v_2434;
  function [0:0] mux_2434(input [0:0] sel);
    case (sel) 0: mux_2434 = 1'h0; 1: mux_2434 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2435;
  wire [0:0] v_2436;
  wire [0:0] v_2437;
  function [0:0] mux_2437(input [0:0] sel);
    case (sel) 0: mux_2437 = 1'h0; 1: mux_2437 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2438;
  wire [0:0] vin0_consume_en_2439;
  wire [0:0] vout_canPeek_2439;
  wire [7:0] vout_peek_2439;
  wire [0:0] v_2440;
  function [0:0] mux_2440(input [0:0] sel);
    case (sel) 0: mux_2440 = 1'h0; 1: mux_2440 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2441;
  wire [0:0] v_2442;
  wire [0:0] v_2443;
  function [0:0] mux_2443(input [0:0] sel);
    case (sel) 0: mux_2443 = 1'h0; 1: mux_2443 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2444;
  wire [0:0] v_2445;
  wire [0:0] v_2446;
  wire [0:0] vin0_consume_en_2447;
  wire [0:0] vout_canPeek_2447;
  wire [7:0] vout_peek_2447;
  wire [0:0] v_2448;
  function [0:0] mux_2448(input [0:0] sel);
    case (sel) 0: mux_2448 = 1'h0; 1: mux_2448 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2449;
  wire [0:0] v_2450;
  wire [0:0] v_2451;
  function [0:0] mux_2451(input [0:0] sel);
    case (sel) 0: mux_2451 = 1'h0; 1: mux_2451 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2452;
  wire [0:0] vin0_consume_en_2453;
  wire [0:0] vout_canPeek_2453;
  wire [7:0] vout_peek_2453;
  wire [0:0] v_2454;
  function [0:0] mux_2454(input [0:0] sel);
    case (sel) 0: mux_2454 = 1'h0; 1: mux_2454 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2455;
  wire [0:0] v_2456;
  wire [0:0] v_2457;
  function [0:0] mux_2457(input [0:0] sel);
    case (sel) 0: mux_2457 = 1'h0; 1: mux_2457 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2458;
  wire [0:0] v_2459;
  wire [0:0] v_2460;
  wire [0:0] vin0_consume_en_2461;
  wire [0:0] vout_canPeek_2461;
  wire [7:0] vout_peek_2461;
  wire [0:0] v_2462;
  function [0:0] mux_2462(input [0:0] sel);
    case (sel) 0: mux_2462 = 1'h0; 1: mux_2462 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2463;
  wire [0:0] v_2464;
  wire [0:0] v_2465;
  function [0:0] mux_2465(input [0:0] sel);
    case (sel) 0: mux_2465 = 1'h0; 1: mux_2465 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2466;
  wire [0:0] vin0_consume_en_2467;
  wire [0:0] vout_canPeek_2467;
  wire [7:0] vout_peek_2467;
  wire [0:0] v_2468;
  function [0:0] mux_2468(input [0:0] sel);
    case (sel) 0: mux_2468 = 1'h0; 1: mux_2468 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2469;
  wire [0:0] v_2470;
  wire [0:0] v_2471;
  function [0:0] mux_2471(input [0:0] sel);
    case (sel) 0: mux_2471 = 1'h0; 1: mux_2471 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2472;
  wire [0:0] v_2473;
  wire [0:0] v_2474;
  wire [0:0] vin0_consume_en_2475;
  wire [0:0] vout_canPeek_2475;
  wire [7:0] vout_peek_2475;
  wire [0:0] v_2476;
  function [0:0] mux_2476(input [0:0] sel);
    case (sel) 0: mux_2476 = 1'h0; 1: mux_2476 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2477;
  wire [0:0] v_2478;
  wire [0:0] v_2479;
  function [0:0] mux_2479(input [0:0] sel);
    case (sel) 0: mux_2479 = 1'h0; 1: mux_2479 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2480;
  wire [0:0] vin0_consume_en_2481;
  wire [0:0] vout_canPeek_2481;
  wire [7:0] vout_peek_2481;
  wire [0:0] v_2482;
  function [0:0] mux_2482(input [0:0] sel);
    case (sel) 0: mux_2482 = 1'h0; 1: mux_2482 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2483;
  wire [0:0] v_2484;
  wire [0:0] v_2485;
  function [0:0] mux_2485(input [0:0] sel);
    case (sel) 0: mux_2485 = 1'h0; 1: mux_2485 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2486;
  wire [0:0] v_2487;
  wire [0:0] v_2488;
  wire [0:0] vin0_consume_en_2489;
  wire [0:0] vout_canPeek_2489;
  wire [7:0] vout_peek_2489;
  wire [0:0] v_2490;
  function [0:0] mux_2490(input [0:0] sel);
    case (sel) 0: mux_2490 = 1'h0; 1: mux_2490 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2491;
  wire [0:0] v_2492;
  wire [0:0] v_2493;
  function [0:0] mux_2493(input [0:0] sel);
    case (sel) 0: mux_2493 = 1'h0; 1: mux_2493 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2494;
  wire [0:0] vin0_consume_en_2495;
  wire [0:0] vout_canPeek_2495;
  wire [7:0] vout_peek_2495;
  wire [0:0] v_2496;
  function [0:0] mux_2496(input [0:0] sel);
    case (sel) 0: mux_2496 = 1'h0; 1: mux_2496 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2497;
  wire [0:0] v_2498;
  wire [0:0] v_2499;
  function [0:0] mux_2499(input [0:0] sel);
    case (sel) 0: mux_2499 = 1'h0; 1: mux_2499 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2500;
  wire [0:0] v_2501;
  wire [0:0] v_2502;
  wire [0:0] vin0_consume_en_2503;
  wire [0:0] vout_canPeek_2503;
  wire [7:0] vout_peek_2503;
  wire [0:0] v_2504;
  function [0:0] mux_2504(input [0:0] sel);
    case (sel) 0: mux_2504 = 1'h0; 1: mux_2504 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2505;
  wire [0:0] v_2506;
  wire [0:0] v_2507;
  function [0:0] mux_2507(input [0:0] sel);
    case (sel) 0: mux_2507 = 1'h0; 1: mux_2507 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2508;
  wire [0:0] vin0_consume_en_2509;
  wire [0:0] vout_canPeek_2509;
  wire [7:0] vout_peek_2509;
  wire [0:0] v_2510;
  function [0:0] mux_2510(input [0:0] sel);
    case (sel) 0: mux_2510 = 1'h0; 1: mux_2510 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2511;
  wire [0:0] v_2512;
  wire [0:0] v_2513;
  function [0:0] mux_2513(input [0:0] sel);
    case (sel) 0: mux_2513 = 1'h0; 1: mux_2513 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2514;
  wire [0:0] v_2515;
  wire [0:0] v_2516;
  wire [0:0] vin0_consume_en_2517;
  wire [0:0] vout_canPeek_2517;
  wire [7:0] vout_peek_2517;
  wire [0:0] v_2518;
  function [0:0] mux_2518(input [0:0] sel);
    case (sel) 0: mux_2518 = 1'h0; 1: mux_2518 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2519;
  wire [0:0] v_2520;
  wire [0:0] v_2521;
  function [0:0] mux_2521(input [0:0] sel);
    case (sel) 0: mux_2521 = 1'h0; 1: mux_2521 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2522;
  wire [0:0] vin0_consume_en_2523;
  wire [0:0] vout_canPeek_2523;
  wire [7:0] vout_peek_2523;
  wire [0:0] v_2524;
  function [0:0] mux_2524(input [0:0] sel);
    case (sel) 0: mux_2524 = 1'h0; 1: mux_2524 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2525;
  wire [0:0] v_2526;
  wire [0:0] v_2527;
  function [0:0] mux_2527(input [0:0] sel);
    case (sel) 0: mux_2527 = 1'h0; 1: mux_2527 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2528;
  wire [0:0] v_2529;
  wire [0:0] v_2530;
  wire [0:0] vin0_consume_en_2531;
  wire [0:0] vout_canPeek_2531;
  wire [7:0] vout_peek_2531;
  wire [0:0] v_2532;
  function [0:0] mux_2532(input [0:0] sel);
    case (sel) 0: mux_2532 = 1'h0; 1: mux_2532 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2533;
  wire [0:0] v_2534;
  wire [0:0] v_2535;
  function [0:0] mux_2535(input [0:0] sel);
    case (sel) 0: mux_2535 = 1'h0; 1: mux_2535 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2536;
  wire [0:0] vin0_consume_en_2537;
  wire [0:0] vout_canPeek_2537;
  wire [7:0] vout_peek_2537;
  wire [0:0] v_2538;
  function [0:0] mux_2538(input [0:0] sel);
    case (sel) 0: mux_2538 = 1'h0; 1: mux_2538 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2539;
  wire [0:0] v_2540;
  wire [0:0] v_2541;
  function [0:0] mux_2541(input [0:0] sel);
    case (sel) 0: mux_2541 = 1'h0; 1: mux_2541 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2542;
  wire [0:0] v_2543;
  wire [0:0] v_2544;
  wire [0:0] vin0_consume_en_2545;
  wire [0:0] vout_canPeek_2545;
  wire [7:0] vout_peek_2545;
  wire [0:0] v_2546;
  function [0:0] mux_2546(input [0:0] sel);
    case (sel) 0: mux_2546 = 1'h0; 1: mux_2546 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2547;
  wire [0:0] v_2548;
  wire [0:0] v_2549;
  function [0:0] mux_2549(input [0:0] sel);
    case (sel) 0: mux_2549 = 1'h0; 1: mux_2549 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2550;
  wire [0:0] vin0_consume_en_2551;
  wire [0:0] vout_canPeek_2551;
  wire [7:0] vout_peek_2551;
  wire [0:0] v_2552;
  function [0:0] mux_2552(input [0:0] sel);
    case (sel) 0: mux_2552 = 1'h0; 1: mux_2552 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2553;
  wire [0:0] v_2554;
  wire [0:0] v_2555;
  function [0:0] mux_2555(input [0:0] sel);
    case (sel) 0: mux_2555 = 1'h0; 1: mux_2555 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2556;
  wire [0:0] v_2557;
  wire [0:0] v_2558;
  wire [0:0] vin0_consume_en_2559;
  wire [0:0] vout_canPeek_2559;
  wire [7:0] vout_peek_2559;
  wire [0:0] v_2560;
  function [0:0] mux_2560(input [0:0] sel);
    case (sel) 0: mux_2560 = 1'h0; 1: mux_2560 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2561;
  wire [0:0] v_2562;
  wire [0:0] v_2563;
  function [0:0] mux_2563(input [0:0] sel);
    case (sel) 0: mux_2563 = 1'h0; 1: mux_2563 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2564;
  wire [0:0] vin0_consume_en_2565;
  wire [0:0] vout_canPeek_2565;
  wire [7:0] vout_peek_2565;
  wire [0:0] v_2566;
  function [0:0] mux_2566(input [0:0] sel);
    case (sel) 0: mux_2566 = 1'h0; 1: mux_2566 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2567;
  wire [0:0] v_2568;
  wire [0:0] v_2569;
  function [0:0] mux_2569(input [0:0] sel);
    case (sel) 0: mux_2569 = 1'h0; 1: mux_2569 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2570;
  wire [0:0] v_2571;
  wire [0:0] v_2572;
  wire [0:0] vin0_consume_en_2573;
  wire [0:0] vout_canPeek_2573;
  wire [7:0] vout_peek_2573;
  wire [0:0] v_2574;
  function [0:0] mux_2574(input [0:0] sel);
    case (sel) 0: mux_2574 = 1'h0; 1: mux_2574 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2575;
  wire [0:0] v_2576;
  wire [0:0] v_2577;
  function [0:0] mux_2577(input [0:0] sel);
    case (sel) 0: mux_2577 = 1'h0; 1: mux_2577 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2578;
  wire [0:0] vin0_consume_en_2579;
  wire [0:0] vout_canPeek_2579;
  wire [7:0] vout_peek_2579;
  wire [0:0] v_2580;
  function [0:0] mux_2580(input [0:0] sel);
    case (sel) 0: mux_2580 = 1'h0; 1: mux_2580 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2581;
  wire [0:0] v_2582;
  wire [0:0] v_2583;
  function [0:0] mux_2583(input [0:0] sel);
    case (sel) 0: mux_2583 = 1'h0; 1: mux_2583 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2584;
  wire [0:0] v_2585;
  wire [0:0] v_2586;
  wire [0:0] vin0_consume_en_2587;
  wire [0:0] vout_canPeek_2587;
  wire [7:0] vout_peek_2587;
  wire [0:0] v_2588;
  function [0:0] mux_2588(input [0:0] sel);
    case (sel) 0: mux_2588 = 1'h0; 1: mux_2588 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2589;
  wire [0:0] v_2590;
  wire [0:0] v_2591;
  function [0:0] mux_2591(input [0:0] sel);
    case (sel) 0: mux_2591 = 1'h0; 1: mux_2591 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2592;
  wire [0:0] vin0_consume_en_2593;
  wire [0:0] vout_canPeek_2593;
  wire [7:0] vout_peek_2593;
  wire [0:0] v_2594;
  function [0:0] mux_2594(input [0:0] sel);
    case (sel) 0: mux_2594 = 1'h0; 1: mux_2594 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2595;
  wire [0:0] v_2596;
  wire [0:0] v_2597;
  function [0:0] mux_2597(input [0:0] sel);
    case (sel) 0: mux_2597 = 1'h0; 1: mux_2597 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2598;
  wire [0:0] v_2599;
  wire [0:0] v_2600;
  wire [0:0] vin0_consume_en_2601;
  wire [0:0] vout_canPeek_2601;
  wire [7:0] vout_peek_2601;
  wire [0:0] v_2602;
  function [0:0] mux_2602(input [0:0] sel);
    case (sel) 0: mux_2602 = 1'h0; 1: mux_2602 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2603;
  wire [0:0] v_2604;
  wire [0:0] v_2605;
  function [0:0] mux_2605(input [0:0] sel);
    case (sel) 0: mux_2605 = 1'h0; 1: mux_2605 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2606;
  wire [0:0] vin0_consume_en_2607;
  wire [0:0] vout_canPeek_2607;
  wire [7:0] vout_peek_2607;
  wire [0:0] v_2608;
  function [0:0] mux_2608(input [0:0] sel);
    case (sel) 0: mux_2608 = 1'h0; 1: mux_2608 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2609;
  wire [0:0] v_2610;
  wire [0:0] v_2611;
  function [0:0] mux_2611(input [0:0] sel);
    case (sel) 0: mux_2611 = 1'h0; 1: mux_2611 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2612;
  wire [0:0] v_2613;
  wire [0:0] v_2614;
  wire [0:0] vin0_consume_en_2615;
  wire [0:0] vout_canPeek_2615;
  wire [7:0] vout_peek_2615;
  wire [0:0] v_2616;
  function [0:0] mux_2616(input [0:0] sel);
    case (sel) 0: mux_2616 = 1'h0; 1: mux_2616 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2617;
  wire [0:0] v_2618;
  wire [0:0] v_2619;
  function [0:0] mux_2619(input [0:0] sel);
    case (sel) 0: mux_2619 = 1'h0; 1: mux_2619 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2620;
  wire [0:0] vin0_consume_en_2621;
  wire [0:0] vout_canPeek_2621;
  wire [7:0] vout_peek_2621;
  wire [0:0] v_2622;
  function [0:0] mux_2622(input [0:0] sel);
    case (sel) 0: mux_2622 = 1'h0; 1: mux_2622 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2623;
  wire [0:0] v_2624;
  wire [0:0] v_2625;
  function [0:0] mux_2625(input [0:0] sel);
    case (sel) 0: mux_2625 = 1'h0; 1: mux_2625 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2626;
  wire [0:0] v_2627;
  wire [0:0] v_2628;
  wire [0:0] vin0_consume_en_2629;
  wire [0:0] vout_canPeek_2629;
  wire [7:0] vout_peek_2629;
  wire [0:0] v_2630;
  function [0:0] mux_2630(input [0:0] sel);
    case (sel) 0: mux_2630 = 1'h0; 1: mux_2630 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2631;
  wire [0:0] v_2632;
  wire [0:0] v_2633;
  function [0:0] mux_2633(input [0:0] sel);
    case (sel) 0: mux_2633 = 1'h0; 1: mux_2633 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2634;
  wire [0:0] vin0_consume_en_2635;
  wire [0:0] vout_canPeek_2635;
  wire [7:0] vout_peek_2635;
  wire [0:0] v_2636;
  function [0:0] mux_2636(input [0:0] sel);
    case (sel) 0: mux_2636 = 1'h0; 1: mux_2636 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2637;
  wire [0:0] v_2638;
  wire [0:0] v_2639;
  function [0:0] mux_2639(input [0:0] sel);
    case (sel) 0: mux_2639 = 1'h0; 1: mux_2639 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2640;
  wire [0:0] v_2641;
  wire [0:0] v_2642;
  wire [0:0] vin0_consume_en_2643;
  wire [0:0] vout_canPeek_2643;
  wire [7:0] vout_peek_2643;
  wire [0:0] v_2644;
  function [0:0] mux_2644(input [0:0] sel);
    case (sel) 0: mux_2644 = 1'h0; 1: mux_2644 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2645;
  wire [0:0] v_2646;
  wire [0:0] v_2647;
  function [0:0] mux_2647(input [0:0] sel);
    case (sel) 0: mux_2647 = 1'h0; 1: mux_2647 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2648;
  wire [0:0] vin0_consume_en_2649;
  wire [0:0] vout_canPeek_2649;
  wire [7:0] vout_peek_2649;
  wire [0:0] v_2650;
  function [0:0] mux_2650(input [0:0] sel);
    case (sel) 0: mux_2650 = 1'h0; 1: mux_2650 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2651;
  wire [0:0] v_2652;
  wire [0:0] v_2653;
  function [0:0] mux_2653(input [0:0] sel);
    case (sel) 0: mux_2653 = 1'h0; 1: mux_2653 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2654;
  wire [0:0] v_2655;
  wire [0:0] v_2656;
  wire [0:0] vin0_consume_en_2657;
  wire [0:0] vout_canPeek_2657;
  wire [7:0] vout_peek_2657;
  wire [0:0] v_2658;
  function [0:0] mux_2658(input [0:0] sel);
    case (sel) 0: mux_2658 = 1'h0; 1: mux_2658 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2659;
  wire [0:0] v_2660;
  wire [0:0] v_2661;
  function [0:0] mux_2661(input [0:0] sel);
    case (sel) 0: mux_2661 = 1'h0; 1: mux_2661 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2662;
  wire [0:0] vin0_consume_en_2663;
  wire [0:0] vout_canPeek_2663;
  wire [7:0] vout_peek_2663;
  wire [0:0] v_2664;
  function [0:0] mux_2664(input [0:0] sel);
    case (sel) 0: mux_2664 = 1'h0; 1: mux_2664 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2665;
  wire [0:0] v_2666;
  wire [0:0] v_2667;
  function [0:0] mux_2667(input [0:0] sel);
    case (sel) 0: mux_2667 = 1'h0; 1: mux_2667 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2668;
  wire [0:0] v_2669;
  wire [0:0] v_2670;
  wire [0:0] vin0_consume_en_2671;
  wire [0:0] vout_canPeek_2671;
  wire [7:0] vout_peek_2671;
  wire [0:0] v_2672;
  function [0:0] mux_2672(input [0:0] sel);
    case (sel) 0: mux_2672 = 1'h0; 1: mux_2672 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2673;
  wire [0:0] v_2674;
  wire [0:0] v_2675;
  function [0:0] mux_2675(input [0:0] sel);
    case (sel) 0: mux_2675 = 1'h0; 1: mux_2675 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2676;
  wire [0:0] vin0_consume_en_2677;
  wire [0:0] vout_canPeek_2677;
  wire [7:0] vout_peek_2677;
  wire [0:0] v_2678;
  function [0:0] mux_2678(input [0:0] sel);
    case (sel) 0: mux_2678 = 1'h0; 1: mux_2678 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2679;
  wire [0:0] v_2680;
  wire [0:0] v_2681;
  function [0:0] mux_2681(input [0:0] sel);
    case (sel) 0: mux_2681 = 1'h0; 1: mux_2681 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2682;
  wire [0:0] v_2683;
  wire [0:0] v_2684;
  wire [0:0] vin0_consume_en_2685;
  wire [0:0] vout_canPeek_2685;
  wire [7:0] vout_peek_2685;
  wire [0:0] v_2686;
  function [0:0] mux_2686(input [0:0] sel);
    case (sel) 0: mux_2686 = 1'h0; 1: mux_2686 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2687;
  wire [0:0] v_2688;
  wire [0:0] v_2689;
  function [0:0] mux_2689(input [0:0] sel);
    case (sel) 0: mux_2689 = 1'h0; 1: mux_2689 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2690;
  wire [0:0] vin0_consume_en_2691;
  wire [0:0] vout_canPeek_2691;
  wire [7:0] vout_peek_2691;
  wire [0:0] v_2692;
  function [0:0] mux_2692(input [0:0] sel);
    case (sel) 0: mux_2692 = 1'h0; 1: mux_2692 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2693;
  wire [0:0] v_2694;
  wire [0:0] v_2695;
  function [0:0] mux_2695(input [0:0] sel);
    case (sel) 0: mux_2695 = 1'h0; 1: mux_2695 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2696;
  wire [0:0] v_2697;
  wire [0:0] v_2698;
  wire [0:0] vin0_consume_en_2699;
  wire [0:0] vout_canPeek_2699;
  wire [7:0] vout_peek_2699;
  wire [0:0] v_2700;
  function [0:0] mux_2700(input [0:0] sel);
    case (sel) 0: mux_2700 = 1'h0; 1: mux_2700 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2701;
  wire [0:0] v_2702;
  wire [0:0] v_2703;
  function [0:0] mux_2703(input [0:0] sel);
    case (sel) 0: mux_2703 = 1'h0; 1: mux_2703 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2704;
  wire [0:0] vin0_consume_en_2705;
  wire [0:0] vout_canPeek_2705;
  wire [7:0] vout_peek_2705;
  wire [0:0] v_2706;
  function [0:0] mux_2706(input [0:0] sel);
    case (sel) 0: mux_2706 = 1'h0; 1: mux_2706 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2707;
  wire [0:0] v_2708;
  wire [0:0] v_2709;
  function [0:0] mux_2709(input [0:0] sel);
    case (sel) 0: mux_2709 = 1'h0; 1: mux_2709 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2710;
  wire [0:0] v_2711;
  wire [0:0] v_2712;
  wire [0:0] vin0_consume_en_2713;
  wire [0:0] vout_canPeek_2713;
  wire [7:0] vout_peek_2713;
  wire [0:0] v_2714;
  function [0:0] mux_2714(input [0:0] sel);
    case (sel) 0: mux_2714 = 1'h0; 1: mux_2714 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2715;
  wire [0:0] v_2716;
  wire [0:0] v_2717;
  function [0:0] mux_2717(input [0:0] sel);
    case (sel) 0: mux_2717 = 1'h0; 1: mux_2717 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2718;
  wire [0:0] vin0_consume_en_2719;
  wire [0:0] vout_canPeek_2719;
  wire [7:0] vout_peek_2719;
  wire [0:0] v_2720;
  function [0:0] mux_2720(input [0:0] sel);
    case (sel) 0: mux_2720 = 1'h0; 1: mux_2720 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2721;
  wire [0:0] v_2722;
  wire [0:0] v_2723;
  function [0:0] mux_2723(input [0:0] sel);
    case (sel) 0: mux_2723 = 1'h0; 1: mux_2723 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2724;
  wire [0:0] v_2725;
  wire [0:0] v_2726;
  wire [0:0] vin0_consume_en_2727;
  wire [0:0] vout_canPeek_2727;
  wire [7:0] vout_peek_2727;
  wire [0:0] v_2728;
  function [0:0] mux_2728(input [0:0] sel);
    case (sel) 0: mux_2728 = 1'h0; 1: mux_2728 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2729;
  wire [0:0] v_2730;
  wire [0:0] v_2731;
  function [0:0] mux_2731(input [0:0] sel);
    case (sel) 0: mux_2731 = 1'h0; 1: mux_2731 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2732;
  wire [0:0] vin0_consume_en_2733;
  wire [0:0] vout_canPeek_2733;
  wire [7:0] vout_peek_2733;
  wire [0:0] v_2734;
  function [0:0] mux_2734(input [0:0] sel);
    case (sel) 0: mux_2734 = 1'h0; 1: mux_2734 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2735;
  wire [0:0] v_2736;
  wire [0:0] v_2737;
  function [0:0] mux_2737(input [0:0] sel);
    case (sel) 0: mux_2737 = 1'h0; 1: mux_2737 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2738;
  wire [0:0] v_2739;
  wire [0:0] v_2740;
  wire [0:0] vin0_consume_en_2741;
  wire [0:0] vout_canPeek_2741;
  wire [7:0] vout_peek_2741;
  wire [0:0] v_2742;
  function [0:0] mux_2742(input [0:0] sel);
    case (sel) 0: mux_2742 = 1'h0; 1: mux_2742 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2743;
  wire [0:0] v_2744;
  wire [0:0] v_2745;
  function [0:0] mux_2745(input [0:0] sel);
    case (sel) 0: mux_2745 = 1'h0; 1: mux_2745 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2746;
  wire [0:0] vin0_consume_en_2747;
  wire [0:0] vout_canPeek_2747;
  wire [7:0] vout_peek_2747;
  wire [0:0] v_2748;
  function [0:0] mux_2748(input [0:0] sel);
    case (sel) 0: mux_2748 = 1'h0; 1: mux_2748 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2749;
  wire [0:0] v_2750;
  wire [0:0] v_2751;
  function [0:0] mux_2751(input [0:0] sel);
    case (sel) 0: mux_2751 = 1'h0; 1: mux_2751 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2752;
  wire [0:0] v_2753;
  wire [0:0] v_2754;
  wire [0:0] vin0_consume_en_2755;
  wire [0:0] vout_canPeek_2755;
  wire [7:0] vout_peek_2755;
  wire [0:0] v_2756;
  function [0:0] mux_2756(input [0:0] sel);
    case (sel) 0: mux_2756 = 1'h0; 1: mux_2756 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2757;
  wire [0:0] v_2758;
  wire [0:0] v_2759;
  function [0:0] mux_2759(input [0:0] sel);
    case (sel) 0: mux_2759 = 1'h0; 1: mux_2759 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2760;
  wire [0:0] vin0_consume_en_2761;
  wire [0:0] vout_canPeek_2761;
  wire [7:0] vout_peek_2761;
  wire [0:0] v_2762;
  function [0:0] mux_2762(input [0:0] sel);
    case (sel) 0: mux_2762 = 1'h0; 1: mux_2762 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2763;
  wire [0:0] v_2764;
  wire [0:0] v_2765;
  function [0:0] mux_2765(input [0:0] sel);
    case (sel) 0: mux_2765 = 1'h0; 1: mux_2765 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2766;
  wire [0:0] v_2767;
  wire [0:0] v_2768;
  wire [0:0] vin0_consume_en_2769;
  wire [0:0] vout_canPeek_2769;
  wire [7:0] vout_peek_2769;
  wire [0:0] v_2770;
  function [0:0] mux_2770(input [0:0] sel);
    case (sel) 0: mux_2770 = 1'h0; 1: mux_2770 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2771;
  wire [0:0] v_2772;
  wire [0:0] v_2773;
  function [0:0] mux_2773(input [0:0] sel);
    case (sel) 0: mux_2773 = 1'h0; 1: mux_2773 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2774;
  wire [0:0] vin0_consume_en_2775;
  wire [0:0] vout_canPeek_2775;
  wire [7:0] vout_peek_2775;
  wire [0:0] v_2776;
  function [0:0] mux_2776(input [0:0] sel);
    case (sel) 0: mux_2776 = 1'h0; 1: mux_2776 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2777;
  wire [0:0] v_2778;
  wire [0:0] v_2779;
  function [0:0] mux_2779(input [0:0] sel);
    case (sel) 0: mux_2779 = 1'h0; 1: mux_2779 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2780;
  wire [0:0] v_2781;
  wire [0:0] v_2782;
  wire [0:0] vin0_consume_en_2783;
  wire [0:0] vout_canPeek_2783;
  wire [7:0] vout_peek_2783;
  wire [0:0] v_2784;
  function [0:0] mux_2784(input [0:0] sel);
    case (sel) 0: mux_2784 = 1'h0; 1: mux_2784 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2785;
  wire [0:0] v_2786;
  wire [0:0] v_2787;
  function [0:0] mux_2787(input [0:0] sel);
    case (sel) 0: mux_2787 = 1'h0; 1: mux_2787 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2788;
  wire [0:0] vin0_consume_en_2789;
  wire [0:0] vout_canPeek_2789;
  wire [7:0] vout_peek_2789;
  wire [0:0] v_2790;
  function [0:0] mux_2790(input [0:0] sel);
    case (sel) 0: mux_2790 = 1'h0; 1: mux_2790 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2791;
  wire [0:0] v_2792;
  wire [0:0] v_2793;
  function [0:0] mux_2793(input [0:0] sel);
    case (sel) 0: mux_2793 = 1'h0; 1: mux_2793 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2794;
  wire [0:0] v_2795;
  wire [0:0] v_2796;
  wire [0:0] vin0_consume_en_2797;
  wire [0:0] vout_canPeek_2797;
  wire [7:0] vout_peek_2797;
  wire [0:0] v_2798;
  function [0:0] mux_2798(input [0:0] sel);
    case (sel) 0: mux_2798 = 1'h0; 1: mux_2798 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2799;
  wire [0:0] v_2801;
  function [0:0] mux_2801(input [0:0] sel);
    case (sel) 0: mux_2801 = 1'h0; 1: mux_2801 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2802;
  reg [0:0] v_2804 = 1'h0;
  wire [0:0] v_2805;
  wire [0:0] v_2806;
  wire [0:0] act_2807;
  wire [0:0] v_2808;
  wire [0:0] v_2809;
  wire [0:0] v_2810;
  reg [0:0] v_2811 = 1'h0;
  wire [0:0] v_2812;
  wire [0:0] v_2813;
  wire [0:0] act_2814;
  wire [0:0] v_2815;
  wire [0:0] v_2816;
  wire [0:0] v_2817;
  reg [0:0] v_2818 = 1'h0;
  wire [0:0] v_2819;
  wire [0:0] v_2820;
  wire [0:0] act_2821;
  wire [0:0] v_2822;
  wire [0:0] v_2823;
  wire [0:0] v_2824;
  reg [0:0] v_2825 = 1'h0;
  wire [0:0] v_2826;
  wire [0:0] v_2827;
  wire [0:0] act_2828;
  wire [0:0] v_2829;
  wire [0:0] v_2830;
  wire [0:0] v_2831;
  reg [0:0] v_2832 = 1'h0;
  wire [0:0] v_2833;
  wire [0:0] v_2834;
  wire [0:0] act_2835;
  wire [0:0] v_2836;
  wire [0:0] v_2837;
  wire [0:0] v_2838;
  reg [0:0] v_2839 = 1'h0;
  wire [0:0] v_2840;
  wire [0:0] v_2841;
  wire [0:0] act_2842;
  wire [0:0] v_2843;
  wire [0:0] v_2844;
  wire [0:0] v_2845;
  reg [0:0] v_2846 = 1'h0;
  wire [0:0] v_2847;
  wire [0:0] v_2848;
  wire [0:0] act_2849;
  wire [0:0] v_2850;
  wire [0:0] v_2851;
  wire [0:0] v_2852;
  reg [0:0] v_2853 = 1'h0;
  wire [0:0] v_2854;
  wire [0:0] v_2855;
  wire [0:0] act_2856;
  wire [0:0] v_2857;
  wire [0:0] v_2858;
  wire [0:0] v_2859;
  wire [0:0] v_2860;
  wire [0:0] v_2861;
  wire [0:0] v_2862;
  function [0:0] mux_2862(input [0:0] sel);
    case (sel) 0: mux_2862 = 1'h0; 1: mux_2862 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2863;
  wire [0:0] v_2864;
  function [0:0] mux_2864(input [0:0] sel);
    case (sel) 0: mux_2864 = 1'h0; 1: mux_2864 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2865;
  wire [0:0] v_2866;
  wire [0:0] v_2867;
  wire [0:0] v_2868;
  function [0:0] mux_2868(input [0:0] sel);
    case (sel) 0: mux_2868 = 1'h0; 1: mux_2868 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2869;
  function [0:0] mux_2869(input [0:0] sel);
    case (sel) 0: mux_2869 = 1'h0; 1: mux_2869 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2870 = 1'h0;
  wire [0:0] v_2871;
  wire [0:0] v_2872;
  wire [0:0] act_2873;
  wire [0:0] v_2874;
  wire [0:0] v_2875;
  wire [0:0] v_2876;
  wire [0:0] v_2877;
  wire [0:0] v_2878;
  wire [0:0] v_2879;
  function [0:0] mux_2879(input [0:0] sel);
    case (sel) 0: mux_2879 = 1'h0; 1: mux_2879 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2880;
  function [0:0] mux_2880(input [0:0] sel);
    case (sel) 0: mux_2880 = 1'h0; 1: mux_2880 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2881;
  wire [0:0] v_2882;
  wire [0:0] v_2883;
  wire [0:0] v_2884;
  function [0:0] mux_2884(input [0:0] sel);
    case (sel) 0: mux_2884 = 1'h0; 1: mux_2884 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2885;
  function [0:0] mux_2885(input [0:0] sel);
    case (sel) 0: mux_2885 = 1'h0; 1: mux_2885 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2886;
  wire [0:0] v_2887;
  wire [0:0] v_2888;
  wire [0:0] v_2889;
  wire [0:0] v_2890;
  wire [0:0] v_2891;
  function [0:0] mux_2891(input [0:0] sel);
    case (sel) 0: mux_2891 = 1'h0; 1: mux_2891 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2892;
  wire [0:0] v_2893;
  function [0:0] mux_2893(input [0:0] sel);
    case (sel) 0: mux_2893 = 1'h0; 1: mux_2893 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2894;
  wire [0:0] v_2895;
  wire [0:0] v_2896;
  wire [0:0] v_2897;
  function [0:0] mux_2897(input [0:0] sel);
    case (sel) 0: mux_2897 = 1'h0; 1: mux_2897 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2898;
  function [0:0] mux_2898(input [0:0] sel);
    case (sel) 0: mux_2898 = 1'h0; 1: mux_2898 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2899 = 1'h0;
  wire [0:0] v_2900;
  wire [0:0] v_2901;
  wire [0:0] act_2902;
  wire [0:0] v_2903;
  wire [0:0] v_2904;
  wire [0:0] v_2905;
  reg [0:0] v_2906 = 1'h0;
  wire [0:0] v_2907;
  wire [0:0] v_2908;
  wire [0:0] act_2909;
  wire [0:0] v_2910;
  wire [0:0] v_2911;
  wire [0:0] v_2912;
  wire [0:0] v_2913;
  wire [0:0] v_2914;
  wire [0:0] v_2915;
  function [0:0] mux_2915(input [0:0] sel);
    case (sel) 0: mux_2915 = 1'h0; 1: mux_2915 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2916;
  wire [0:0] v_2917;
  function [0:0] mux_2917(input [0:0] sel);
    case (sel) 0: mux_2917 = 1'h0; 1: mux_2917 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2918;
  wire [0:0] v_2919;
  wire [0:0] v_2920;
  wire [0:0] v_2921;
  function [0:0] mux_2921(input [0:0] sel);
    case (sel) 0: mux_2921 = 1'h0; 1: mux_2921 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2922;
  function [0:0] mux_2922(input [0:0] sel);
    case (sel) 0: mux_2922 = 1'h0; 1: mux_2922 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2923 = 1'h0;
  wire [0:0] v_2924;
  wire [0:0] v_2925;
  wire [0:0] act_2926;
  wire [0:0] v_2927;
  wire [0:0] v_2928;
  wire [0:0] v_2929;
  wire [0:0] v_2930;
  wire [0:0] v_2931;
  wire [0:0] v_2932;
  function [0:0] mux_2932(input [0:0] sel);
    case (sel) 0: mux_2932 = 1'h0; 1: mux_2932 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2933;
  function [0:0] mux_2933(input [0:0] sel);
    case (sel) 0: mux_2933 = 1'h0; 1: mux_2933 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2934;
  wire [0:0] v_2935;
  wire [0:0] v_2936;
  wire [0:0] v_2937;
  function [0:0] mux_2937(input [0:0] sel);
    case (sel) 0: mux_2937 = 1'h0; 1: mux_2937 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2938;
  function [0:0] mux_2938(input [0:0] sel);
    case (sel) 0: mux_2938 = 1'h0; 1: mux_2938 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2939;
  wire [0:0] v_2940;
  wire [0:0] v_2941;
  wire [0:0] v_2942;
  wire [0:0] v_2943;
  wire [0:0] v_2944;
  function [0:0] mux_2944(input [0:0] sel);
    case (sel) 0: mux_2944 = 1'h0; 1: mux_2944 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2945;
  function [0:0] mux_2945(input [0:0] sel);
    case (sel) 0: mux_2945 = 1'h0; 1: mux_2945 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2946;
  wire [0:0] v_2947;
  wire [0:0] v_2948;
  wire [0:0] v_2949;
  function [0:0] mux_2949(input [0:0] sel);
    case (sel) 0: mux_2949 = 1'h0; 1: mux_2949 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2950;
  function [0:0] mux_2950(input [0:0] sel);
    case (sel) 0: mux_2950 = 1'h0; 1: mux_2950 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2951;
  wire [0:0] v_2952;
  wire [0:0] v_2953;
  wire [0:0] v_2954;
  wire [0:0] v_2955;
  wire [0:0] v_2956;
  function [0:0] mux_2956(input [0:0] sel);
    case (sel) 0: mux_2956 = 1'h0; 1: mux_2956 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2957;
  wire [0:0] v_2958;
  function [0:0] mux_2958(input [0:0] sel);
    case (sel) 0: mux_2958 = 1'h0; 1: mux_2958 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2959;
  wire [0:0] v_2960;
  wire [0:0] v_2961;
  wire [0:0] v_2962;
  function [0:0] mux_2962(input [0:0] sel);
    case (sel) 0: mux_2962 = 1'h0; 1: mux_2962 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2963;
  function [0:0] mux_2963(input [0:0] sel);
    case (sel) 0: mux_2963 = 1'h0; 1: mux_2963 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2964 = 1'h0;
  wire [0:0] v_2965;
  wire [0:0] v_2966;
  wire [0:0] act_2967;
  wire [0:0] v_2968;
  wire [0:0] v_2969;
  wire [0:0] v_2970;
  reg [0:0] v_2971 = 1'h0;
  wire [0:0] v_2972;
  wire [0:0] v_2973;
  wire [0:0] act_2974;
  wire [0:0] v_2975;
  wire [0:0] v_2976;
  wire [0:0] v_2977;
  reg [0:0] v_2978 = 1'h0;
  wire [0:0] v_2979;
  wire [0:0] v_2980;
  wire [0:0] act_2981;
  wire [0:0] v_2982;
  wire [0:0] v_2983;
  wire [0:0] v_2984;
  wire [0:0] v_2985;
  wire [0:0] v_2986;
  wire [0:0] v_2987;
  function [0:0] mux_2987(input [0:0] sel);
    case (sel) 0: mux_2987 = 1'h0; 1: mux_2987 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2988;
  wire [0:0] v_2989;
  function [0:0] mux_2989(input [0:0] sel);
    case (sel) 0: mux_2989 = 1'h0; 1: mux_2989 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_2990;
  wire [0:0] v_2991;
  wire [0:0] v_2992;
  wire [0:0] v_2993;
  function [0:0] mux_2993(input [0:0] sel);
    case (sel) 0: mux_2993 = 1'h0; 1: mux_2993 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_2994;
  function [0:0] mux_2994(input [0:0] sel);
    case (sel) 0: mux_2994 = 1'h0; 1: mux_2994 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_2995 = 1'h0;
  wire [0:0] v_2996;
  wire [0:0] v_2997;
  wire [0:0] act_2998;
  wire [0:0] v_2999;
  wire [0:0] v_3000;
  wire [0:0] v_3001;
  wire [0:0] v_3002;
  wire [0:0] v_3003;
  wire [0:0] v_3004;
  function [0:0] mux_3004(input [0:0] sel);
    case (sel) 0: mux_3004 = 1'h0; 1: mux_3004 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3005;
  function [0:0] mux_3005(input [0:0] sel);
    case (sel) 0: mux_3005 = 1'h0; 1: mux_3005 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3006;
  wire [0:0] v_3007;
  wire [0:0] v_3008;
  wire [0:0] v_3009;
  function [0:0] mux_3009(input [0:0] sel);
    case (sel) 0: mux_3009 = 1'h0; 1: mux_3009 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3010;
  function [0:0] mux_3010(input [0:0] sel);
    case (sel) 0: mux_3010 = 1'h0; 1: mux_3010 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3011;
  wire [0:0] v_3012;
  wire [0:0] v_3013;
  wire [0:0] v_3014;
  wire [0:0] v_3015;
  wire [0:0] v_3016;
  function [0:0] mux_3016(input [0:0] sel);
    case (sel) 0: mux_3016 = 1'h0; 1: mux_3016 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3017;
  wire [0:0] v_3018;
  function [0:0] mux_3018(input [0:0] sel);
    case (sel) 0: mux_3018 = 1'h0; 1: mux_3018 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3019;
  wire [0:0] v_3020;
  wire [0:0] v_3021;
  wire [0:0] v_3022;
  function [0:0] mux_3022(input [0:0] sel);
    case (sel) 0: mux_3022 = 1'h0; 1: mux_3022 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3023;
  function [0:0] mux_3023(input [0:0] sel);
    case (sel) 0: mux_3023 = 1'h0; 1: mux_3023 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3024 = 1'h0;
  wire [0:0] v_3025;
  wire [0:0] v_3026;
  wire [0:0] act_3027;
  wire [0:0] v_3028;
  wire [0:0] v_3029;
  wire [0:0] v_3030;
  reg [0:0] v_3031 = 1'h0;
  wire [0:0] v_3032;
  wire [0:0] v_3033;
  wire [0:0] act_3034;
  wire [0:0] v_3035;
  wire [0:0] v_3036;
  wire [0:0] v_3037;
  wire [0:0] v_3038;
  wire [0:0] v_3039;
  wire [0:0] v_3040;
  function [0:0] mux_3040(input [0:0] sel);
    case (sel) 0: mux_3040 = 1'h0; 1: mux_3040 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3041;
  wire [0:0] v_3042;
  function [0:0] mux_3042(input [0:0] sel);
    case (sel) 0: mux_3042 = 1'h0; 1: mux_3042 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3043;
  wire [0:0] v_3044;
  wire [0:0] v_3045;
  wire [0:0] v_3046;
  function [0:0] mux_3046(input [0:0] sel);
    case (sel) 0: mux_3046 = 1'h0; 1: mux_3046 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3047;
  function [0:0] mux_3047(input [0:0] sel);
    case (sel) 0: mux_3047 = 1'h0; 1: mux_3047 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3048 = 1'h0;
  wire [0:0] v_3049;
  wire [0:0] v_3050;
  wire [0:0] act_3051;
  wire [0:0] v_3052;
  wire [0:0] v_3053;
  wire [0:0] v_3054;
  wire [0:0] v_3055;
  wire [0:0] v_3056;
  wire [0:0] v_3057;
  function [0:0] mux_3057(input [0:0] sel);
    case (sel) 0: mux_3057 = 1'h0; 1: mux_3057 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3058;
  function [0:0] mux_3058(input [0:0] sel);
    case (sel) 0: mux_3058 = 1'h0; 1: mux_3058 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3059;
  wire [0:0] v_3060;
  wire [0:0] v_3061;
  wire [0:0] v_3062;
  function [0:0] mux_3062(input [0:0] sel);
    case (sel) 0: mux_3062 = 1'h0; 1: mux_3062 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3063;
  function [0:0] mux_3063(input [0:0] sel);
    case (sel) 0: mux_3063 = 1'h0; 1: mux_3063 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3064;
  wire [0:0] v_3065;
  wire [0:0] v_3066;
  wire [0:0] v_3067;
  wire [0:0] v_3068;
  wire [0:0] v_3069;
  function [0:0] mux_3069(input [0:0] sel);
    case (sel) 0: mux_3069 = 1'h0; 1: mux_3069 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3070;
  function [0:0] mux_3070(input [0:0] sel);
    case (sel) 0: mux_3070 = 1'h0; 1: mux_3070 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3071;
  wire [0:0] v_3072;
  wire [0:0] v_3073;
  wire [0:0] v_3074;
  function [0:0] mux_3074(input [0:0] sel);
    case (sel) 0: mux_3074 = 1'h0; 1: mux_3074 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3075;
  function [0:0] mux_3075(input [0:0] sel);
    case (sel) 0: mux_3075 = 1'h0; 1: mux_3075 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3076;
  wire [0:0] v_3077;
  wire [0:0] v_3078;
  wire [0:0] v_3079;
  wire [0:0] v_3080;
  wire [0:0] v_3081;
  function [0:0] mux_3081(input [0:0] sel);
    case (sel) 0: mux_3081 = 1'h0; 1: mux_3081 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3082;
  function [0:0] mux_3082(input [0:0] sel);
    case (sel) 0: mux_3082 = 1'h0; 1: mux_3082 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3083;
  wire [0:0] v_3084;
  wire [0:0] v_3085;
  wire [0:0] v_3086;
  function [0:0] mux_3086(input [0:0] sel);
    case (sel) 0: mux_3086 = 1'h0; 1: mux_3086 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3087;
  function [0:0] mux_3087(input [0:0] sel);
    case (sel) 0: mux_3087 = 1'h0; 1: mux_3087 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3088;
  wire [0:0] v_3089;
  wire [0:0] v_3090;
  wire [0:0] v_3091;
  wire [0:0] v_3092;
  wire [0:0] v_3093;
  function [0:0] mux_3093(input [0:0] sel);
    case (sel) 0: mux_3093 = 1'h0; 1: mux_3093 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3094;
  wire [0:0] v_3095;
  function [0:0] mux_3095(input [0:0] sel);
    case (sel) 0: mux_3095 = 1'h0; 1: mux_3095 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3096;
  wire [0:0] v_3097;
  wire [0:0] v_3098;
  wire [0:0] v_3099;
  function [0:0] mux_3099(input [0:0] sel);
    case (sel) 0: mux_3099 = 1'h0; 1: mux_3099 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3100;
  function [0:0] mux_3100(input [0:0] sel);
    case (sel) 0: mux_3100 = 1'h0; 1: mux_3100 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3101 = 1'h0;
  wire [0:0] v_3102;
  wire [0:0] v_3103;
  wire [0:0] act_3104;
  wire [0:0] v_3105;
  wire [0:0] v_3106;
  wire [0:0] v_3107;
  reg [0:0] v_3108 = 1'h0;
  wire [0:0] v_3109;
  wire [0:0] v_3110;
  wire [0:0] act_3111;
  wire [0:0] v_3112;
  wire [0:0] v_3113;
  wire [0:0] v_3114;
  reg [0:0] v_3115 = 1'h0;
  wire [0:0] v_3116;
  wire [0:0] v_3117;
  wire [0:0] act_3118;
  wire [0:0] v_3119;
  wire [0:0] v_3120;
  wire [0:0] v_3121;
  reg [0:0] v_3122 = 1'h0;
  wire [0:0] v_3123;
  wire [0:0] v_3124;
  wire [0:0] act_3125;
  wire [0:0] v_3126;
  wire [0:0] v_3127;
  wire [0:0] v_3128;
  wire [0:0] v_3129;
  wire [0:0] v_3130;
  wire [0:0] v_3131;
  function [0:0] mux_3131(input [0:0] sel);
    case (sel) 0: mux_3131 = 1'h0; 1: mux_3131 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3132;
  wire [0:0] v_3133;
  function [0:0] mux_3133(input [0:0] sel);
    case (sel) 0: mux_3133 = 1'h0; 1: mux_3133 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3134;
  wire [0:0] v_3135;
  wire [0:0] v_3136;
  wire [0:0] v_3137;
  function [0:0] mux_3137(input [0:0] sel);
    case (sel) 0: mux_3137 = 1'h0; 1: mux_3137 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3138;
  function [0:0] mux_3138(input [0:0] sel);
    case (sel) 0: mux_3138 = 1'h0; 1: mux_3138 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3139 = 1'h0;
  wire [0:0] v_3140;
  wire [0:0] v_3141;
  wire [0:0] act_3142;
  wire [0:0] v_3143;
  wire [0:0] v_3144;
  wire [0:0] v_3145;
  wire [0:0] v_3146;
  wire [0:0] v_3147;
  wire [0:0] v_3148;
  function [0:0] mux_3148(input [0:0] sel);
    case (sel) 0: mux_3148 = 1'h0; 1: mux_3148 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3149;
  function [0:0] mux_3149(input [0:0] sel);
    case (sel) 0: mux_3149 = 1'h0; 1: mux_3149 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3150;
  wire [0:0] v_3151;
  wire [0:0] v_3152;
  wire [0:0] v_3153;
  function [0:0] mux_3153(input [0:0] sel);
    case (sel) 0: mux_3153 = 1'h0; 1: mux_3153 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3154;
  function [0:0] mux_3154(input [0:0] sel);
    case (sel) 0: mux_3154 = 1'h0; 1: mux_3154 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3155;
  wire [0:0] v_3156;
  wire [0:0] v_3157;
  wire [0:0] v_3158;
  wire [0:0] v_3159;
  wire [0:0] v_3160;
  function [0:0] mux_3160(input [0:0] sel);
    case (sel) 0: mux_3160 = 1'h0; 1: mux_3160 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3161;
  wire [0:0] v_3162;
  function [0:0] mux_3162(input [0:0] sel);
    case (sel) 0: mux_3162 = 1'h0; 1: mux_3162 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3163;
  wire [0:0] v_3164;
  wire [0:0] v_3165;
  wire [0:0] v_3166;
  function [0:0] mux_3166(input [0:0] sel);
    case (sel) 0: mux_3166 = 1'h0; 1: mux_3166 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3167;
  function [0:0] mux_3167(input [0:0] sel);
    case (sel) 0: mux_3167 = 1'h0; 1: mux_3167 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3168 = 1'h0;
  wire [0:0] v_3169;
  wire [0:0] v_3170;
  wire [0:0] act_3171;
  wire [0:0] v_3172;
  wire [0:0] v_3173;
  wire [0:0] v_3174;
  reg [0:0] v_3175 = 1'h0;
  wire [0:0] v_3176;
  wire [0:0] v_3177;
  wire [0:0] act_3178;
  wire [0:0] v_3179;
  wire [0:0] v_3180;
  wire [0:0] v_3181;
  wire [0:0] v_3182;
  wire [0:0] v_3183;
  wire [0:0] v_3184;
  function [0:0] mux_3184(input [0:0] sel);
    case (sel) 0: mux_3184 = 1'h0; 1: mux_3184 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3185;
  wire [0:0] v_3186;
  function [0:0] mux_3186(input [0:0] sel);
    case (sel) 0: mux_3186 = 1'h0; 1: mux_3186 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3187;
  wire [0:0] v_3188;
  wire [0:0] v_3189;
  wire [0:0] v_3190;
  function [0:0] mux_3190(input [0:0] sel);
    case (sel) 0: mux_3190 = 1'h0; 1: mux_3190 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3191;
  function [0:0] mux_3191(input [0:0] sel);
    case (sel) 0: mux_3191 = 1'h0; 1: mux_3191 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3192 = 1'h0;
  wire [0:0] v_3193;
  wire [0:0] v_3194;
  wire [0:0] act_3195;
  wire [0:0] v_3196;
  wire [0:0] v_3197;
  wire [0:0] v_3198;
  wire [0:0] v_3199;
  wire [0:0] v_3200;
  wire [0:0] v_3201;
  function [0:0] mux_3201(input [0:0] sel);
    case (sel) 0: mux_3201 = 1'h0; 1: mux_3201 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3202;
  function [0:0] mux_3202(input [0:0] sel);
    case (sel) 0: mux_3202 = 1'h0; 1: mux_3202 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3203;
  wire [0:0] v_3204;
  wire [0:0] v_3205;
  wire [0:0] v_3206;
  function [0:0] mux_3206(input [0:0] sel);
    case (sel) 0: mux_3206 = 1'h0; 1: mux_3206 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3207;
  function [0:0] mux_3207(input [0:0] sel);
    case (sel) 0: mux_3207 = 1'h0; 1: mux_3207 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3208;
  wire [0:0] v_3209;
  wire [0:0] v_3210;
  wire [0:0] v_3211;
  wire [0:0] v_3212;
  wire [0:0] v_3213;
  function [0:0] mux_3213(input [0:0] sel);
    case (sel) 0: mux_3213 = 1'h0; 1: mux_3213 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3214;
  function [0:0] mux_3214(input [0:0] sel);
    case (sel) 0: mux_3214 = 1'h0; 1: mux_3214 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3215;
  wire [0:0] v_3216;
  wire [0:0] v_3217;
  wire [0:0] v_3218;
  function [0:0] mux_3218(input [0:0] sel);
    case (sel) 0: mux_3218 = 1'h0; 1: mux_3218 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3219;
  function [0:0] mux_3219(input [0:0] sel);
    case (sel) 0: mux_3219 = 1'h0; 1: mux_3219 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3220;
  wire [0:0] v_3221;
  wire [0:0] v_3222;
  wire [0:0] v_3223;
  wire [0:0] v_3224;
  wire [0:0] v_3225;
  function [0:0] mux_3225(input [0:0] sel);
    case (sel) 0: mux_3225 = 1'h0; 1: mux_3225 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3226;
  wire [0:0] v_3227;
  function [0:0] mux_3227(input [0:0] sel);
    case (sel) 0: mux_3227 = 1'h0; 1: mux_3227 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3228;
  wire [0:0] v_3229;
  wire [0:0] v_3230;
  wire [0:0] v_3231;
  function [0:0] mux_3231(input [0:0] sel);
    case (sel) 0: mux_3231 = 1'h0; 1: mux_3231 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3232;
  function [0:0] mux_3232(input [0:0] sel);
    case (sel) 0: mux_3232 = 1'h0; 1: mux_3232 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3233 = 1'h0;
  wire [0:0] v_3234;
  wire [0:0] v_3235;
  wire [0:0] act_3236;
  wire [0:0] v_3237;
  wire [0:0] v_3238;
  wire [0:0] v_3239;
  reg [0:0] v_3240 = 1'h0;
  wire [0:0] v_3241;
  wire [0:0] v_3242;
  wire [0:0] act_3243;
  wire [0:0] v_3244;
  wire [0:0] v_3245;
  wire [0:0] v_3246;
  reg [0:0] v_3247 = 1'h0;
  wire [0:0] v_3248;
  wire [0:0] v_3249;
  wire [0:0] act_3250;
  wire [0:0] v_3251;
  wire [0:0] v_3252;
  wire [0:0] v_3253;
  wire [0:0] v_3254;
  wire [0:0] v_3255;
  wire [0:0] v_3256;
  function [0:0] mux_3256(input [0:0] sel);
    case (sel) 0: mux_3256 = 1'h0; 1: mux_3256 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3257;
  wire [0:0] v_3258;
  function [0:0] mux_3258(input [0:0] sel);
    case (sel) 0: mux_3258 = 1'h0; 1: mux_3258 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3259;
  wire [0:0] v_3260;
  wire [0:0] v_3261;
  wire [0:0] v_3262;
  function [0:0] mux_3262(input [0:0] sel);
    case (sel) 0: mux_3262 = 1'h0; 1: mux_3262 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3263;
  function [0:0] mux_3263(input [0:0] sel);
    case (sel) 0: mux_3263 = 1'h0; 1: mux_3263 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3264 = 1'h0;
  wire [0:0] v_3265;
  wire [0:0] v_3266;
  wire [0:0] act_3267;
  wire [0:0] v_3268;
  wire [0:0] v_3269;
  wire [0:0] v_3270;
  wire [0:0] v_3271;
  wire [0:0] v_3272;
  wire [0:0] v_3273;
  function [0:0] mux_3273(input [0:0] sel);
    case (sel) 0: mux_3273 = 1'h0; 1: mux_3273 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3274;
  function [0:0] mux_3274(input [0:0] sel);
    case (sel) 0: mux_3274 = 1'h0; 1: mux_3274 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3275;
  wire [0:0] v_3276;
  wire [0:0] v_3277;
  wire [0:0] v_3278;
  function [0:0] mux_3278(input [0:0] sel);
    case (sel) 0: mux_3278 = 1'h0; 1: mux_3278 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3279;
  function [0:0] mux_3279(input [0:0] sel);
    case (sel) 0: mux_3279 = 1'h0; 1: mux_3279 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3280;
  wire [0:0] v_3281;
  wire [0:0] v_3282;
  wire [0:0] v_3283;
  wire [0:0] v_3284;
  wire [0:0] v_3285;
  function [0:0] mux_3285(input [0:0] sel);
    case (sel) 0: mux_3285 = 1'h0; 1: mux_3285 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3286;
  wire [0:0] v_3287;
  function [0:0] mux_3287(input [0:0] sel);
    case (sel) 0: mux_3287 = 1'h0; 1: mux_3287 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3288;
  wire [0:0] v_3289;
  wire [0:0] v_3290;
  wire [0:0] v_3291;
  function [0:0] mux_3291(input [0:0] sel);
    case (sel) 0: mux_3291 = 1'h0; 1: mux_3291 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3292;
  function [0:0] mux_3292(input [0:0] sel);
    case (sel) 0: mux_3292 = 1'h0; 1: mux_3292 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3293 = 1'h0;
  wire [0:0] v_3294;
  wire [0:0] v_3295;
  wire [0:0] act_3296;
  wire [0:0] v_3297;
  wire [0:0] v_3298;
  wire [0:0] v_3299;
  reg [0:0] v_3300 = 1'h0;
  wire [0:0] v_3301;
  wire [0:0] v_3302;
  wire [0:0] act_3303;
  wire [0:0] v_3304;
  wire [0:0] v_3305;
  wire [0:0] v_3306;
  wire [0:0] v_3307;
  wire [0:0] v_3308;
  wire [0:0] v_3309;
  function [0:0] mux_3309(input [0:0] sel);
    case (sel) 0: mux_3309 = 1'h0; 1: mux_3309 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3310;
  wire [0:0] v_3311;
  function [0:0] mux_3311(input [0:0] sel);
    case (sel) 0: mux_3311 = 1'h0; 1: mux_3311 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3312;
  wire [0:0] v_3313;
  wire [0:0] v_3314;
  wire [0:0] v_3315;
  function [0:0] mux_3315(input [0:0] sel);
    case (sel) 0: mux_3315 = 1'h0; 1: mux_3315 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3316;
  function [0:0] mux_3316(input [0:0] sel);
    case (sel) 0: mux_3316 = 1'h0; 1: mux_3316 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3317 = 1'h0;
  wire [0:0] v_3318;
  wire [0:0] v_3319;
  wire [0:0] act_3320;
  wire [0:0] v_3321;
  wire [0:0] v_3322;
  wire [0:0] v_3323;
  wire [0:0] v_3324;
  wire [0:0] v_3325;
  wire [0:0] v_3326;
  function [0:0] mux_3326(input [0:0] sel);
    case (sel) 0: mux_3326 = 1'h0; 1: mux_3326 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3327;
  function [0:0] mux_3327(input [0:0] sel);
    case (sel) 0: mux_3327 = 1'h0; 1: mux_3327 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3328;
  wire [0:0] v_3329;
  wire [0:0] v_3330;
  wire [0:0] v_3331;
  function [0:0] mux_3331(input [0:0] sel);
    case (sel) 0: mux_3331 = 1'h0; 1: mux_3331 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3332;
  function [0:0] mux_3332(input [0:0] sel);
    case (sel) 0: mux_3332 = 1'h0; 1: mux_3332 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3333;
  wire [0:0] v_3334;
  wire [0:0] v_3335;
  wire [0:0] v_3336;
  wire [0:0] v_3337;
  wire [0:0] v_3338;
  function [0:0] mux_3338(input [0:0] sel);
    case (sel) 0: mux_3338 = 1'h0; 1: mux_3338 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3339;
  function [0:0] mux_3339(input [0:0] sel);
    case (sel) 0: mux_3339 = 1'h0; 1: mux_3339 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3340;
  wire [0:0] v_3341;
  wire [0:0] v_3342;
  wire [0:0] v_3343;
  function [0:0] mux_3343(input [0:0] sel);
    case (sel) 0: mux_3343 = 1'h0; 1: mux_3343 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3344;
  function [0:0] mux_3344(input [0:0] sel);
    case (sel) 0: mux_3344 = 1'h0; 1: mux_3344 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3345;
  wire [0:0] v_3346;
  wire [0:0] v_3347;
  wire [0:0] v_3348;
  wire [0:0] v_3349;
  wire [0:0] v_3350;
  function [0:0] mux_3350(input [0:0] sel);
    case (sel) 0: mux_3350 = 1'h0; 1: mux_3350 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3351;
  function [0:0] mux_3351(input [0:0] sel);
    case (sel) 0: mux_3351 = 1'h0; 1: mux_3351 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3352;
  wire [0:0] v_3353;
  wire [0:0] v_3354;
  wire [0:0] v_3355;
  function [0:0] mux_3355(input [0:0] sel);
    case (sel) 0: mux_3355 = 1'h0; 1: mux_3355 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3356;
  function [0:0] mux_3356(input [0:0] sel);
    case (sel) 0: mux_3356 = 1'h0; 1: mux_3356 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3357;
  wire [0:0] v_3358;
  wire [0:0] v_3359;
  wire [0:0] v_3360;
  wire [0:0] v_3361;
  wire [0:0] v_3362;
  function [0:0] mux_3362(input [0:0] sel);
    case (sel) 0: mux_3362 = 1'h0; 1: mux_3362 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3363;
  function [0:0] mux_3363(input [0:0] sel);
    case (sel) 0: mux_3363 = 1'h0; 1: mux_3363 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3364;
  wire [0:0] v_3365;
  wire [0:0] v_3366;
  wire [0:0] v_3367;
  function [0:0] mux_3367(input [0:0] sel);
    case (sel) 0: mux_3367 = 1'h0; 1: mux_3367 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3368;
  function [0:0] mux_3368(input [0:0] sel);
    case (sel) 0: mux_3368 = 1'h0; 1: mux_3368 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3369;
  wire [0:0] v_3370;
  wire [0:0] v_3371;
  wire [0:0] v_3372;
  wire [0:0] v_3373;
  wire [0:0] v_3374;
  function [0:0] mux_3374(input [0:0] sel);
    case (sel) 0: mux_3374 = 1'h0; 1: mux_3374 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3375;
  wire [0:0] v_3376;
  function [0:0] mux_3376(input [0:0] sel);
    case (sel) 0: mux_3376 = 1'h0; 1: mux_3376 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3377;
  wire [0:0] v_3378;
  wire [0:0] v_3379;
  wire [0:0] v_3380;
  function [0:0] mux_3380(input [0:0] sel);
    case (sel) 0: mux_3380 = 1'h0; 1: mux_3380 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3381;
  function [0:0] mux_3381(input [0:0] sel);
    case (sel) 0: mux_3381 = 1'h0; 1: mux_3381 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3382 = 1'h0;
  wire [0:0] v_3383;
  wire [0:0] v_3384;
  wire [0:0] act_3385;
  wire [0:0] v_3386;
  wire [0:0] v_3387;
  wire [0:0] v_3388;
  reg [0:0] v_3389 = 1'h0;
  wire [0:0] v_3390;
  wire [0:0] v_3391;
  wire [0:0] act_3392;
  wire [0:0] v_3393;
  wire [0:0] v_3394;
  wire [0:0] v_3395;
  reg [0:0] v_3396 = 1'h0;
  wire [0:0] v_3397;
  wire [0:0] v_3398;
  wire [0:0] act_3399;
  wire [0:0] v_3400;
  wire [0:0] v_3401;
  wire [0:0] v_3402;
  reg [0:0] v_3403 = 1'h0;
  wire [0:0] v_3404;
  wire [0:0] v_3405;
  wire [0:0] act_3406;
  wire [0:0] v_3407;
  wire [0:0] v_3408;
  wire [0:0] v_3409;
  reg [0:0] v_3410 = 1'h0;
  wire [0:0] v_3411;
  wire [0:0] v_3412;
  wire [0:0] act_3413;
  wire [0:0] v_3414;
  wire [0:0] v_3415;
  wire [0:0] v_3416;
  wire [0:0] v_3417;
  wire [0:0] v_3418;
  wire [0:0] v_3419;
  function [0:0] mux_3419(input [0:0] sel);
    case (sel) 0: mux_3419 = 1'h0; 1: mux_3419 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3420;
  wire [0:0] v_3421;
  function [0:0] mux_3421(input [0:0] sel);
    case (sel) 0: mux_3421 = 1'h0; 1: mux_3421 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3422;
  wire [0:0] v_3423;
  wire [0:0] v_3424;
  wire [0:0] v_3425;
  function [0:0] mux_3425(input [0:0] sel);
    case (sel) 0: mux_3425 = 1'h0; 1: mux_3425 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3426;
  function [0:0] mux_3426(input [0:0] sel);
    case (sel) 0: mux_3426 = 1'h0; 1: mux_3426 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3427 = 1'h0;
  wire [0:0] v_3428;
  wire [0:0] v_3429;
  wire [0:0] act_3430;
  wire [0:0] v_3431;
  wire [0:0] v_3432;
  wire [0:0] v_3433;
  wire [0:0] v_3434;
  wire [0:0] v_3435;
  wire [0:0] v_3436;
  function [0:0] mux_3436(input [0:0] sel);
    case (sel) 0: mux_3436 = 1'h0; 1: mux_3436 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3437;
  function [0:0] mux_3437(input [0:0] sel);
    case (sel) 0: mux_3437 = 1'h0; 1: mux_3437 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3438;
  wire [0:0] v_3439;
  wire [0:0] v_3440;
  wire [0:0] v_3441;
  function [0:0] mux_3441(input [0:0] sel);
    case (sel) 0: mux_3441 = 1'h0; 1: mux_3441 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3442;
  function [0:0] mux_3442(input [0:0] sel);
    case (sel) 0: mux_3442 = 1'h0; 1: mux_3442 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3443;
  wire [0:0] v_3444;
  wire [0:0] v_3445;
  wire [0:0] v_3446;
  wire [0:0] v_3447;
  wire [0:0] v_3448;
  function [0:0] mux_3448(input [0:0] sel);
    case (sel) 0: mux_3448 = 1'h0; 1: mux_3448 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3449;
  wire [0:0] v_3450;
  function [0:0] mux_3450(input [0:0] sel);
    case (sel) 0: mux_3450 = 1'h0; 1: mux_3450 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3451;
  wire [0:0] v_3452;
  wire [0:0] v_3453;
  wire [0:0] v_3454;
  function [0:0] mux_3454(input [0:0] sel);
    case (sel) 0: mux_3454 = 1'h0; 1: mux_3454 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3455;
  function [0:0] mux_3455(input [0:0] sel);
    case (sel) 0: mux_3455 = 1'h0; 1: mux_3455 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3456 = 1'h0;
  wire [0:0] v_3457;
  wire [0:0] v_3458;
  wire [0:0] act_3459;
  wire [0:0] v_3460;
  wire [0:0] v_3461;
  wire [0:0] v_3462;
  reg [0:0] v_3463 = 1'h0;
  wire [0:0] v_3464;
  wire [0:0] v_3465;
  wire [0:0] act_3466;
  wire [0:0] v_3467;
  wire [0:0] v_3468;
  wire [0:0] v_3469;
  wire [0:0] v_3470;
  wire [0:0] v_3471;
  wire [0:0] v_3472;
  function [0:0] mux_3472(input [0:0] sel);
    case (sel) 0: mux_3472 = 1'h0; 1: mux_3472 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3473;
  wire [0:0] v_3474;
  function [0:0] mux_3474(input [0:0] sel);
    case (sel) 0: mux_3474 = 1'h0; 1: mux_3474 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3475;
  wire [0:0] v_3476;
  wire [0:0] v_3477;
  wire [0:0] v_3478;
  function [0:0] mux_3478(input [0:0] sel);
    case (sel) 0: mux_3478 = 1'h0; 1: mux_3478 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3479;
  function [0:0] mux_3479(input [0:0] sel);
    case (sel) 0: mux_3479 = 1'h0; 1: mux_3479 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3480 = 1'h0;
  wire [0:0] v_3481;
  wire [0:0] v_3482;
  wire [0:0] act_3483;
  wire [0:0] v_3484;
  wire [0:0] v_3485;
  wire [0:0] v_3486;
  wire [0:0] v_3487;
  wire [0:0] v_3488;
  wire [0:0] v_3489;
  function [0:0] mux_3489(input [0:0] sel);
    case (sel) 0: mux_3489 = 1'h0; 1: mux_3489 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3490;
  function [0:0] mux_3490(input [0:0] sel);
    case (sel) 0: mux_3490 = 1'h0; 1: mux_3490 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3491;
  wire [0:0] v_3492;
  wire [0:0] v_3493;
  wire [0:0] v_3494;
  function [0:0] mux_3494(input [0:0] sel);
    case (sel) 0: mux_3494 = 1'h0; 1: mux_3494 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3495;
  function [0:0] mux_3495(input [0:0] sel);
    case (sel) 0: mux_3495 = 1'h0; 1: mux_3495 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3496;
  wire [0:0] v_3497;
  wire [0:0] v_3498;
  wire [0:0] v_3499;
  wire [0:0] v_3500;
  wire [0:0] v_3501;
  function [0:0] mux_3501(input [0:0] sel);
    case (sel) 0: mux_3501 = 1'h0; 1: mux_3501 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3502;
  function [0:0] mux_3502(input [0:0] sel);
    case (sel) 0: mux_3502 = 1'h0; 1: mux_3502 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3503;
  wire [0:0] v_3504;
  wire [0:0] v_3505;
  wire [0:0] v_3506;
  function [0:0] mux_3506(input [0:0] sel);
    case (sel) 0: mux_3506 = 1'h0; 1: mux_3506 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3507;
  function [0:0] mux_3507(input [0:0] sel);
    case (sel) 0: mux_3507 = 1'h0; 1: mux_3507 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3508;
  wire [0:0] v_3509;
  wire [0:0] v_3510;
  wire [0:0] v_3511;
  wire [0:0] v_3512;
  wire [0:0] v_3513;
  function [0:0] mux_3513(input [0:0] sel);
    case (sel) 0: mux_3513 = 1'h0; 1: mux_3513 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3514;
  wire [0:0] v_3515;
  function [0:0] mux_3515(input [0:0] sel);
    case (sel) 0: mux_3515 = 1'h0; 1: mux_3515 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3516;
  wire [0:0] v_3517;
  wire [0:0] v_3518;
  wire [0:0] v_3519;
  function [0:0] mux_3519(input [0:0] sel);
    case (sel) 0: mux_3519 = 1'h0; 1: mux_3519 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3520;
  function [0:0] mux_3520(input [0:0] sel);
    case (sel) 0: mux_3520 = 1'h0; 1: mux_3520 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3521 = 1'h0;
  wire [0:0] v_3522;
  wire [0:0] v_3523;
  wire [0:0] act_3524;
  wire [0:0] v_3525;
  wire [0:0] v_3526;
  wire [0:0] v_3527;
  reg [0:0] v_3528 = 1'h0;
  wire [0:0] v_3529;
  wire [0:0] v_3530;
  wire [0:0] act_3531;
  wire [0:0] v_3532;
  wire [0:0] v_3533;
  wire [0:0] v_3534;
  reg [0:0] v_3535 = 1'h0;
  wire [0:0] v_3536;
  wire [0:0] v_3537;
  wire [0:0] act_3538;
  wire [0:0] v_3539;
  wire [0:0] v_3540;
  wire [0:0] v_3541;
  wire [0:0] v_3542;
  wire [0:0] v_3543;
  wire [0:0] v_3544;
  function [0:0] mux_3544(input [0:0] sel);
    case (sel) 0: mux_3544 = 1'h0; 1: mux_3544 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3545;
  wire [0:0] v_3546;
  function [0:0] mux_3546(input [0:0] sel);
    case (sel) 0: mux_3546 = 1'h0; 1: mux_3546 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3547;
  wire [0:0] v_3548;
  wire [0:0] v_3549;
  wire [0:0] v_3550;
  function [0:0] mux_3550(input [0:0] sel);
    case (sel) 0: mux_3550 = 1'h0; 1: mux_3550 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3551;
  function [0:0] mux_3551(input [0:0] sel);
    case (sel) 0: mux_3551 = 1'h0; 1: mux_3551 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3552 = 1'h0;
  wire [0:0] v_3553;
  wire [0:0] v_3554;
  wire [0:0] act_3555;
  wire [0:0] v_3556;
  wire [0:0] v_3557;
  wire [0:0] v_3558;
  wire [0:0] v_3559;
  wire [0:0] v_3560;
  wire [0:0] v_3561;
  function [0:0] mux_3561(input [0:0] sel);
    case (sel) 0: mux_3561 = 1'h0; 1: mux_3561 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3562;
  function [0:0] mux_3562(input [0:0] sel);
    case (sel) 0: mux_3562 = 1'h0; 1: mux_3562 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3563;
  wire [0:0] v_3564;
  wire [0:0] v_3565;
  wire [0:0] v_3566;
  function [0:0] mux_3566(input [0:0] sel);
    case (sel) 0: mux_3566 = 1'h0; 1: mux_3566 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3567;
  function [0:0] mux_3567(input [0:0] sel);
    case (sel) 0: mux_3567 = 1'h0; 1: mux_3567 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3568;
  wire [0:0] v_3569;
  wire [0:0] v_3570;
  wire [0:0] v_3571;
  wire [0:0] v_3572;
  wire [0:0] v_3573;
  function [0:0] mux_3573(input [0:0] sel);
    case (sel) 0: mux_3573 = 1'h0; 1: mux_3573 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3574;
  wire [0:0] v_3575;
  function [0:0] mux_3575(input [0:0] sel);
    case (sel) 0: mux_3575 = 1'h0; 1: mux_3575 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3576;
  wire [0:0] v_3577;
  wire [0:0] v_3578;
  wire [0:0] v_3579;
  function [0:0] mux_3579(input [0:0] sel);
    case (sel) 0: mux_3579 = 1'h0; 1: mux_3579 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3580;
  function [0:0] mux_3580(input [0:0] sel);
    case (sel) 0: mux_3580 = 1'h0; 1: mux_3580 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3581 = 1'h0;
  wire [0:0] v_3582;
  wire [0:0] v_3583;
  wire [0:0] act_3584;
  wire [0:0] v_3585;
  wire [0:0] v_3586;
  wire [0:0] v_3587;
  reg [0:0] v_3588 = 1'h0;
  wire [0:0] v_3589;
  wire [0:0] v_3590;
  wire [0:0] act_3591;
  wire [0:0] v_3592;
  wire [0:0] v_3593;
  wire [0:0] v_3594;
  wire [0:0] v_3595;
  wire [0:0] v_3596;
  wire [0:0] v_3597;
  function [0:0] mux_3597(input [0:0] sel);
    case (sel) 0: mux_3597 = 1'h0; 1: mux_3597 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3598;
  wire [0:0] v_3599;
  function [0:0] mux_3599(input [0:0] sel);
    case (sel) 0: mux_3599 = 1'h0; 1: mux_3599 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3600;
  wire [0:0] v_3601;
  wire [0:0] v_3602;
  wire [0:0] v_3603;
  function [0:0] mux_3603(input [0:0] sel);
    case (sel) 0: mux_3603 = 1'h0; 1: mux_3603 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3604;
  function [0:0] mux_3604(input [0:0] sel);
    case (sel) 0: mux_3604 = 1'h0; 1: mux_3604 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3605 = 1'h0;
  wire [0:0] v_3606;
  wire [0:0] v_3607;
  wire [0:0] act_3608;
  wire [0:0] v_3609;
  wire [0:0] v_3610;
  wire [0:0] v_3611;
  wire [0:0] v_3612;
  wire [0:0] v_3613;
  wire [0:0] v_3614;
  function [0:0] mux_3614(input [0:0] sel);
    case (sel) 0: mux_3614 = 1'h0; 1: mux_3614 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3615;
  function [0:0] mux_3615(input [0:0] sel);
    case (sel) 0: mux_3615 = 1'h0; 1: mux_3615 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3616;
  wire [0:0] v_3617;
  wire [0:0] v_3618;
  wire [0:0] v_3619;
  function [0:0] mux_3619(input [0:0] sel);
    case (sel) 0: mux_3619 = 1'h0; 1: mux_3619 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3620;
  function [0:0] mux_3620(input [0:0] sel);
    case (sel) 0: mux_3620 = 1'h0; 1: mux_3620 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3621;
  wire [0:0] v_3622;
  wire [0:0] v_3623;
  wire [0:0] v_3624;
  wire [0:0] v_3625;
  wire [0:0] v_3626;
  function [0:0] mux_3626(input [0:0] sel);
    case (sel) 0: mux_3626 = 1'h0; 1: mux_3626 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3627;
  function [0:0] mux_3627(input [0:0] sel);
    case (sel) 0: mux_3627 = 1'h0; 1: mux_3627 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3628;
  wire [0:0] v_3629;
  wire [0:0] v_3630;
  wire [0:0] v_3631;
  function [0:0] mux_3631(input [0:0] sel);
    case (sel) 0: mux_3631 = 1'h0; 1: mux_3631 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3632;
  function [0:0] mux_3632(input [0:0] sel);
    case (sel) 0: mux_3632 = 1'h0; 1: mux_3632 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3633;
  wire [0:0] v_3634;
  wire [0:0] v_3635;
  wire [0:0] v_3636;
  wire [0:0] v_3637;
  wire [0:0] v_3638;
  function [0:0] mux_3638(input [0:0] sel);
    case (sel) 0: mux_3638 = 1'h0; 1: mux_3638 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3639;
  function [0:0] mux_3639(input [0:0] sel);
    case (sel) 0: mux_3639 = 1'h0; 1: mux_3639 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3640;
  wire [0:0] v_3641;
  wire [0:0] v_3642;
  wire [0:0] v_3643;
  function [0:0] mux_3643(input [0:0] sel);
    case (sel) 0: mux_3643 = 1'h0; 1: mux_3643 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3644;
  function [0:0] mux_3644(input [0:0] sel);
    case (sel) 0: mux_3644 = 1'h0; 1: mux_3644 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3645;
  wire [0:0] v_3646;
  wire [0:0] v_3647;
  wire [0:0] v_3648;
  wire [0:0] v_3649;
  wire [0:0] v_3650;
  function [0:0] mux_3650(input [0:0] sel);
    case (sel) 0: mux_3650 = 1'h0; 1: mux_3650 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3651;
  wire [0:0] v_3652;
  function [0:0] mux_3652(input [0:0] sel);
    case (sel) 0: mux_3652 = 1'h0; 1: mux_3652 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3653;
  wire [0:0] v_3654;
  wire [0:0] v_3655;
  wire [0:0] v_3656;
  function [0:0] mux_3656(input [0:0] sel);
    case (sel) 0: mux_3656 = 1'h0; 1: mux_3656 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3657;
  function [0:0] mux_3657(input [0:0] sel);
    case (sel) 0: mux_3657 = 1'h0; 1: mux_3657 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3658 = 1'h0;
  wire [0:0] v_3659;
  wire [0:0] v_3660;
  wire [0:0] act_3661;
  wire [0:0] v_3662;
  wire [0:0] v_3663;
  wire [0:0] v_3664;
  reg [0:0] v_3665 = 1'h0;
  wire [0:0] v_3666;
  wire [0:0] v_3667;
  wire [0:0] act_3668;
  wire [0:0] v_3669;
  wire [0:0] v_3670;
  wire [0:0] v_3671;
  reg [0:0] v_3672 = 1'h0;
  wire [0:0] v_3673;
  wire [0:0] v_3674;
  wire [0:0] act_3675;
  wire [0:0] v_3676;
  wire [0:0] v_3677;
  wire [0:0] v_3678;
  reg [0:0] v_3679 = 1'h0;
  wire [0:0] v_3680;
  wire [0:0] v_3681;
  wire [0:0] act_3682;
  wire [0:0] v_3683;
  wire [0:0] v_3684;
  wire [0:0] v_3685;
  wire [0:0] v_3686;
  wire [0:0] v_3687;
  wire [0:0] v_3688;
  function [0:0] mux_3688(input [0:0] sel);
    case (sel) 0: mux_3688 = 1'h0; 1: mux_3688 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3689;
  wire [0:0] v_3690;
  function [0:0] mux_3690(input [0:0] sel);
    case (sel) 0: mux_3690 = 1'h0; 1: mux_3690 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3691;
  wire [0:0] v_3692;
  wire [0:0] v_3693;
  wire [0:0] v_3694;
  function [0:0] mux_3694(input [0:0] sel);
    case (sel) 0: mux_3694 = 1'h0; 1: mux_3694 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3695;
  function [0:0] mux_3695(input [0:0] sel);
    case (sel) 0: mux_3695 = 1'h0; 1: mux_3695 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3696 = 1'h0;
  wire [0:0] v_3697;
  wire [0:0] v_3698;
  wire [0:0] act_3699;
  wire [0:0] v_3700;
  wire [0:0] v_3701;
  wire [0:0] v_3702;
  wire [0:0] v_3703;
  wire [0:0] v_3704;
  wire [0:0] v_3705;
  function [0:0] mux_3705(input [0:0] sel);
    case (sel) 0: mux_3705 = 1'h0; 1: mux_3705 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3706;
  function [0:0] mux_3706(input [0:0] sel);
    case (sel) 0: mux_3706 = 1'h0; 1: mux_3706 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3707;
  wire [0:0] v_3708;
  wire [0:0] v_3709;
  wire [0:0] v_3710;
  function [0:0] mux_3710(input [0:0] sel);
    case (sel) 0: mux_3710 = 1'h0; 1: mux_3710 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3711;
  function [0:0] mux_3711(input [0:0] sel);
    case (sel) 0: mux_3711 = 1'h0; 1: mux_3711 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3712;
  wire [0:0] v_3713;
  wire [0:0] v_3714;
  wire [0:0] v_3715;
  wire [0:0] v_3716;
  wire [0:0] v_3717;
  function [0:0] mux_3717(input [0:0] sel);
    case (sel) 0: mux_3717 = 1'h0; 1: mux_3717 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3718;
  wire [0:0] v_3719;
  function [0:0] mux_3719(input [0:0] sel);
    case (sel) 0: mux_3719 = 1'h0; 1: mux_3719 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3720;
  wire [0:0] v_3721;
  wire [0:0] v_3722;
  wire [0:0] v_3723;
  function [0:0] mux_3723(input [0:0] sel);
    case (sel) 0: mux_3723 = 1'h0; 1: mux_3723 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3724;
  function [0:0] mux_3724(input [0:0] sel);
    case (sel) 0: mux_3724 = 1'h0; 1: mux_3724 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3725 = 1'h0;
  wire [0:0] v_3726;
  wire [0:0] v_3727;
  wire [0:0] act_3728;
  wire [0:0] v_3729;
  wire [0:0] v_3730;
  wire [0:0] v_3731;
  reg [0:0] v_3732 = 1'h0;
  wire [0:0] v_3733;
  wire [0:0] v_3734;
  wire [0:0] act_3735;
  wire [0:0] v_3736;
  wire [0:0] v_3737;
  wire [0:0] v_3738;
  wire [0:0] v_3739;
  wire [0:0] v_3740;
  wire [0:0] v_3741;
  function [0:0] mux_3741(input [0:0] sel);
    case (sel) 0: mux_3741 = 1'h0; 1: mux_3741 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3742;
  wire [0:0] v_3743;
  function [0:0] mux_3743(input [0:0] sel);
    case (sel) 0: mux_3743 = 1'h0; 1: mux_3743 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3744;
  wire [0:0] v_3745;
  wire [0:0] v_3746;
  wire [0:0] v_3747;
  function [0:0] mux_3747(input [0:0] sel);
    case (sel) 0: mux_3747 = 1'h0; 1: mux_3747 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3748;
  function [0:0] mux_3748(input [0:0] sel);
    case (sel) 0: mux_3748 = 1'h0; 1: mux_3748 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3749 = 1'h0;
  wire [0:0] v_3750;
  wire [0:0] v_3751;
  wire [0:0] act_3752;
  wire [0:0] v_3753;
  wire [0:0] v_3754;
  wire [0:0] v_3755;
  wire [0:0] v_3756;
  wire [0:0] v_3757;
  wire [0:0] v_3758;
  function [0:0] mux_3758(input [0:0] sel);
    case (sel) 0: mux_3758 = 1'h0; 1: mux_3758 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3759;
  function [0:0] mux_3759(input [0:0] sel);
    case (sel) 0: mux_3759 = 1'h0; 1: mux_3759 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3760;
  wire [0:0] v_3761;
  wire [0:0] v_3762;
  wire [0:0] v_3763;
  function [0:0] mux_3763(input [0:0] sel);
    case (sel) 0: mux_3763 = 1'h0; 1: mux_3763 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3764;
  function [0:0] mux_3764(input [0:0] sel);
    case (sel) 0: mux_3764 = 1'h0; 1: mux_3764 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3765;
  wire [0:0] v_3766;
  wire [0:0] v_3767;
  wire [0:0] v_3768;
  wire [0:0] v_3769;
  wire [0:0] v_3770;
  function [0:0] mux_3770(input [0:0] sel);
    case (sel) 0: mux_3770 = 1'h0; 1: mux_3770 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3771;
  function [0:0] mux_3771(input [0:0] sel);
    case (sel) 0: mux_3771 = 1'h0; 1: mux_3771 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3772;
  wire [0:0] v_3773;
  wire [0:0] v_3774;
  wire [0:0] v_3775;
  function [0:0] mux_3775(input [0:0] sel);
    case (sel) 0: mux_3775 = 1'h0; 1: mux_3775 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3776;
  function [0:0] mux_3776(input [0:0] sel);
    case (sel) 0: mux_3776 = 1'h0; 1: mux_3776 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3777;
  wire [0:0] v_3778;
  wire [0:0] v_3779;
  wire [0:0] v_3780;
  wire [0:0] v_3781;
  wire [0:0] v_3782;
  function [0:0] mux_3782(input [0:0] sel);
    case (sel) 0: mux_3782 = 1'h0; 1: mux_3782 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3783;
  wire [0:0] v_3784;
  function [0:0] mux_3784(input [0:0] sel);
    case (sel) 0: mux_3784 = 1'h0; 1: mux_3784 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3785;
  wire [0:0] v_3786;
  wire [0:0] v_3787;
  wire [0:0] v_3788;
  function [0:0] mux_3788(input [0:0] sel);
    case (sel) 0: mux_3788 = 1'h0; 1: mux_3788 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3789;
  function [0:0] mux_3789(input [0:0] sel);
    case (sel) 0: mux_3789 = 1'h0; 1: mux_3789 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3790 = 1'h0;
  wire [0:0] v_3791;
  wire [0:0] v_3792;
  wire [0:0] act_3793;
  wire [0:0] v_3794;
  wire [0:0] v_3795;
  wire [0:0] v_3796;
  reg [0:0] v_3797 = 1'h0;
  wire [0:0] v_3798;
  wire [0:0] v_3799;
  wire [0:0] act_3800;
  wire [0:0] v_3801;
  wire [0:0] v_3802;
  wire [0:0] v_3803;
  reg [0:0] v_3804 = 1'h0;
  wire [0:0] v_3805;
  wire [0:0] v_3806;
  wire [0:0] act_3807;
  wire [0:0] v_3808;
  wire [0:0] v_3809;
  wire [0:0] v_3810;
  wire [0:0] v_3811;
  wire [0:0] v_3812;
  wire [0:0] v_3813;
  function [0:0] mux_3813(input [0:0] sel);
    case (sel) 0: mux_3813 = 1'h0; 1: mux_3813 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3814;
  wire [0:0] v_3815;
  function [0:0] mux_3815(input [0:0] sel);
    case (sel) 0: mux_3815 = 1'h0; 1: mux_3815 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3816;
  wire [0:0] v_3817;
  wire [0:0] v_3818;
  wire [0:0] v_3819;
  function [0:0] mux_3819(input [0:0] sel);
    case (sel) 0: mux_3819 = 1'h0; 1: mux_3819 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3820;
  function [0:0] mux_3820(input [0:0] sel);
    case (sel) 0: mux_3820 = 1'h0; 1: mux_3820 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3821 = 1'h0;
  wire [0:0] v_3822;
  wire [0:0] v_3823;
  wire [0:0] act_3824;
  wire [0:0] v_3825;
  wire [0:0] v_3826;
  wire [0:0] v_3827;
  wire [0:0] v_3828;
  wire [0:0] v_3829;
  wire [0:0] v_3830;
  function [0:0] mux_3830(input [0:0] sel);
    case (sel) 0: mux_3830 = 1'h0; 1: mux_3830 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3831;
  function [0:0] mux_3831(input [0:0] sel);
    case (sel) 0: mux_3831 = 1'h0; 1: mux_3831 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3832;
  wire [0:0] v_3833;
  wire [0:0] v_3834;
  wire [0:0] v_3835;
  function [0:0] mux_3835(input [0:0] sel);
    case (sel) 0: mux_3835 = 1'h0; 1: mux_3835 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3836;
  function [0:0] mux_3836(input [0:0] sel);
    case (sel) 0: mux_3836 = 1'h0; 1: mux_3836 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3837;
  wire [0:0] v_3838;
  wire [0:0] v_3839;
  wire [0:0] v_3840;
  wire [0:0] v_3841;
  wire [0:0] v_3842;
  function [0:0] mux_3842(input [0:0] sel);
    case (sel) 0: mux_3842 = 1'h0; 1: mux_3842 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3843;
  wire [0:0] v_3844;
  function [0:0] mux_3844(input [0:0] sel);
    case (sel) 0: mux_3844 = 1'h0; 1: mux_3844 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3845;
  wire [0:0] v_3846;
  wire [0:0] v_3847;
  wire [0:0] v_3848;
  function [0:0] mux_3848(input [0:0] sel);
    case (sel) 0: mux_3848 = 1'h0; 1: mux_3848 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3849;
  function [0:0] mux_3849(input [0:0] sel);
    case (sel) 0: mux_3849 = 1'h0; 1: mux_3849 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3850 = 1'h0;
  wire [0:0] v_3851;
  wire [0:0] v_3852;
  wire [0:0] act_3853;
  wire [0:0] v_3854;
  wire [0:0] v_3855;
  wire [0:0] v_3856;
  reg [0:0] v_3857 = 1'h0;
  wire [0:0] v_3858;
  wire [0:0] v_3859;
  wire [0:0] act_3860;
  wire [0:0] v_3861;
  wire [0:0] v_3862;
  wire [0:0] v_3863;
  wire [0:0] v_3864;
  wire [0:0] v_3865;
  wire [0:0] v_3866;
  function [0:0] mux_3866(input [0:0] sel);
    case (sel) 0: mux_3866 = 1'h0; 1: mux_3866 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3867;
  wire [0:0] v_3868;
  function [0:0] mux_3868(input [0:0] sel);
    case (sel) 0: mux_3868 = 1'h0; 1: mux_3868 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3869;
  wire [0:0] v_3870;
  wire [0:0] v_3871;
  wire [0:0] v_3872;
  function [0:0] mux_3872(input [0:0] sel);
    case (sel) 0: mux_3872 = 1'h0; 1: mux_3872 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3873;
  function [0:0] mux_3873(input [0:0] sel);
    case (sel) 0: mux_3873 = 1'h0; 1: mux_3873 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3874 = 1'h0;
  wire [0:0] v_3875;
  wire [0:0] v_3876;
  wire [0:0] act_3877;
  wire [0:0] v_3878;
  wire [0:0] v_3879;
  wire [0:0] v_3880;
  wire [0:0] v_3881;
  wire [0:0] v_3882;
  wire [0:0] v_3883;
  function [0:0] mux_3883(input [0:0] sel);
    case (sel) 0: mux_3883 = 1'h0; 1: mux_3883 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3884;
  function [0:0] mux_3884(input [0:0] sel);
    case (sel) 0: mux_3884 = 1'h0; 1: mux_3884 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3885;
  wire [0:0] v_3886;
  wire [0:0] v_3887;
  wire [0:0] v_3888;
  function [0:0] mux_3888(input [0:0] sel);
    case (sel) 0: mux_3888 = 1'h0; 1: mux_3888 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3889;
  function [0:0] mux_3889(input [0:0] sel);
    case (sel) 0: mux_3889 = 1'h0; 1: mux_3889 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3890;
  wire [0:0] v_3891;
  wire [0:0] v_3892;
  wire [0:0] v_3893;
  wire [0:0] v_3894;
  wire [0:0] v_3895;
  function [0:0] mux_3895(input [0:0] sel);
    case (sel) 0: mux_3895 = 1'h0; 1: mux_3895 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3896;
  function [0:0] mux_3896(input [0:0] sel);
    case (sel) 0: mux_3896 = 1'h0; 1: mux_3896 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3897;
  wire [0:0] v_3898;
  wire [0:0] v_3899;
  wire [0:0] v_3900;
  function [0:0] mux_3900(input [0:0] sel);
    case (sel) 0: mux_3900 = 1'h0; 1: mux_3900 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3901;
  function [0:0] mux_3901(input [0:0] sel);
    case (sel) 0: mux_3901 = 1'h0; 1: mux_3901 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3902;
  wire [0:0] v_3903;
  wire [0:0] v_3904;
  wire [0:0] v_3905;
  wire [0:0] v_3906;
  wire [0:0] v_3907;
  function [0:0] mux_3907(input [0:0] sel);
    case (sel) 0: mux_3907 = 1'h0; 1: mux_3907 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3908;
  function [0:0] mux_3908(input [0:0] sel);
    case (sel) 0: mux_3908 = 1'h0; 1: mux_3908 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3909;
  wire [0:0] v_3910;
  wire [0:0] v_3911;
  wire [0:0] v_3912;
  function [0:0] mux_3912(input [0:0] sel);
    case (sel) 0: mux_3912 = 1'h0; 1: mux_3912 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3913;
  function [0:0] mux_3913(input [0:0] sel);
    case (sel) 0: mux_3913 = 1'h0; 1: mux_3913 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3914;
  wire [0:0] v_3915;
  wire [0:0] v_3916;
  wire [0:0] v_3917;
  wire [0:0] v_3918;
  wire [0:0] v_3919;
  function [0:0] mux_3919(input [0:0] sel);
    case (sel) 0: mux_3919 = 1'h0; 1: mux_3919 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3920;
  function [0:0] mux_3920(input [0:0] sel);
    case (sel) 0: mux_3920 = 1'h0; 1: mux_3920 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3921;
  wire [0:0] v_3922;
  wire [0:0] v_3923;
  wire [0:0] v_3924;
  function [0:0] mux_3924(input [0:0] sel);
    case (sel) 0: mux_3924 = 1'h0; 1: mux_3924 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3925;
  function [0:0] mux_3925(input [0:0] sel);
    case (sel) 0: mux_3925 = 1'h0; 1: mux_3925 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3926;
  wire [0:0] v_3927;
  wire [0:0] v_3928;
  wire [0:0] v_3929;
  wire [0:0] v_3930;
  wire [0:0] v_3931;
  function [0:0] mux_3931(input [0:0] sel);
    case (sel) 0: mux_3931 = 1'h0; 1: mux_3931 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3932;
  function [0:0] mux_3932(input [0:0] sel);
    case (sel) 0: mux_3932 = 1'h0; 1: mux_3932 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3933;
  wire [0:0] v_3934;
  wire [0:0] v_3935;
  wire [0:0] v_3936;
  function [0:0] mux_3936(input [0:0] sel);
    case (sel) 0: mux_3936 = 1'h0; 1: mux_3936 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3937;
  function [0:0] mux_3937(input [0:0] sel);
    case (sel) 0: mux_3937 = 1'h0; 1: mux_3937 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3938;
  wire [0:0] v_3939;
  wire [0:0] v_3940;
  wire [0:0] v_3941;
  wire [0:0] v_3942;
  wire [0:0] v_3943;
  function [0:0] mux_3943(input [0:0] sel);
    case (sel) 0: mux_3943 = 1'h0; 1: mux_3943 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3944;
  wire [0:0] v_3945;
  function [0:0] mux_3945(input [0:0] sel);
    case (sel) 0: mux_3945 = 1'h0; 1: mux_3945 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3946;
  wire [0:0] v_3947;
  wire [0:0] v_3948;
  wire [0:0] v_3949;
  function [0:0] mux_3949(input [0:0] sel);
    case (sel) 0: mux_3949 = 1'h0; 1: mux_3949 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3950;
  function [0:0] mux_3950(input [0:0] sel);
    case (sel) 0: mux_3950 = 1'h0; 1: mux_3950 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_3951 = 1'h0;
  wire [0:0] v_3952;
  wire [0:0] v_3953;
  wire [0:0] act_3954;
  wire [0:0] v_3955;
  wire [0:0] v_3956;
  wire [0:0] v_3957;
  reg [0:0] v_3958 = 1'h0;
  wire [0:0] v_3959;
  wire [0:0] v_3960;
  wire [0:0] act_3961;
  wire [0:0] v_3962;
  wire [0:0] v_3963;
  wire [0:0] v_3964;
  reg [0:0] v_3965 = 1'h0;
  wire [0:0] v_3966;
  wire [0:0] v_3967;
  wire [0:0] act_3968;
  wire [0:0] v_3969;
  wire [0:0] v_3970;
  wire [0:0] v_3971;
  reg [0:0] v_3972 = 1'h0;
  wire [0:0] v_3973;
  wire [0:0] v_3974;
  wire [0:0] act_3975;
  wire [0:0] v_3976;
  wire [0:0] v_3977;
  wire [0:0] v_3978;
  reg [0:0] v_3979 = 1'h0;
  wire [0:0] v_3980;
  wire [0:0] v_3981;
  wire [0:0] act_3982;
  wire [0:0] v_3983;
  wire [0:0] v_3984;
  wire [0:0] v_3985;
  reg [0:0] v_3986 = 1'h0;
  wire [0:0] v_3987;
  wire [0:0] v_3988;
  wire [0:0] act_3989;
  wire [0:0] v_3990;
  wire [0:0] v_3991;
  wire [0:0] v_3992;
  wire [0:0] v_3993;
  wire [0:0] v_3994;
  wire [0:0] v_3995;
  function [0:0] mux_3995(input [0:0] sel);
    case (sel) 0: mux_3995 = 1'h0; 1: mux_3995 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_3996;
  wire [0:0] v_3997;
  function [0:0] mux_3997(input [0:0] sel);
    case (sel) 0: mux_3997 = 1'h0; 1: mux_3997 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_3998;
  wire [0:0] v_3999;
  wire [0:0] v_4000;
  wire [0:0] v_4001;
  function [0:0] mux_4001(input [0:0] sel);
    case (sel) 0: mux_4001 = 1'h0; 1: mux_4001 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4002;
  function [0:0] mux_4002(input [0:0] sel);
    case (sel) 0: mux_4002 = 1'h0; 1: mux_4002 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4003 = 1'h0;
  wire [0:0] v_4004;
  wire [0:0] v_4005;
  wire [0:0] act_4006;
  wire [0:0] v_4007;
  wire [0:0] v_4008;
  wire [0:0] v_4009;
  wire [0:0] v_4010;
  wire [0:0] v_4011;
  wire [0:0] v_4012;
  function [0:0] mux_4012(input [0:0] sel);
    case (sel) 0: mux_4012 = 1'h0; 1: mux_4012 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4013;
  function [0:0] mux_4013(input [0:0] sel);
    case (sel) 0: mux_4013 = 1'h0; 1: mux_4013 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4014;
  wire [0:0] v_4015;
  wire [0:0] v_4016;
  wire [0:0] v_4017;
  function [0:0] mux_4017(input [0:0] sel);
    case (sel) 0: mux_4017 = 1'h0; 1: mux_4017 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4018;
  function [0:0] mux_4018(input [0:0] sel);
    case (sel) 0: mux_4018 = 1'h0; 1: mux_4018 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4019;
  wire [0:0] v_4020;
  wire [0:0] v_4021;
  wire [0:0] v_4022;
  wire [0:0] v_4023;
  wire [0:0] v_4024;
  function [0:0] mux_4024(input [0:0] sel);
    case (sel) 0: mux_4024 = 1'h0; 1: mux_4024 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4025;
  wire [0:0] v_4026;
  function [0:0] mux_4026(input [0:0] sel);
    case (sel) 0: mux_4026 = 1'h0; 1: mux_4026 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4027;
  wire [0:0] v_4028;
  wire [0:0] v_4029;
  wire [0:0] v_4030;
  function [0:0] mux_4030(input [0:0] sel);
    case (sel) 0: mux_4030 = 1'h0; 1: mux_4030 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4031;
  function [0:0] mux_4031(input [0:0] sel);
    case (sel) 0: mux_4031 = 1'h0; 1: mux_4031 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4032 = 1'h0;
  wire [0:0] v_4033;
  wire [0:0] v_4034;
  wire [0:0] act_4035;
  wire [0:0] v_4036;
  wire [0:0] v_4037;
  wire [0:0] v_4038;
  reg [0:0] v_4039 = 1'h0;
  wire [0:0] v_4040;
  wire [0:0] v_4041;
  wire [0:0] act_4042;
  wire [0:0] v_4043;
  wire [0:0] v_4044;
  wire [0:0] v_4045;
  wire [0:0] v_4046;
  wire [0:0] v_4047;
  wire [0:0] v_4048;
  function [0:0] mux_4048(input [0:0] sel);
    case (sel) 0: mux_4048 = 1'h0; 1: mux_4048 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4049;
  wire [0:0] v_4050;
  function [0:0] mux_4050(input [0:0] sel);
    case (sel) 0: mux_4050 = 1'h0; 1: mux_4050 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4051;
  wire [0:0] v_4052;
  wire [0:0] v_4053;
  wire [0:0] v_4054;
  function [0:0] mux_4054(input [0:0] sel);
    case (sel) 0: mux_4054 = 1'h0; 1: mux_4054 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4055;
  function [0:0] mux_4055(input [0:0] sel);
    case (sel) 0: mux_4055 = 1'h0; 1: mux_4055 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4056 = 1'h0;
  wire [0:0] v_4057;
  wire [0:0] v_4058;
  wire [0:0] act_4059;
  wire [0:0] v_4060;
  wire [0:0] v_4061;
  wire [0:0] v_4062;
  wire [0:0] v_4063;
  wire [0:0] v_4064;
  wire [0:0] v_4065;
  function [0:0] mux_4065(input [0:0] sel);
    case (sel) 0: mux_4065 = 1'h0; 1: mux_4065 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4066;
  function [0:0] mux_4066(input [0:0] sel);
    case (sel) 0: mux_4066 = 1'h0; 1: mux_4066 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4067;
  wire [0:0] v_4068;
  wire [0:0] v_4069;
  wire [0:0] v_4070;
  function [0:0] mux_4070(input [0:0] sel);
    case (sel) 0: mux_4070 = 1'h0; 1: mux_4070 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4071;
  function [0:0] mux_4071(input [0:0] sel);
    case (sel) 0: mux_4071 = 1'h0; 1: mux_4071 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4072;
  wire [0:0] v_4073;
  wire [0:0] v_4074;
  wire [0:0] v_4075;
  wire [0:0] v_4076;
  wire [0:0] v_4077;
  function [0:0] mux_4077(input [0:0] sel);
    case (sel) 0: mux_4077 = 1'h0; 1: mux_4077 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4078;
  function [0:0] mux_4078(input [0:0] sel);
    case (sel) 0: mux_4078 = 1'h0; 1: mux_4078 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4079;
  wire [0:0] v_4080;
  wire [0:0] v_4081;
  wire [0:0] v_4082;
  function [0:0] mux_4082(input [0:0] sel);
    case (sel) 0: mux_4082 = 1'h0; 1: mux_4082 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4083;
  function [0:0] mux_4083(input [0:0] sel);
    case (sel) 0: mux_4083 = 1'h0; 1: mux_4083 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4084;
  wire [0:0] v_4085;
  wire [0:0] v_4086;
  wire [0:0] v_4087;
  wire [0:0] v_4088;
  wire [0:0] v_4089;
  function [0:0] mux_4089(input [0:0] sel);
    case (sel) 0: mux_4089 = 1'h0; 1: mux_4089 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4090;
  wire [0:0] v_4091;
  function [0:0] mux_4091(input [0:0] sel);
    case (sel) 0: mux_4091 = 1'h0; 1: mux_4091 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4092;
  wire [0:0] v_4093;
  wire [0:0] v_4094;
  wire [0:0] v_4095;
  function [0:0] mux_4095(input [0:0] sel);
    case (sel) 0: mux_4095 = 1'h0; 1: mux_4095 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4096;
  function [0:0] mux_4096(input [0:0] sel);
    case (sel) 0: mux_4096 = 1'h0; 1: mux_4096 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4097 = 1'h0;
  wire [0:0] v_4098;
  wire [0:0] v_4099;
  wire [0:0] act_4100;
  wire [0:0] v_4101;
  wire [0:0] v_4102;
  wire [0:0] v_4103;
  reg [0:0] v_4104 = 1'h0;
  wire [0:0] v_4105;
  wire [0:0] v_4106;
  wire [0:0] act_4107;
  wire [0:0] v_4108;
  wire [0:0] v_4109;
  wire [0:0] v_4110;
  reg [0:0] v_4111 = 1'h0;
  wire [0:0] v_4112;
  wire [0:0] v_4113;
  wire [0:0] act_4114;
  wire [0:0] v_4115;
  wire [0:0] v_4116;
  wire [0:0] v_4117;
  wire [0:0] v_4118;
  wire [0:0] v_4119;
  wire [0:0] v_4120;
  function [0:0] mux_4120(input [0:0] sel);
    case (sel) 0: mux_4120 = 1'h0; 1: mux_4120 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4121;
  wire [0:0] v_4122;
  function [0:0] mux_4122(input [0:0] sel);
    case (sel) 0: mux_4122 = 1'h0; 1: mux_4122 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4123;
  wire [0:0] v_4124;
  wire [0:0] v_4125;
  wire [0:0] v_4126;
  function [0:0] mux_4126(input [0:0] sel);
    case (sel) 0: mux_4126 = 1'h0; 1: mux_4126 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4127;
  function [0:0] mux_4127(input [0:0] sel);
    case (sel) 0: mux_4127 = 1'h0; 1: mux_4127 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4128 = 1'h0;
  wire [0:0] v_4129;
  wire [0:0] v_4130;
  wire [0:0] act_4131;
  wire [0:0] v_4132;
  wire [0:0] v_4133;
  wire [0:0] v_4134;
  wire [0:0] v_4135;
  wire [0:0] v_4136;
  wire [0:0] v_4137;
  function [0:0] mux_4137(input [0:0] sel);
    case (sel) 0: mux_4137 = 1'h0; 1: mux_4137 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4138;
  function [0:0] mux_4138(input [0:0] sel);
    case (sel) 0: mux_4138 = 1'h0; 1: mux_4138 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4139;
  wire [0:0] v_4140;
  wire [0:0] v_4141;
  wire [0:0] v_4142;
  function [0:0] mux_4142(input [0:0] sel);
    case (sel) 0: mux_4142 = 1'h0; 1: mux_4142 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4143;
  function [0:0] mux_4143(input [0:0] sel);
    case (sel) 0: mux_4143 = 1'h0; 1: mux_4143 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4144;
  wire [0:0] v_4145;
  wire [0:0] v_4146;
  wire [0:0] v_4147;
  wire [0:0] v_4148;
  wire [0:0] v_4149;
  function [0:0] mux_4149(input [0:0] sel);
    case (sel) 0: mux_4149 = 1'h0; 1: mux_4149 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4150;
  wire [0:0] v_4151;
  function [0:0] mux_4151(input [0:0] sel);
    case (sel) 0: mux_4151 = 1'h0; 1: mux_4151 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4152;
  wire [0:0] v_4153;
  wire [0:0] v_4154;
  wire [0:0] v_4155;
  function [0:0] mux_4155(input [0:0] sel);
    case (sel) 0: mux_4155 = 1'h0; 1: mux_4155 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4156;
  function [0:0] mux_4156(input [0:0] sel);
    case (sel) 0: mux_4156 = 1'h0; 1: mux_4156 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4157 = 1'h0;
  wire [0:0] v_4158;
  wire [0:0] v_4159;
  wire [0:0] act_4160;
  wire [0:0] v_4161;
  wire [0:0] v_4162;
  wire [0:0] v_4163;
  reg [0:0] v_4164 = 1'h0;
  wire [0:0] v_4165;
  wire [0:0] v_4166;
  wire [0:0] act_4167;
  wire [0:0] v_4168;
  wire [0:0] v_4169;
  wire [0:0] v_4170;
  wire [0:0] v_4171;
  wire [0:0] v_4172;
  wire [0:0] v_4173;
  function [0:0] mux_4173(input [0:0] sel);
    case (sel) 0: mux_4173 = 1'h0; 1: mux_4173 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4174;
  wire [0:0] v_4175;
  function [0:0] mux_4175(input [0:0] sel);
    case (sel) 0: mux_4175 = 1'h0; 1: mux_4175 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4176;
  wire [0:0] v_4177;
  wire [0:0] v_4178;
  wire [0:0] v_4179;
  function [0:0] mux_4179(input [0:0] sel);
    case (sel) 0: mux_4179 = 1'h0; 1: mux_4179 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4180;
  function [0:0] mux_4180(input [0:0] sel);
    case (sel) 0: mux_4180 = 1'h0; 1: mux_4180 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4181 = 1'h0;
  wire [0:0] v_4182;
  wire [0:0] v_4183;
  wire [0:0] act_4184;
  wire [0:0] v_4185;
  wire [0:0] v_4186;
  wire [0:0] v_4187;
  wire [0:0] v_4188;
  wire [0:0] v_4189;
  wire [0:0] v_4190;
  function [0:0] mux_4190(input [0:0] sel);
    case (sel) 0: mux_4190 = 1'h0; 1: mux_4190 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4191;
  function [0:0] mux_4191(input [0:0] sel);
    case (sel) 0: mux_4191 = 1'h0; 1: mux_4191 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4192;
  wire [0:0] v_4193;
  wire [0:0] v_4194;
  wire [0:0] v_4195;
  function [0:0] mux_4195(input [0:0] sel);
    case (sel) 0: mux_4195 = 1'h0; 1: mux_4195 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4196;
  function [0:0] mux_4196(input [0:0] sel);
    case (sel) 0: mux_4196 = 1'h0; 1: mux_4196 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4197;
  wire [0:0] v_4198;
  wire [0:0] v_4199;
  wire [0:0] v_4200;
  wire [0:0] v_4201;
  wire [0:0] v_4202;
  function [0:0] mux_4202(input [0:0] sel);
    case (sel) 0: mux_4202 = 1'h0; 1: mux_4202 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4203;
  function [0:0] mux_4203(input [0:0] sel);
    case (sel) 0: mux_4203 = 1'h0; 1: mux_4203 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4204;
  wire [0:0] v_4205;
  wire [0:0] v_4206;
  wire [0:0] v_4207;
  function [0:0] mux_4207(input [0:0] sel);
    case (sel) 0: mux_4207 = 1'h0; 1: mux_4207 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4208;
  function [0:0] mux_4208(input [0:0] sel);
    case (sel) 0: mux_4208 = 1'h0; 1: mux_4208 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4209;
  wire [0:0] v_4210;
  wire [0:0] v_4211;
  wire [0:0] v_4212;
  wire [0:0] v_4213;
  wire [0:0] v_4214;
  function [0:0] mux_4214(input [0:0] sel);
    case (sel) 0: mux_4214 = 1'h0; 1: mux_4214 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4215;
  function [0:0] mux_4215(input [0:0] sel);
    case (sel) 0: mux_4215 = 1'h0; 1: mux_4215 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4216;
  wire [0:0] v_4217;
  wire [0:0] v_4218;
  wire [0:0] v_4219;
  function [0:0] mux_4219(input [0:0] sel);
    case (sel) 0: mux_4219 = 1'h0; 1: mux_4219 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4220;
  function [0:0] mux_4220(input [0:0] sel);
    case (sel) 0: mux_4220 = 1'h0; 1: mux_4220 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4221;
  wire [0:0] v_4222;
  wire [0:0] v_4223;
  wire [0:0] v_4224;
  wire [0:0] v_4225;
  wire [0:0] v_4226;
  function [0:0] mux_4226(input [0:0] sel);
    case (sel) 0: mux_4226 = 1'h0; 1: mux_4226 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4227;
  wire [0:0] v_4228;
  function [0:0] mux_4228(input [0:0] sel);
    case (sel) 0: mux_4228 = 1'h0; 1: mux_4228 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4229;
  wire [0:0] v_4230;
  wire [0:0] v_4231;
  wire [0:0] v_4232;
  function [0:0] mux_4232(input [0:0] sel);
    case (sel) 0: mux_4232 = 1'h0; 1: mux_4232 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4233;
  function [0:0] mux_4233(input [0:0] sel);
    case (sel) 0: mux_4233 = 1'h0; 1: mux_4233 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4234 = 1'h0;
  wire [0:0] v_4235;
  wire [0:0] v_4236;
  wire [0:0] act_4237;
  wire [0:0] v_4238;
  wire [0:0] v_4239;
  wire [0:0] v_4240;
  reg [0:0] v_4241 = 1'h0;
  wire [0:0] v_4242;
  wire [0:0] v_4243;
  wire [0:0] act_4244;
  wire [0:0] v_4245;
  wire [0:0] v_4246;
  wire [0:0] v_4247;
  reg [0:0] v_4248 = 1'h0;
  wire [0:0] v_4249;
  wire [0:0] v_4250;
  wire [0:0] act_4251;
  wire [0:0] v_4252;
  wire [0:0] v_4253;
  wire [0:0] v_4254;
  reg [0:0] v_4255 = 1'h0;
  wire [0:0] v_4256;
  wire [0:0] v_4257;
  wire [0:0] act_4258;
  wire [0:0] v_4259;
  wire [0:0] v_4260;
  wire [0:0] v_4261;
  wire [0:0] v_4262;
  wire [0:0] v_4263;
  wire [0:0] v_4264;
  function [0:0] mux_4264(input [0:0] sel);
    case (sel) 0: mux_4264 = 1'h0; 1: mux_4264 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4265;
  wire [0:0] v_4266;
  function [0:0] mux_4266(input [0:0] sel);
    case (sel) 0: mux_4266 = 1'h0; 1: mux_4266 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4267;
  wire [0:0] v_4268;
  wire [0:0] v_4269;
  wire [0:0] v_4270;
  function [0:0] mux_4270(input [0:0] sel);
    case (sel) 0: mux_4270 = 1'h0; 1: mux_4270 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4271;
  function [0:0] mux_4271(input [0:0] sel);
    case (sel) 0: mux_4271 = 1'h0; 1: mux_4271 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4272 = 1'h0;
  wire [0:0] v_4273;
  wire [0:0] v_4274;
  wire [0:0] act_4275;
  wire [0:0] v_4276;
  wire [0:0] v_4277;
  wire [0:0] v_4278;
  wire [0:0] v_4279;
  wire [0:0] v_4280;
  wire [0:0] v_4281;
  function [0:0] mux_4281(input [0:0] sel);
    case (sel) 0: mux_4281 = 1'h0; 1: mux_4281 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4282;
  function [0:0] mux_4282(input [0:0] sel);
    case (sel) 0: mux_4282 = 1'h0; 1: mux_4282 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4283;
  wire [0:0] v_4284;
  wire [0:0] v_4285;
  wire [0:0] v_4286;
  function [0:0] mux_4286(input [0:0] sel);
    case (sel) 0: mux_4286 = 1'h0; 1: mux_4286 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4287;
  function [0:0] mux_4287(input [0:0] sel);
    case (sel) 0: mux_4287 = 1'h0; 1: mux_4287 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4288;
  wire [0:0] v_4289;
  wire [0:0] v_4290;
  wire [0:0] v_4291;
  wire [0:0] v_4292;
  wire [0:0] v_4293;
  function [0:0] mux_4293(input [0:0] sel);
    case (sel) 0: mux_4293 = 1'h0; 1: mux_4293 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4294;
  wire [0:0] v_4295;
  function [0:0] mux_4295(input [0:0] sel);
    case (sel) 0: mux_4295 = 1'h0; 1: mux_4295 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4296;
  wire [0:0] v_4297;
  wire [0:0] v_4298;
  wire [0:0] v_4299;
  function [0:0] mux_4299(input [0:0] sel);
    case (sel) 0: mux_4299 = 1'h0; 1: mux_4299 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4300;
  function [0:0] mux_4300(input [0:0] sel);
    case (sel) 0: mux_4300 = 1'h0; 1: mux_4300 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4301 = 1'h0;
  wire [0:0] v_4302;
  wire [0:0] v_4303;
  wire [0:0] act_4304;
  wire [0:0] v_4305;
  wire [0:0] v_4306;
  wire [0:0] v_4307;
  reg [0:0] v_4308 = 1'h0;
  wire [0:0] v_4309;
  wire [0:0] v_4310;
  wire [0:0] act_4311;
  wire [0:0] v_4312;
  wire [0:0] v_4313;
  wire [0:0] v_4314;
  wire [0:0] v_4315;
  wire [0:0] v_4316;
  wire [0:0] v_4317;
  function [0:0] mux_4317(input [0:0] sel);
    case (sel) 0: mux_4317 = 1'h0; 1: mux_4317 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4318;
  wire [0:0] v_4319;
  function [0:0] mux_4319(input [0:0] sel);
    case (sel) 0: mux_4319 = 1'h0; 1: mux_4319 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4320;
  wire [0:0] v_4321;
  wire [0:0] v_4322;
  wire [0:0] v_4323;
  function [0:0] mux_4323(input [0:0] sel);
    case (sel) 0: mux_4323 = 1'h0; 1: mux_4323 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4324;
  function [0:0] mux_4324(input [0:0] sel);
    case (sel) 0: mux_4324 = 1'h0; 1: mux_4324 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4325 = 1'h0;
  wire [0:0] v_4326;
  wire [0:0] v_4327;
  wire [0:0] act_4328;
  wire [0:0] v_4329;
  wire [0:0] v_4330;
  wire [0:0] v_4331;
  wire [0:0] v_4332;
  wire [0:0] v_4333;
  wire [0:0] v_4334;
  function [0:0] mux_4334(input [0:0] sel);
    case (sel) 0: mux_4334 = 1'h0; 1: mux_4334 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4335;
  function [0:0] mux_4335(input [0:0] sel);
    case (sel) 0: mux_4335 = 1'h0; 1: mux_4335 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4336;
  wire [0:0] v_4337;
  wire [0:0] v_4338;
  wire [0:0] v_4339;
  function [0:0] mux_4339(input [0:0] sel);
    case (sel) 0: mux_4339 = 1'h0; 1: mux_4339 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4340;
  function [0:0] mux_4340(input [0:0] sel);
    case (sel) 0: mux_4340 = 1'h0; 1: mux_4340 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4341;
  wire [0:0] v_4342;
  wire [0:0] v_4343;
  wire [0:0] v_4344;
  wire [0:0] v_4345;
  wire [0:0] v_4346;
  function [0:0] mux_4346(input [0:0] sel);
    case (sel) 0: mux_4346 = 1'h0; 1: mux_4346 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4347;
  function [0:0] mux_4347(input [0:0] sel);
    case (sel) 0: mux_4347 = 1'h0; 1: mux_4347 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4348;
  wire [0:0] v_4349;
  wire [0:0] v_4350;
  wire [0:0] v_4351;
  function [0:0] mux_4351(input [0:0] sel);
    case (sel) 0: mux_4351 = 1'h0; 1: mux_4351 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4352;
  function [0:0] mux_4352(input [0:0] sel);
    case (sel) 0: mux_4352 = 1'h0; 1: mux_4352 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4353;
  wire [0:0] v_4354;
  wire [0:0] v_4355;
  wire [0:0] v_4356;
  wire [0:0] v_4357;
  wire [0:0] v_4358;
  function [0:0] mux_4358(input [0:0] sel);
    case (sel) 0: mux_4358 = 1'h0; 1: mux_4358 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4359;
  wire [0:0] v_4360;
  function [0:0] mux_4360(input [0:0] sel);
    case (sel) 0: mux_4360 = 1'h0; 1: mux_4360 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4361;
  wire [0:0] v_4362;
  wire [0:0] v_4363;
  wire [0:0] v_4364;
  function [0:0] mux_4364(input [0:0] sel);
    case (sel) 0: mux_4364 = 1'h0; 1: mux_4364 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4365;
  function [0:0] mux_4365(input [0:0] sel);
    case (sel) 0: mux_4365 = 1'h0; 1: mux_4365 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4366 = 1'h0;
  wire [0:0] v_4367;
  wire [0:0] v_4368;
  wire [0:0] act_4369;
  wire [0:0] v_4370;
  wire [0:0] v_4371;
  wire [0:0] v_4372;
  reg [0:0] v_4373 = 1'h0;
  wire [0:0] v_4374;
  wire [0:0] v_4375;
  wire [0:0] act_4376;
  wire [0:0] v_4377;
  wire [0:0] v_4378;
  wire [0:0] v_4379;
  reg [0:0] v_4380 = 1'h0;
  wire [0:0] v_4381;
  wire [0:0] v_4382;
  wire [0:0] act_4383;
  wire [0:0] v_4384;
  wire [0:0] v_4385;
  wire [0:0] v_4386;
  wire [0:0] v_4387;
  wire [0:0] v_4388;
  wire [0:0] v_4389;
  function [0:0] mux_4389(input [0:0] sel);
    case (sel) 0: mux_4389 = 1'h0; 1: mux_4389 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4390;
  wire [0:0] v_4391;
  function [0:0] mux_4391(input [0:0] sel);
    case (sel) 0: mux_4391 = 1'h0; 1: mux_4391 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4392;
  wire [0:0] v_4393;
  wire [0:0] v_4394;
  wire [0:0] v_4395;
  function [0:0] mux_4395(input [0:0] sel);
    case (sel) 0: mux_4395 = 1'h0; 1: mux_4395 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4396;
  function [0:0] mux_4396(input [0:0] sel);
    case (sel) 0: mux_4396 = 1'h0; 1: mux_4396 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4397 = 1'h0;
  wire [0:0] v_4398;
  wire [0:0] v_4399;
  wire [0:0] act_4400;
  wire [0:0] v_4401;
  wire [0:0] v_4402;
  wire [0:0] v_4403;
  wire [0:0] v_4404;
  wire [0:0] v_4405;
  wire [0:0] v_4406;
  function [0:0] mux_4406(input [0:0] sel);
    case (sel) 0: mux_4406 = 1'h0; 1: mux_4406 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4407;
  function [0:0] mux_4407(input [0:0] sel);
    case (sel) 0: mux_4407 = 1'h0; 1: mux_4407 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4408;
  wire [0:0] v_4409;
  wire [0:0] v_4410;
  wire [0:0] v_4411;
  function [0:0] mux_4411(input [0:0] sel);
    case (sel) 0: mux_4411 = 1'h0; 1: mux_4411 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4412;
  function [0:0] mux_4412(input [0:0] sel);
    case (sel) 0: mux_4412 = 1'h0; 1: mux_4412 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4413;
  wire [0:0] v_4414;
  wire [0:0] v_4415;
  wire [0:0] v_4416;
  wire [0:0] v_4417;
  wire [0:0] v_4418;
  function [0:0] mux_4418(input [0:0] sel);
    case (sel) 0: mux_4418 = 1'h0; 1: mux_4418 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4419;
  wire [0:0] v_4420;
  function [0:0] mux_4420(input [0:0] sel);
    case (sel) 0: mux_4420 = 1'h0; 1: mux_4420 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4421;
  wire [0:0] v_4422;
  wire [0:0] v_4423;
  wire [0:0] v_4424;
  function [0:0] mux_4424(input [0:0] sel);
    case (sel) 0: mux_4424 = 1'h0; 1: mux_4424 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4425;
  function [0:0] mux_4425(input [0:0] sel);
    case (sel) 0: mux_4425 = 1'h0; 1: mux_4425 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4426 = 1'h0;
  wire [0:0] v_4427;
  wire [0:0] v_4428;
  wire [0:0] act_4429;
  wire [0:0] v_4430;
  wire [0:0] v_4431;
  wire [0:0] v_4432;
  reg [0:0] v_4433 = 1'h0;
  wire [0:0] v_4434;
  wire [0:0] v_4435;
  wire [0:0] act_4436;
  wire [0:0] v_4437;
  wire [0:0] v_4438;
  wire [0:0] v_4439;
  wire [0:0] v_4440;
  wire [0:0] v_4441;
  wire [0:0] v_4442;
  function [0:0] mux_4442(input [0:0] sel);
    case (sel) 0: mux_4442 = 1'h0; 1: mux_4442 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4443;
  wire [0:0] v_4444;
  function [0:0] mux_4444(input [0:0] sel);
    case (sel) 0: mux_4444 = 1'h0; 1: mux_4444 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4445;
  wire [0:0] v_4446;
  wire [0:0] v_4447;
  wire [0:0] v_4448;
  function [0:0] mux_4448(input [0:0] sel);
    case (sel) 0: mux_4448 = 1'h0; 1: mux_4448 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4449;
  function [0:0] mux_4449(input [0:0] sel);
    case (sel) 0: mux_4449 = 1'h0; 1: mux_4449 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4450 = 1'h0;
  wire [0:0] v_4451;
  wire [0:0] v_4452;
  wire [0:0] act_4453;
  wire [0:0] v_4454;
  wire [0:0] v_4455;
  wire [0:0] v_4456;
  wire [0:0] v_4457;
  wire [0:0] v_4458;
  wire [0:0] v_4459;
  function [0:0] mux_4459(input [0:0] sel);
    case (sel) 0: mux_4459 = 1'h0; 1: mux_4459 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4460;
  function [0:0] mux_4460(input [0:0] sel);
    case (sel) 0: mux_4460 = 1'h0; 1: mux_4460 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4461;
  wire [0:0] v_4462;
  wire [0:0] v_4463;
  wire [0:0] v_4464;
  function [0:0] mux_4464(input [0:0] sel);
    case (sel) 0: mux_4464 = 1'h0; 1: mux_4464 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4465;
  function [0:0] mux_4465(input [0:0] sel);
    case (sel) 0: mux_4465 = 1'h0; 1: mux_4465 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4466;
  wire [0:0] v_4467;
  wire [0:0] v_4468;
  wire [0:0] v_4469;
  wire [0:0] v_4470;
  wire [0:0] v_4471;
  function [0:0] mux_4471(input [0:0] sel);
    case (sel) 0: mux_4471 = 1'h0; 1: mux_4471 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4472;
  function [0:0] mux_4472(input [0:0] sel);
    case (sel) 0: mux_4472 = 1'h0; 1: mux_4472 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4473;
  wire [0:0] v_4474;
  wire [0:0] v_4475;
  wire [0:0] v_4476;
  function [0:0] mux_4476(input [0:0] sel);
    case (sel) 0: mux_4476 = 1'h0; 1: mux_4476 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4477;
  function [0:0] mux_4477(input [0:0] sel);
    case (sel) 0: mux_4477 = 1'h0; 1: mux_4477 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4478;
  wire [0:0] v_4479;
  wire [0:0] v_4480;
  wire [0:0] v_4481;
  wire [0:0] v_4482;
  wire [0:0] v_4483;
  function [0:0] mux_4483(input [0:0] sel);
    case (sel) 0: mux_4483 = 1'h0; 1: mux_4483 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4484;
  function [0:0] mux_4484(input [0:0] sel);
    case (sel) 0: mux_4484 = 1'h0; 1: mux_4484 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4485;
  wire [0:0] v_4486;
  wire [0:0] v_4487;
  wire [0:0] v_4488;
  function [0:0] mux_4488(input [0:0] sel);
    case (sel) 0: mux_4488 = 1'h0; 1: mux_4488 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4489;
  function [0:0] mux_4489(input [0:0] sel);
    case (sel) 0: mux_4489 = 1'h0; 1: mux_4489 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4490;
  wire [0:0] v_4491;
  wire [0:0] v_4492;
  wire [0:0] v_4493;
  wire [0:0] v_4494;
  wire [0:0] v_4495;
  function [0:0] mux_4495(input [0:0] sel);
    case (sel) 0: mux_4495 = 1'h0; 1: mux_4495 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4496;
  function [0:0] mux_4496(input [0:0] sel);
    case (sel) 0: mux_4496 = 1'h0; 1: mux_4496 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4497;
  wire [0:0] v_4498;
  wire [0:0] v_4499;
  wire [0:0] v_4500;
  function [0:0] mux_4500(input [0:0] sel);
    case (sel) 0: mux_4500 = 1'h0; 1: mux_4500 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4501;
  function [0:0] mux_4501(input [0:0] sel);
    case (sel) 0: mux_4501 = 1'h0; 1: mux_4501 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4502;
  wire [0:0] v_4503;
  wire [0:0] v_4504;
  wire [0:0] v_4505;
  wire [0:0] v_4506;
  wire [0:0] v_4507;
  function [0:0] mux_4507(input [0:0] sel);
    case (sel) 0: mux_4507 = 1'h0; 1: mux_4507 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4508;
  wire [0:0] v_4509;
  function [0:0] mux_4509(input [0:0] sel);
    case (sel) 0: mux_4509 = 1'h0; 1: mux_4509 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4510;
  wire [0:0] v_4511;
  wire [0:0] v_4512;
  wire [0:0] v_4513;
  function [0:0] mux_4513(input [0:0] sel);
    case (sel) 0: mux_4513 = 1'h0; 1: mux_4513 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4514;
  function [0:0] mux_4514(input [0:0] sel);
    case (sel) 0: mux_4514 = 1'h0; 1: mux_4514 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4515 = 1'h0;
  wire [0:0] v_4516;
  wire [0:0] v_4517;
  wire [0:0] act_4518;
  wire [0:0] v_4519;
  wire [0:0] v_4520;
  wire [0:0] v_4521;
  reg [0:0] v_4522 = 1'h0;
  wire [0:0] v_4523;
  wire [0:0] v_4524;
  wire [0:0] act_4525;
  wire [0:0] v_4526;
  wire [0:0] v_4527;
  wire [0:0] v_4528;
  reg [0:0] v_4529 = 1'h0;
  wire [0:0] v_4530;
  wire [0:0] v_4531;
  wire [0:0] act_4532;
  wire [0:0] v_4533;
  wire [0:0] v_4534;
  wire [0:0] v_4535;
  reg [0:0] v_4536 = 1'h0;
  wire [0:0] v_4537;
  wire [0:0] v_4538;
  wire [0:0] act_4539;
  wire [0:0] v_4540;
  wire [0:0] v_4541;
  wire [0:0] v_4542;
  reg [0:0] v_4543 = 1'h0;
  wire [0:0] v_4544;
  wire [0:0] v_4545;
  wire [0:0] act_4546;
  wire [0:0] v_4547;
  wire [0:0] v_4548;
  wire [0:0] v_4549;
  wire [0:0] v_4550;
  wire [0:0] v_4551;
  wire [0:0] v_4552;
  function [0:0] mux_4552(input [0:0] sel);
    case (sel) 0: mux_4552 = 1'h0; 1: mux_4552 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4553;
  wire [0:0] v_4554;
  function [0:0] mux_4554(input [0:0] sel);
    case (sel) 0: mux_4554 = 1'h0; 1: mux_4554 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4555;
  wire [0:0] v_4556;
  wire [0:0] v_4557;
  wire [0:0] v_4558;
  function [0:0] mux_4558(input [0:0] sel);
    case (sel) 0: mux_4558 = 1'h0; 1: mux_4558 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4559;
  function [0:0] mux_4559(input [0:0] sel);
    case (sel) 0: mux_4559 = 1'h0; 1: mux_4559 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4560 = 1'h0;
  wire [0:0] v_4561;
  wire [0:0] v_4562;
  wire [0:0] act_4563;
  wire [0:0] v_4564;
  wire [0:0] v_4565;
  wire [0:0] v_4566;
  wire [0:0] v_4567;
  wire [0:0] v_4568;
  wire [0:0] v_4569;
  function [0:0] mux_4569(input [0:0] sel);
    case (sel) 0: mux_4569 = 1'h0; 1: mux_4569 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4570;
  function [0:0] mux_4570(input [0:0] sel);
    case (sel) 0: mux_4570 = 1'h0; 1: mux_4570 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4571;
  wire [0:0] v_4572;
  wire [0:0] v_4573;
  wire [0:0] v_4574;
  function [0:0] mux_4574(input [0:0] sel);
    case (sel) 0: mux_4574 = 1'h0; 1: mux_4574 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4575;
  function [0:0] mux_4575(input [0:0] sel);
    case (sel) 0: mux_4575 = 1'h0; 1: mux_4575 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4576;
  wire [0:0] v_4577;
  wire [0:0] v_4578;
  wire [0:0] v_4579;
  wire [0:0] v_4580;
  wire [0:0] v_4581;
  function [0:0] mux_4581(input [0:0] sel);
    case (sel) 0: mux_4581 = 1'h0; 1: mux_4581 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4582;
  wire [0:0] v_4583;
  function [0:0] mux_4583(input [0:0] sel);
    case (sel) 0: mux_4583 = 1'h0; 1: mux_4583 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4584;
  wire [0:0] v_4585;
  wire [0:0] v_4586;
  wire [0:0] v_4587;
  function [0:0] mux_4587(input [0:0] sel);
    case (sel) 0: mux_4587 = 1'h0; 1: mux_4587 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4588;
  function [0:0] mux_4588(input [0:0] sel);
    case (sel) 0: mux_4588 = 1'h0; 1: mux_4588 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4589 = 1'h0;
  wire [0:0] v_4590;
  wire [0:0] v_4591;
  wire [0:0] act_4592;
  wire [0:0] v_4593;
  wire [0:0] v_4594;
  wire [0:0] v_4595;
  reg [0:0] v_4596 = 1'h0;
  wire [0:0] v_4597;
  wire [0:0] v_4598;
  wire [0:0] act_4599;
  wire [0:0] v_4600;
  wire [0:0] v_4601;
  wire [0:0] v_4602;
  wire [0:0] v_4603;
  wire [0:0] v_4604;
  wire [0:0] v_4605;
  function [0:0] mux_4605(input [0:0] sel);
    case (sel) 0: mux_4605 = 1'h0; 1: mux_4605 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4606;
  wire [0:0] v_4607;
  function [0:0] mux_4607(input [0:0] sel);
    case (sel) 0: mux_4607 = 1'h0; 1: mux_4607 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4608;
  wire [0:0] v_4609;
  wire [0:0] v_4610;
  wire [0:0] v_4611;
  function [0:0] mux_4611(input [0:0] sel);
    case (sel) 0: mux_4611 = 1'h0; 1: mux_4611 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4612;
  function [0:0] mux_4612(input [0:0] sel);
    case (sel) 0: mux_4612 = 1'h0; 1: mux_4612 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4613 = 1'h0;
  wire [0:0] v_4614;
  wire [0:0] v_4615;
  wire [0:0] act_4616;
  wire [0:0] v_4617;
  wire [0:0] v_4618;
  wire [0:0] v_4619;
  wire [0:0] v_4620;
  wire [0:0] v_4621;
  wire [0:0] v_4622;
  function [0:0] mux_4622(input [0:0] sel);
    case (sel) 0: mux_4622 = 1'h0; 1: mux_4622 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4623;
  function [0:0] mux_4623(input [0:0] sel);
    case (sel) 0: mux_4623 = 1'h0; 1: mux_4623 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4624;
  wire [0:0] v_4625;
  wire [0:0] v_4626;
  wire [0:0] v_4627;
  function [0:0] mux_4627(input [0:0] sel);
    case (sel) 0: mux_4627 = 1'h0; 1: mux_4627 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4628;
  function [0:0] mux_4628(input [0:0] sel);
    case (sel) 0: mux_4628 = 1'h0; 1: mux_4628 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4629;
  wire [0:0] v_4630;
  wire [0:0] v_4631;
  wire [0:0] v_4632;
  wire [0:0] v_4633;
  wire [0:0] v_4634;
  function [0:0] mux_4634(input [0:0] sel);
    case (sel) 0: mux_4634 = 1'h0; 1: mux_4634 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4635;
  function [0:0] mux_4635(input [0:0] sel);
    case (sel) 0: mux_4635 = 1'h0; 1: mux_4635 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4636;
  wire [0:0] v_4637;
  wire [0:0] v_4638;
  wire [0:0] v_4639;
  function [0:0] mux_4639(input [0:0] sel);
    case (sel) 0: mux_4639 = 1'h0; 1: mux_4639 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4640;
  function [0:0] mux_4640(input [0:0] sel);
    case (sel) 0: mux_4640 = 1'h0; 1: mux_4640 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4641;
  wire [0:0] v_4642;
  wire [0:0] v_4643;
  wire [0:0] v_4644;
  wire [0:0] v_4645;
  wire [0:0] v_4646;
  function [0:0] mux_4646(input [0:0] sel);
    case (sel) 0: mux_4646 = 1'h0; 1: mux_4646 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4647;
  wire [0:0] v_4648;
  function [0:0] mux_4648(input [0:0] sel);
    case (sel) 0: mux_4648 = 1'h0; 1: mux_4648 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4649;
  wire [0:0] v_4650;
  wire [0:0] v_4651;
  wire [0:0] v_4652;
  function [0:0] mux_4652(input [0:0] sel);
    case (sel) 0: mux_4652 = 1'h0; 1: mux_4652 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4653;
  function [0:0] mux_4653(input [0:0] sel);
    case (sel) 0: mux_4653 = 1'h0; 1: mux_4653 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4654 = 1'h0;
  wire [0:0] v_4655;
  wire [0:0] v_4656;
  wire [0:0] act_4657;
  wire [0:0] v_4658;
  wire [0:0] v_4659;
  wire [0:0] v_4660;
  reg [0:0] v_4661 = 1'h0;
  wire [0:0] v_4662;
  wire [0:0] v_4663;
  wire [0:0] act_4664;
  wire [0:0] v_4665;
  wire [0:0] v_4666;
  wire [0:0] v_4667;
  reg [0:0] v_4668 = 1'h0;
  wire [0:0] v_4669;
  wire [0:0] v_4670;
  wire [0:0] act_4671;
  wire [0:0] v_4672;
  wire [0:0] v_4673;
  wire [0:0] v_4674;
  wire [0:0] v_4675;
  wire [0:0] v_4676;
  wire [0:0] v_4677;
  function [0:0] mux_4677(input [0:0] sel);
    case (sel) 0: mux_4677 = 1'h0; 1: mux_4677 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4678;
  wire [0:0] v_4679;
  function [0:0] mux_4679(input [0:0] sel);
    case (sel) 0: mux_4679 = 1'h0; 1: mux_4679 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4680;
  wire [0:0] v_4681;
  wire [0:0] v_4682;
  wire [0:0] v_4683;
  function [0:0] mux_4683(input [0:0] sel);
    case (sel) 0: mux_4683 = 1'h0; 1: mux_4683 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4684;
  function [0:0] mux_4684(input [0:0] sel);
    case (sel) 0: mux_4684 = 1'h0; 1: mux_4684 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4685 = 1'h0;
  wire [0:0] v_4686;
  wire [0:0] v_4687;
  wire [0:0] act_4688;
  wire [0:0] v_4689;
  wire [0:0] v_4690;
  wire [0:0] v_4691;
  wire [0:0] v_4692;
  wire [0:0] v_4693;
  wire [0:0] v_4694;
  function [0:0] mux_4694(input [0:0] sel);
    case (sel) 0: mux_4694 = 1'h0; 1: mux_4694 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4695;
  function [0:0] mux_4695(input [0:0] sel);
    case (sel) 0: mux_4695 = 1'h0; 1: mux_4695 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4696;
  wire [0:0] v_4697;
  wire [0:0] v_4698;
  wire [0:0] v_4699;
  function [0:0] mux_4699(input [0:0] sel);
    case (sel) 0: mux_4699 = 1'h0; 1: mux_4699 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4700;
  function [0:0] mux_4700(input [0:0] sel);
    case (sel) 0: mux_4700 = 1'h0; 1: mux_4700 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4701;
  wire [0:0] v_4702;
  wire [0:0] v_4703;
  wire [0:0] v_4704;
  wire [0:0] v_4705;
  wire [0:0] v_4706;
  function [0:0] mux_4706(input [0:0] sel);
    case (sel) 0: mux_4706 = 1'h0; 1: mux_4706 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4707;
  wire [0:0] v_4708;
  function [0:0] mux_4708(input [0:0] sel);
    case (sel) 0: mux_4708 = 1'h0; 1: mux_4708 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4709;
  wire [0:0] v_4710;
  wire [0:0] v_4711;
  wire [0:0] v_4712;
  function [0:0] mux_4712(input [0:0] sel);
    case (sel) 0: mux_4712 = 1'h0; 1: mux_4712 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4713;
  function [0:0] mux_4713(input [0:0] sel);
    case (sel) 0: mux_4713 = 1'h0; 1: mux_4713 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4714 = 1'h0;
  wire [0:0] v_4715;
  wire [0:0] v_4716;
  wire [0:0] act_4717;
  wire [0:0] v_4718;
  wire [0:0] v_4719;
  wire [0:0] v_4720;
  reg [0:0] v_4721 = 1'h0;
  wire [0:0] v_4722;
  wire [0:0] v_4723;
  wire [0:0] act_4724;
  wire [0:0] v_4725;
  wire [0:0] v_4726;
  wire [0:0] v_4727;
  wire [0:0] v_4728;
  wire [0:0] v_4729;
  wire [0:0] v_4730;
  function [0:0] mux_4730(input [0:0] sel);
    case (sel) 0: mux_4730 = 1'h0; 1: mux_4730 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4731;
  wire [0:0] v_4732;
  function [0:0] mux_4732(input [0:0] sel);
    case (sel) 0: mux_4732 = 1'h0; 1: mux_4732 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4733;
  wire [0:0] v_4734;
  wire [0:0] v_4735;
  wire [0:0] v_4736;
  function [0:0] mux_4736(input [0:0] sel);
    case (sel) 0: mux_4736 = 1'h0; 1: mux_4736 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4737;
  function [0:0] mux_4737(input [0:0] sel);
    case (sel) 0: mux_4737 = 1'h0; 1: mux_4737 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4738 = 1'h0;
  wire [0:0] v_4739;
  wire [0:0] v_4740;
  wire [0:0] act_4741;
  wire [0:0] v_4742;
  wire [0:0] v_4743;
  wire [0:0] v_4744;
  wire [0:0] v_4745;
  wire [0:0] v_4746;
  wire [0:0] v_4747;
  function [0:0] mux_4747(input [0:0] sel);
    case (sel) 0: mux_4747 = 1'h0; 1: mux_4747 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4748;
  function [0:0] mux_4748(input [0:0] sel);
    case (sel) 0: mux_4748 = 1'h0; 1: mux_4748 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4749;
  wire [0:0] v_4750;
  wire [0:0] v_4751;
  wire [0:0] v_4752;
  function [0:0] mux_4752(input [0:0] sel);
    case (sel) 0: mux_4752 = 1'h0; 1: mux_4752 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4753;
  function [0:0] mux_4753(input [0:0] sel);
    case (sel) 0: mux_4753 = 1'h0; 1: mux_4753 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4754;
  wire [0:0] v_4755;
  wire [0:0] v_4756;
  wire [0:0] v_4757;
  wire [0:0] v_4758;
  wire [0:0] v_4759;
  function [0:0] mux_4759(input [0:0] sel);
    case (sel) 0: mux_4759 = 1'h0; 1: mux_4759 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4760;
  function [0:0] mux_4760(input [0:0] sel);
    case (sel) 0: mux_4760 = 1'h0; 1: mux_4760 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4761;
  wire [0:0] v_4762;
  wire [0:0] v_4763;
  wire [0:0] v_4764;
  function [0:0] mux_4764(input [0:0] sel);
    case (sel) 0: mux_4764 = 1'h0; 1: mux_4764 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4765;
  function [0:0] mux_4765(input [0:0] sel);
    case (sel) 0: mux_4765 = 1'h0; 1: mux_4765 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4766;
  wire [0:0] v_4767;
  wire [0:0] v_4768;
  wire [0:0] v_4769;
  wire [0:0] v_4770;
  wire [0:0] v_4771;
  function [0:0] mux_4771(input [0:0] sel);
    case (sel) 0: mux_4771 = 1'h0; 1: mux_4771 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4772;
  function [0:0] mux_4772(input [0:0] sel);
    case (sel) 0: mux_4772 = 1'h0; 1: mux_4772 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4773;
  wire [0:0] v_4774;
  wire [0:0] v_4775;
  wire [0:0] v_4776;
  function [0:0] mux_4776(input [0:0] sel);
    case (sel) 0: mux_4776 = 1'h0; 1: mux_4776 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4777;
  function [0:0] mux_4777(input [0:0] sel);
    case (sel) 0: mux_4777 = 1'h0; 1: mux_4777 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4778;
  wire [0:0] v_4779;
  wire [0:0] v_4780;
  wire [0:0] v_4781;
  wire [0:0] v_4782;
  wire [0:0] v_4783;
  function [0:0] mux_4783(input [0:0] sel);
    case (sel) 0: mux_4783 = 1'h0; 1: mux_4783 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4784;
  wire [0:0] v_4785;
  function [0:0] mux_4785(input [0:0] sel);
    case (sel) 0: mux_4785 = 1'h0; 1: mux_4785 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4786;
  wire [0:0] v_4787;
  wire [0:0] v_4788;
  wire [0:0] v_4789;
  function [0:0] mux_4789(input [0:0] sel);
    case (sel) 0: mux_4789 = 1'h0; 1: mux_4789 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4790;
  function [0:0] mux_4790(input [0:0] sel);
    case (sel) 0: mux_4790 = 1'h0; 1: mux_4790 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4791 = 1'h0;
  wire [0:0] v_4792;
  wire [0:0] v_4793;
  wire [0:0] act_4794;
  wire [0:0] v_4795;
  wire [0:0] v_4796;
  wire [0:0] v_4797;
  reg [0:0] v_4798 = 1'h0;
  wire [0:0] v_4799;
  wire [0:0] v_4800;
  wire [0:0] act_4801;
  wire [0:0] v_4802;
  wire [0:0] v_4803;
  wire [0:0] v_4804;
  reg [0:0] v_4805 = 1'h0;
  wire [0:0] v_4806;
  wire [0:0] v_4807;
  wire [0:0] act_4808;
  wire [0:0] v_4809;
  wire [0:0] v_4810;
  wire [0:0] v_4811;
  reg [0:0] v_4812 = 1'h0;
  wire [0:0] v_4813;
  wire [0:0] v_4814;
  wire [0:0] act_4815;
  wire [0:0] v_4816;
  wire [0:0] v_4817;
  wire [0:0] v_4818;
  reg [0:0] v_4819 = 1'h0;
  wire [0:0] v_4820;
  wire [0:0] v_4821;
  wire [0:0] act_4822;
  wire [0:0] v_4823;
  wire [0:0] v_4824;
  wire [0:0] v_4825;
  wire [0:0] v_4826;
  wire [0:0] v_4827;
  wire [0:0] v_4828;
  function [0:0] mux_4828(input [0:0] sel);
    case (sel) 0: mux_4828 = 1'h0; 1: mux_4828 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4829;
  wire [0:0] v_4830;
  function [0:0] mux_4830(input [0:0] sel);
    case (sel) 0: mux_4830 = 1'h0; 1: mux_4830 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4831;
  wire [0:0] v_4832;
  wire [0:0] v_4833;
  wire [0:0] v_4834;
  function [0:0] mux_4834(input [0:0] sel);
    case (sel) 0: mux_4834 = 1'h0; 1: mux_4834 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4835;
  function [0:0] mux_4835(input [0:0] sel);
    case (sel) 0: mux_4835 = 1'h0; 1: mux_4835 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4836 = 1'h0;
  wire [0:0] v_4837;
  wire [0:0] v_4838;
  wire [0:0] act_4839;
  wire [0:0] v_4840;
  wire [0:0] v_4841;
  wire [0:0] v_4842;
  wire [0:0] v_4843;
  wire [0:0] v_4844;
  wire [0:0] v_4845;
  function [0:0] mux_4845(input [0:0] sel);
    case (sel) 0: mux_4845 = 1'h0; 1: mux_4845 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4846;
  function [0:0] mux_4846(input [0:0] sel);
    case (sel) 0: mux_4846 = 1'h0; 1: mux_4846 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4847;
  wire [0:0] v_4848;
  wire [0:0] v_4849;
  wire [0:0] v_4850;
  function [0:0] mux_4850(input [0:0] sel);
    case (sel) 0: mux_4850 = 1'h0; 1: mux_4850 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4851;
  function [0:0] mux_4851(input [0:0] sel);
    case (sel) 0: mux_4851 = 1'h0; 1: mux_4851 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4852;
  wire [0:0] v_4853;
  wire [0:0] v_4854;
  wire [0:0] v_4855;
  wire [0:0] v_4856;
  wire [0:0] v_4857;
  function [0:0] mux_4857(input [0:0] sel);
    case (sel) 0: mux_4857 = 1'h0; 1: mux_4857 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4858;
  wire [0:0] v_4859;
  function [0:0] mux_4859(input [0:0] sel);
    case (sel) 0: mux_4859 = 1'h0; 1: mux_4859 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4860;
  wire [0:0] v_4861;
  wire [0:0] v_4862;
  wire [0:0] v_4863;
  function [0:0] mux_4863(input [0:0] sel);
    case (sel) 0: mux_4863 = 1'h0; 1: mux_4863 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4864;
  function [0:0] mux_4864(input [0:0] sel);
    case (sel) 0: mux_4864 = 1'h0; 1: mux_4864 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4865 = 1'h0;
  wire [0:0] v_4866;
  wire [0:0] v_4867;
  wire [0:0] act_4868;
  wire [0:0] v_4869;
  wire [0:0] v_4870;
  wire [0:0] v_4871;
  reg [0:0] v_4872 = 1'h0;
  wire [0:0] v_4873;
  wire [0:0] v_4874;
  wire [0:0] act_4875;
  wire [0:0] v_4876;
  wire [0:0] v_4877;
  wire [0:0] v_4878;
  wire [0:0] v_4879;
  wire [0:0] v_4880;
  wire [0:0] v_4881;
  function [0:0] mux_4881(input [0:0] sel);
    case (sel) 0: mux_4881 = 1'h0; 1: mux_4881 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4882;
  wire [0:0] v_4883;
  function [0:0] mux_4883(input [0:0] sel);
    case (sel) 0: mux_4883 = 1'h0; 1: mux_4883 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4884;
  wire [0:0] v_4885;
  wire [0:0] v_4886;
  wire [0:0] v_4887;
  function [0:0] mux_4887(input [0:0] sel);
    case (sel) 0: mux_4887 = 1'h0; 1: mux_4887 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4888;
  function [0:0] mux_4888(input [0:0] sel);
    case (sel) 0: mux_4888 = 1'h0; 1: mux_4888 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4889 = 1'h0;
  wire [0:0] v_4890;
  wire [0:0] v_4891;
  wire [0:0] act_4892;
  wire [0:0] v_4893;
  wire [0:0] v_4894;
  wire [0:0] v_4895;
  wire [0:0] v_4896;
  wire [0:0] v_4897;
  wire [0:0] v_4898;
  function [0:0] mux_4898(input [0:0] sel);
    case (sel) 0: mux_4898 = 1'h0; 1: mux_4898 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4899;
  function [0:0] mux_4899(input [0:0] sel);
    case (sel) 0: mux_4899 = 1'h0; 1: mux_4899 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4900;
  wire [0:0] v_4901;
  wire [0:0] v_4902;
  wire [0:0] v_4903;
  function [0:0] mux_4903(input [0:0] sel);
    case (sel) 0: mux_4903 = 1'h0; 1: mux_4903 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4904;
  function [0:0] mux_4904(input [0:0] sel);
    case (sel) 0: mux_4904 = 1'h0; 1: mux_4904 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4905;
  wire [0:0] v_4906;
  wire [0:0] v_4907;
  wire [0:0] v_4908;
  wire [0:0] v_4909;
  wire [0:0] v_4910;
  function [0:0] mux_4910(input [0:0] sel);
    case (sel) 0: mux_4910 = 1'h0; 1: mux_4910 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4911;
  function [0:0] mux_4911(input [0:0] sel);
    case (sel) 0: mux_4911 = 1'h0; 1: mux_4911 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4912;
  wire [0:0] v_4913;
  wire [0:0] v_4914;
  wire [0:0] v_4915;
  function [0:0] mux_4915(input [0:0] sel);
    case (sel) 0: mux_4915 = 1'h0; 1: mux_4915 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4916;
  function [0:0] mux_4916(input [0:0] sel);
    case (sel) 0: mux_4916 = 1'h0; 1: mux_4916 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4917;
  wire [0:0] v_4918;
  wire [0:0] v_4919;
  wire [0:0] v_4920;
  wire [0:0] v_4921;
  wire [0:0] v_4922;
  function [0:0] mux_4922(input [0:0] sel);
    case (sel) 0: mux_4922 = 1'h0; 1: mux_4922 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4923;
  wire [0:0] v_4924;
  function [0:0] mux_4924(input [0:0] sel);
    case (sel) 0: mux_4924 = 1'h0; 1: mux_4924 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4925;
  wire [0:0] v_4926;
  wire [0:0] v_4927;
  wire [0:0] v_4928;
  function [0:0] mux_4928(input [0:0] sel);
    case (sel) 0: mux_4928 = 1'h0; 1: mux_4928 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4929;
  function [0:0] mux_4929(input [0:0] sel);
    case (sel) 0: mux_4929 = 1'h0; 1: mux_4929 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4930 = 1'h0;
  wire [0:0] v_4931;
  wire [0:0] v_4932;
  wire [0:0] act_4933;
  wire [0:0] v_4934;
  wire [0:0] v_4935;
  wire [0:0] v_4936;
  reg [0:0] v_4937 = 1'h0;
  wire [0:0] v_4938;
  wire [0:0] v_4939;
  wire [0:0] act_4940;
  wire [0:0] v_4941;
  wire [0:0] v_4942;
  wire [0:0] v_4943;
  reg [0:0] v_4944 = 1'h0;
  wire [0:0] v_4945;
  wire [0:0] v_4946;
  wire [0:0] act_4947;
  wire [0:0] v_4948;
  wire [0:0] v_4949;
  wire [0:0] v_4950;
  wire [0:0] v_4951;
  wire [0:0] v_4952;
  wire [0:0] v_4953;
  function [0:0] mux_4953(input [0:0] sel);
    case (sel) 0: mux_4953 = 1'h0; 1: mux_4953 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4954;
  wire [0:0] v_4955;
  function [0:0] mux_4955(input [0:0] sel);
    case (sel) 0: mux_4955 = 1'h0; 1: mux_4955 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4956;
  wire [0:0] v_4957;
  wire [0:0] v_4958;
  wire [0:0] v_4959;
  function [0:0] mux_4959(input [0:0] sel);
    case (sel) 0: mux_4959 = 1'h0; 1: mux_4959 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4960;
  function [0:0] mux_4960(input [0:0] sel);
    case (sel) 0: mux_4960 = 1'h0; 1: mux_4960 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4961 = 1'h0;
  wire [0:0] v_4962;
  wire [0:0] v_4963;
  wire [0:0] act_4964;
  wire [0:0] v_4965;
  wire [0:0] v_4966;
  wire [0:0] v_4967;
  wire [0:0] v_4968;
  wire [0:0] v_4969;
  wire [0:0] v_4970;
  function [0:0] mux_4970(input [0:0] sel);
    case (sel) 0: mux_4970 = 1'h0; 1: mux_4970 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4971;
  function [0:0] mux_4971(input [0:0] sel);
    case (sel) 0: mux_4971 = 1'h0; 1: mux_4971 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4972;
  wire [0:0] v_4973;
  wire [0:0] v_4974;
  wire [0:0] v_4975;
  function [0:0] mux_4975(input [0:0] sel);
    case (sel) 0: mux_4975 = 1'h0; 1: mux_4975 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4976;
  function [0:0] mux_4976(input [0:0] sel);
    case (sel) 0: mux_4976 = 1'h0; 1: mux_4976 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4977;
  wire [0:0] v_4978;
  wire [0:0] v_4979;
  wire [0:0] v_4980;
  wire [0:0] v_4981;
  wire [0:0] v_4982;
  function [0:0] mux_4982(input [0:0] sel);
    case (sel) 0: mux_4982 = 1'h0; 1: mux_4982 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4983;
  wire [0:0] v_4984;
  function [0:0] mux_4984(input [0:0] sel);
    case (sel) 0: mux_4984 = 1'h0; 1: mux_4984 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_4985;
  wire [0:0] v_4986;
  wire [0:0] v_4987;
  wire [0:0] v_4988;
  function [0:0] mux_4988(input [0:0] sel);
    case (sel) 0: mux_4988 = 1'h0; 1: mux_4988 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_4989;
  function [0:0] mux_4989(input [0:0] sel);
    case (sel) 0: mux_4989 = 1'h0; 1: mux_4989 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_4990 = 1'h0;
  wire [0:0] v_4991;
  wire [0:0] v_4992;
  wire [0:0] act_4993;
  wire [0:0] v_4994;
  wire [0:0] v_4995;
  wire [0:0] v_4996;
  reg [0:0] v_4997 = 1'h0;
  wire [0:0] v_4998;
  wire [0:0] v_4999;
  wire [0:0] act_5000;
  wire [0:0] v_5001;
  wire [0:0] v_5002;
  wire [0:0] v_5003;
  wire [0:0] v_5004;
  wire [0:0] v_5005;
  wire [0:0] v_5006;
  function [0:0] mux_5006(input [0:0] sel);
    case (sel) 0: mux_5006 = 1'h0; 1: mux_5006 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5007;
  wire [0:0] v_5008;
  function [0:0] mux_5008(input [0:0] sel);
    case (sel) 0: mux_5008 = 1'h0; 1: mux_5008 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5009;
  wire [0:0] v_5010;
  wire [0:0] v_5011;
  wire [0:0] v_5012;
  function [0:0] mux_5012(input [0:0] sel);
    case (sel) 0: mux_5012 = 1'h0; 1: mux_5012 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5013;
  function [0:0] mux_5013(input [0:0] sel);
    case (sel) 0: mux_5013 = 1'h0; 1: mux_5013 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5014 = 1'h0;
  wire [0:0] v_5015;
  wire [0:0] v_5016;
  wire [0:0] act_5017;
  wire [0:0] v_5018;
  wire [0:0] v_5019;
  wire [0:0] v_5020;
  wire [0:0] v_5021;
  wire [0:0] v_5022;
  wire [0:0] v_5023;
  function [0:0] mux_5023(input [0:0] sel);
    case (sel) 0: mux_5023 = 1'h0; 1: mux_5023 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5024;
  function [0:0] mux_5024(input [0:0] sel);
    case (sel) 0: mux_5024 = 1'h0; 1: mux_5024 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5025;
  wire [0:0] v_5026;
  wire [0:0] v_5027;
  wire [0:0] v_5028;
  function [0:0] mux_5028(input [0:0] sel);
    case (sel) 0: mux_5028 = 1'h0; 1: mux_5028 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5029;
  function [0:0] mux_5029(input [0:0] sel);
    case (sel) 0: mux_5029 = 1'h0; 1: mux_5029 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5030;
  wire [0:0] v_5031;
  wire [0:0] v_5032;
  wire [0:0] v_5033;
  wire [0:0] v_5034;
  wire [0:0] v_5035;
  function [0:0] mux_5035(input [0:0] sel);
    case (sel) 0: mux_5035 = 1'h0; 1: mux_5035 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5036;
  function [0:0] mux_5036(input [0:0] sel);
    case (sel) 0: mux_5036 = 1'h0; 1: mux_5036 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5037;
  wire [0:0] v_5038;
  wire [0:0] v_5039;
  wire [0:0] v_5040;
  function [0:0] mux_5040(input [0:0] sel);
    case (sel) 0: mux_5040 = 1'h0; 1: mux_5040 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5041;
  function [0:0] mux_5041(input [0:0] sel);
    case (sel) 0: mux_5041 = 1'h0; 1: mux_5041 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5042;
  wire [0:0] v_5043;
  wire [0:0] v_5044;
  wire [0:0] v_5045;
  wire [0:0] v_5046;
  wire [0:0] v_5047;
  function [0:0] mux_5047(input [0:0] sel);
    case (sel) 0: mux_5047 = 1'h0; 1: mux_5047 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5048;
  function [0:0] mux_5048(input [0:0] sel);
    case (sel) 0: mux_5048 = 1'h0; 1: mux_5048 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5049;
  wire [0:0] v_5050;
  wire [0:0] v_5051;
  wire [0:0] v_5052;
  function [0:0] mux_5052(input [0:0] sel);
    case (sel) 0: mux_5052 = 1'h0; 1: mux_5052 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5053;
  function [0:0] mux_5053(input [0:0] sel);
    case (sel) 0: mux_5053 = 1'h0; 1: mux_5053 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5054;
  wire [0:0] v_5055;
  wire [0:0] v_5056;
  wire [0:0] v_5057;
  wire [0:0] v_5058;
  wire [0:0] v_5059;
  function [0:0] mux_5059(input [0:0] sel);
    case (sel) 0: mux_5059 = 1'h0; 1: mux_5059 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5060;
  wire [0:0] v_5061;
  function [0:0] mux_5061(input [0:0] sel);
    case (sel) 0: mux_5061 = 1'h0; 1: mux_5061 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5062;
  wire [0:0] v_5063;
  wire [0:0] v_5064;
  wire [0:0] v_5065;
  function [0:0] mux_5065(input [0:0] sel);
    case (sel) 0: mux_5065 = 1'h0; 1: mux_5065 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5066;
  function [0:0] mux_5066(input [0:0] sel);
    case (sel) 0: mux_5066 = 1'h0; 1: mux_5066 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5067 = 1'h0;
  wire [0:0] v_5068;
  wire [0:0] v_5069;
  wire [0:0] act_5070;
  wire [0:0] v_5071;
  wire [0:0] v_5072;
  wire [0:0] v_5073;
  reg [0:0] v_5074 = 1'h0;
  wire [0:0] v_5075;
  wire [0:0] v_5076;
  wire [0:0] act_5077;
  wire [0:0] v_5078;
  wire [0:0] v_5079;
  wire [0:0] v_5080;
  reg [0:0] v_5081 = 1'h0;
  wire [0:0] v_5082;
  wire [0:0] v_5083;
  wire [0:0] act_5084;
  wire [0:0] v_5085;
  wire [0:0] v_5086;
  wire [0:0] v_5087;
  reg [0:0] v_5088 = 1'h0;
  wire [0:0] v_5089;
  wire [0:0] v_5090;
  wire [0:0] act_5091;
  wire [0:0] v_5092;
  wire [0:0] v_5093;
  wire [0:0] v_5094;
  wire [0:0] v_5095;
  wire [0:0] v_5096;
  wire [0:0] v_5097;
  function [0:0] mux_5097(input [0:0] sel);
    case (sel) 0: mux_5097 = 1'h0; 1: mux_5097 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5098;
  wire [0:0] v_5099;
  function [0:0] mux_5099(input [0:0] sel);
    case (sel) 0: mux_5099 = 1'h0; 1: mux_5099 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5100;
  wire [0:0] v_5101;
  wire [0:0] v_5102;
  wire [0:0] v_5103;
  function [0:0] mux_5103(input [0:0] sel);
    case (sel) 0: mux_5103 = 1'h0; 1: mux_5103 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5104;
  function [0:0] mux_5104(input [0:0] sel);
    case (sel) 0: mux_5104 = 1'h0; 1: mux_5104 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5105 = 1'h0;
  wire [0:0] v_5106;
  wire [0:0] v_5107;
  wire [0:0] act_5108;
  wire [0:0] v_5109;
  wire [0:0] v_5110;
  wire [0:0] v_5111;
  wire [0:0] v_5112;
  wire [0:0] v_5113;
  wire [0:0] v_5114;
  function [0:0] mux_5114(input [0:0] sel);
    case (sel) 0: mux_5114 = 1'h0; 1: mux_5114 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5115;
  function [0:0] mux_5115(input [0:0] sel);
    case (sel) 0: mux_5115 = 1'h0; 1: mux_5115 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5116;
  wire [0:0] v_5117;
  wire [0:0] v_5118;
  wire [0:0] v_5119;
  function [0:0] mux_5119(input [0:0] sel);
    case (sel) 0: mux_5119 = 1'h0; 1: mux_5119 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5120;
  function [0:0] mux_5120(input [0:0] sel);
    case (sel) 0: mux_5120 = 1'h0; 1: mux_5120 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5121;
  wire [0:0] v_5122;
  wire [0:0] v_5123;
  wire [0:0] v_5124;
  wire [0:0] v_5125;
  wire [0:0] v_5126;
  function [0:0] mux_5126(input [0:0] sel);
    case (sel) 0: mux_5126 = 1'h0; 1: mux_5126 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5127;
  wire [0:0] v_5128;
  function [0:0] mux_5128(input [0:0] sel);
    case (sel) 0: mux_5128 = 1'h0; 1: mux_5128 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5129;
  wire [0:0] v_5130;
  wire [0:0] v_5131;
  wire [0:0] v_5132;
  function [0:0] mux_5132(input [0:0] sel);
    case (sel) 0: mux_5132 = 1'h0; 1: mux_5132 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5133;
  function [0:0] mux_5133(input [0:0] sel);
    case (sel) 0: mux_5133 = 1'h0; 1: mux_5133 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5134 = 1'h0;
  wire [0:0] v_5135;
  wire [0:0] v_5136;
  wire [0:0] act_5137;
  wire [0:0] v_5138;
  wire [0:0] v_5139;
  wire [0:0] v_5140;
  reg [0:0] v_5141 = 1'h0;
  wire [0:0] v_5142;
  wire [0:0] v_5143;
  wire [0:0] act_5144;
  wire [0:0] v_5145;
  wire [0:0] v_5146;
  wire [0:0] v_5147;
  wire [0:0] v_5148;
  wire [0:0] v_5149;
  wire [0:0] v_5150;
  function [0:0] mux_5150(input [0:0] sel);
    case (sel) 0: mux_5150 = 1'h0; 1: mux_5150 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5151;
  wire [0:0] v_5152;
  function [0:0] mux_5152(input [0:0] sel);
    case (sel) 0: mux_5152 = 1'h0; 1: mux_5152 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5153;
  wire [0:0] v_5154;
  wire [0:0] v_5155;
  wire [0:0] v_5156;
  function [0:0] mux_5156(input [0:0] sel);
    case (sel) 0: mux_5156 = 1'h0; 1: mux_5156 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5157;
  function [0:0] mux_5157(input [0:0] sel);
    case (sel) 0: mux_5157 = 1'h0; 1: mux_5157 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5158 = 1'h0;
  wire [0:0] v_5159;
  wire [0:0] v_5160;
  wire [0:0] act_5161;
  wire [0:0] v_5162;
  wire [0:0] v_5163;
  wire [0:0] v_5164;
  wire [0:0] v_5165;
  wire [0:0] v_5166;
  wire [0:0] v_5167;
  function [0:0] mux_5167(input [0:0] sel);
    case (sel) 0: mux_5167 = 1'h0; 1: mux_5167 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5168;
  function [0:0] mux_5168(input [0:0] sel);
    case (sel) 0: mux_5168 = 1'h0; 1: mux_5168 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5169;
  wire [0:0] v_5170;
  wire [0:0] v_5171;
  wire [0:0] v_5172;
  function [0:0] mux_5172(input [0:0] sel);
    case (sel) 0: mux_5172 = 1'h0; 1: mux_5172 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5173;
  function [0:0] mux_5173(input [0:0] sel);
    case (sel) 0: mux_5173 = 1'h0; 1: mux_5173 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5174;
  wire [0:0] v_5175;
  wire [0:0] v_5176;
  wire [0:0] v_5177;
  wire [0:0] v_5178;
  wire [0:0] v_5179;
  function [0:0] mux_5179(input [0:0] sel);
    case (sel) 0: mux_5179 = 1'h0; 1: mux_5179 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5180;
  function [0:0] mux_5180(input [0:0] sel);
    case (sel) 0: mux_5180 = 1'h0; 1: mux_5180 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5181;
  wire [0:0] v_5182;
  wire [0:0] v_5183;
  wire [0:0] v_5184;
  function [0:0] mux_5184(input [0:0] sel);
    case (sel) 0: mux_5184 = 1'h0; 1: mux_5184 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5185;
  function [0:0] mux_5185(input [0:0] sel);
    case (sel) 0: mux_5185 = 1'h0; 1: mux_5185 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5186;
  wire [0:0] v_5187;
  wire [0:0] v_5188;
  wire [0:0] v_5189;
  wire [0:0] v_5190;
  wire [0:0] v_5191;
  function [0:0] mux_5191(input [0:0] sel);
    case (sel) 0: mux_5191 = 1'h0; 1: mux_5191 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5192;
  wire [0:0] v_5193;
  function [0:0] mux_5193(input [0:0] sel);
    case (sel) 0: mux_5193 = 1'h0; 1: mux_5193 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5194;
  wire [0:0] v_5195;
  wire [0:0] v_5196;
  wire [0:0] v_5197;
  function [0:0] mux_5197(input [0:0] sel);
    case (sel) 0: mux_5197 = 1'h0; 1: mux_5197 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5198;
  function [0:0] mux_5198(input [0:0] sel);
    case (sel) 0: mux_5198 = 1'h0; 1: mux_5198 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5199 = 1'h0;
  wire [0:0] v_5200;
  wire [0:0] v_5201;
  wire [0:0] act_5202;
  wire [0:0] v_5203;
  wire [0:0] v_5204;
  wire [0:0] v_5205;
  reg [0:0] v_5206 = 1'h0;
  wire [0:0] v_5207;
  wire [0:0] v_5208;
  wire [0:0] act_5209;
  wire [0:0] v_5210;
  wire [0:0] v_5211;
  wire [0:0] v_5212;
  reg [0:0] v_5213 = 1'h0;
  wire [0:0] v_5214;
  wire [0:0] v_5215;
  wire [0:0] act_5216;
  wire [0:0] v_5217;
  wire [0:0] v_5218;
  wire [0:0] v_5219;
  wire [0:0] v_5220;
  wire [0:0] v_5221;
  wire [0:0] v_5222;
  function [0:0] mux_5222(input [0:0] sel);
    case (sel) 0: mux_5222 = 1'h0; 1: mux_5222 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5223;
  wire [0:0] v_5224;
  function [0:0] mux_5224(input [0:0] sel);
    case (sel) 0: mux_5224 = 1'h0; 1: mux_5224 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5225;
  wire [0:0] v_5226;
  wire [0:0] v_5227;
  wire [0:0] v_5228;
  function [0:0] mux_5228(input [0:0] sel);
    case (sel) 0: mux_5228 = 1'h0; 1: mux_5228 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5229;
  function [0:0] mux_5229(input [0:0] sel);
    case (sel) 0: mux_5229 = 1'h0; 1: mux_5229 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5230 = 1'h0;
  wire [0:0] v_5231;
  wire [0:0] v_5232;
  wire [0:0] act_5233;
  wire [0:0] v_5234;
  wire [0:0] v_5235;
  wire [0:0] v_5236;
  wire [0:0] v_5237;
  wire [0:0] v_5238;
  wire [0:0] v_5239;
  function [0:0] mux_5239(input [0:0] sel);
    case (sel) 0: mux_5239 = 1'h0; 1: mux_5239 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5240;
  function [0:0] mux_5240(input [0:0] sel);
    case (sel) 0: mux_5240 = 1'h0; 1: mux_5240 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5241;
  wire [0:0] v_5242;
  wire [0:0] v_5243;
  wire [0:0] v_5244;
  function [0:0] mux_5244(input [0:0] sel);
    case (sel) 0: mux_5244 = 1'h0; 1: mux_5244 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5245;
  function [0:0] mux_5245(input [0:0] sel);
    case (sel) 0: mux_5245 = 1'h0; 1: mux_5245 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5246;
  wire [0:0] v_5247;
  wire [0:0] v_5248;
  wire [0:0] v_5249;
  wire [0:0] v_5250;
  wire [0:0] v_5251;
  function [0:0] mux_5251(input [0:0] sel);
    case (sel) 0: mux_5251 = 1'h0; 1: mux_5251 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5252;
  wire [0:0] v_5253;
  function [0:0] mux_5253(input [0:0] sel);
    case (sel) 0: mux_5253 = 1'h0; 1: mux_5253 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5254;
  wire [0:0] v_5255;
  wire [0:0] v_5256;
  wire [0:0] v_5257;
  function [0:0] mux_5257(input [0:0] sel);
    case (sel) 0: mux_5257 = 1'h0; 1: mux_5257 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5258;
  function [0:0] mux_5258(input [0:0] sel);
    case (sel) 0: mux_5258 = 1'h0; 1: mux_5258 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5259 = 1'h0;
  wire [0:0] v_5260;
  wire [0:0] v_5261;
  wire [0:0] act_5262;
  wire [0:0] v_5263;
  wire [0:0] v_5264;
  wire [0:0] v_5265;
  reg [0:0] v_5266 = 1'h0;
  wire [0:0] v_5267;
  wire [0:0] v_5268;
  wire [0:0] act_5269;
  wire [0:0] v_5270;
  wire [0:0] v_5271;
  wire [0:0] v_5272;
  wire [0:0] v_5273;
  wire [0:0] v_5274;
  wire [0:0] v_5275;
  function [0:0] mux_5275(input [0:0] sel);
    case (sel) 0: mux_5275 = 1'h0; 1: mux_5275 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5276;
  wire [0:0] v_5277;
  function [0:0] mux_5277(input [0:0] sel);
    case (sel) 0: mux_5277 = 1'h0; 1: mux_5277 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5278;
  wire [0:0] v_5279;
  wire [0:0] v_5280;
  wire [0:0] v_5281;
  function [0:0] mux_5281(input [0:0] sel);
    case (sel) 0: mux_5281 = 1'h0; 1: mux_5281 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5282;
  function [0:0] mux_5282(input [0:0] sel);
    case (sel) 0: mux_5282 = 1'h0; 1: mux_5282 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5283 = 1'h0;
  wire [0:0] v_5284;
  wire [0:0] v_5285;
  wire [0:0] act_5286;
  wire [0:0] v_5287;
  wire [0:0] v_5288;
  wire [0:0] v_5289;
  wire [0:0] v_5290;
  wire [0:0] v_5291;
  wire [0:0] v_5292;
  function [0:0] mux_5292(input [0:0] sel);
    case (sel) 0: mux_5292 = 1'h0; 1: mux_5292 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5293;
  function [0:0] mux_5293(input [0:0] sel);
    case (sel) 0: mux_5293 = 1'h0; 1: mux_5293 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5294;
  wire [0:0] v_5295;
  wire [0:0] v_5296;
  wire [0:0] v_5297;
  function [0:0] mux_5297(input [0:0] sel);
    case (sel) 0: mux_5297 = 1'h0; 1: mux_5297 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5298;
  function [0:0] mux_5298(input [0:0] sel);
    case (sel) 0: mux_5298 = 1'h0; 1: mux_5298 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5299;
  wire [0:0] v_5300;
  wire [0:0] v_5301;
  wire [0:0] v_5302;
  wire [0:0] v_5303;
  wire [0:0] v_5304;
  function [0:0] mux_5304(input [0:0] sel);
    case (sel) 0: mux_5304 = 1'h0; 1: mux_5304 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5305;
  function [0:0] mux_5305(input [0:0] sel);
    case (sel) 0: mux_5305 = 1'h0; 1: mux_5305 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5306;
  wire [0:0] v_5307;
  wire [0:0] v_5308;
  wire [0:0] v_5309;
  function [0:0] mux_5309(input [0:0] sel);
    case (sel) 0: mux_5309 = 1'h0; 1: mux_5309 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5310;
  function [0:0] mux_5310(input [0:0] sel);
    case (sel) 0: mux_5310 = 1'h0; 1: mux_5310 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5311;
  wire [0:0] v_5312;
  wire [0:0] v_5313;
  wire [0:0] v_5314;
  wire [0:0] v_5315;
  wire [0:0] v_5316;
  function [0:0] mux_5316(input [0:0] sel);
    case (sel) 0: mux_5316 = 1'h0; 1: mux_5316 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5317;
  function [0:0] mux_5317(input [0:0] sel);
    case (sel) 0: mux_5317 = 1'h0; 1: mux_5317 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5318;
  wire [0:0] v_5319;
  wire [0:0] v_5320;
  wire [0:0] v_5321;
  function [0:0] mux_5321(input [0:0] sel);
    case (sel) 0: mux_5321 = 1'h0; 1: mux_5321 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5322;
  function [0:0] mux_5322(input [0:0] sel);
    case (sel) 0: mux_5322 = 1'h0; 1: mux_5322 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5323;
  wire [0:0] v_5324;
  wire [0:0] v_5325;
  wire [0:0] v_5326;
  wire [0:0] v_5327;
  wire [0:0] v_5328;
  function [0:0] mux_5328(input [0:0] sel);
    case (sel) 0: mux_5328 = 1'h0; 1: mux_5328 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5329;
  function [0:0] mux_5329(input [0:0] sel);
    case (sel) 0: mux_5329 = 1'h0; 1: mux_5329 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5330;
  wire [0:0] v_5331;
  wire [0:0] v_5332;
  wire [0:0] v_5333;
  function [0:0] mux_5333(input [0:0] sel);
    case (sel) 0: mux_5333 = 1'h0; 1: mux_5333 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5334;
  function [0:0] mux_5334(input [0:0] sel);
    case (sel) 0: mux_5334 = 1'h0; 1: mux_5334 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5335;
  wire [0:0] v_5336;
  wire [0:0] v_5337;
  wire [0:0] v_5338;
  wire [0:0] v_5339;
  wire [0:0] v_5340;
  function [0:0] mux_5340(input [0:0] sel);
    case (sel) 0: mux_5340 = 1'h0; 1: mux_5340 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5341;
  function [0:0] mux_5341(input [0:0] sel);
    case (sel) 0: mux_5341 = 1'h0; 1: mux_5341 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5342;
  wire [0:0] v_5343;
  wire [0:0] v_5344;
  wire [0:0] v_5345;
  function [0:0] mux_5345(input [0:0] sel);
    case (sel) 0: mux_5345 = 1'h0; 1: mux_5345 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5346;
  function [0:0] mux_5346(input [0:0] sel);
    case (sel) 0: mux_5346 = 1'h0; 1: mux_5346 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5347;
  wire [0:0] v_5348;
  wire [0:0] v_5349;
  wire [0:0] v_5350;
  wire [0:0] v_5351;
  wire [0:0] v_5352;
  function [0:0] mux_5352(input [0:0] sel);
    case (sel) 0: mux_5352 = 1'h0; 1: mux_5352 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5353;
  function [0:0] mux_5353(input [0:0] sel);
    case (sel) 0: mux_5353 = 1'h0; 1: mux_5353 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5354;
  wire [0:0] v_5355;
  wire [0:0] v_5356;
  wire [0:0] v_5357;
  function [0:0] mux_5357(input [0:0] sel);
    case (sel) 0: mux_5357 = 1'h0; 1: mux_5357 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5358;
  function [0:0] mux_5358(input [0:0] sel);
    case (sel) 0: mux_5358 = 1'h0; 1: mux_5358 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5359;
  wire [0:0] v_5360;
  wire [0:0] v_5361;
  wire [0:0] v_5362;
  wire [0:0] v_5363;
  wire [0:0] v_5364;
  function [0:0] mux_5364(input [0:0] sel);
    case (sel) 0: mux_5364 = 1'h0; 1: mux_5364 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5365;
  function [0:0] mux_5365(input [0:0] sel);
    case (sel) 0: mux_5365 = 1'h0; 1: mux_5365 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5366;
  wire [0:0] v_5367;
  wire [0:0] v_5368;
  wire [0:0] v_5369;
  function [0:0] mux_5369(input [0:0] sel);
    case (sel) 0: mux_5369 = 1'h0; 1: mux_5369 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5370;
  function [0:0] mux_5370(input [0:0] sel);
    case (sel) 0: mux_5370 = 1'h0; 1: mux_5370 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5371;
  wire [0:0] v_5372;
  wire [0:0] v_5373;
  wire [0:0] v_5374;
  wire [0:0] v_5375;
  wire [0:0] v_5376;
  function [0:0] mux_5376(input [0:0] sel);
    case (sel) 0: mux_5376 = 1'h0; 1: mux_5376 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5377;
  wire [0:0] v_5378;
  function [0:0] mux_5378(input [0:0] sel);
    case (sel) 0: mux_5378 = 1'h0; 1: mux_5378 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5379;
  wire [0:0] v_5380;
  wire [0:0] v_5381;
  wire [0:0] v_5382;
  function [0:0] mux_5382(input [0:0] sel);
    case (sel) 0: mux_5382 = 1'h0; 1: mux_5382 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5383;
  function [0:0] mux_5383(input [0:0] sel);
    case (sel) 0: mux_5383 = 1'h0; 1: mux_5383 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5384 = 1'h0;
  wire [0:0] v_5385;
  wire [0:0] v_5386;
  wire [0:0] act_5387;
  wire [0:0] v_5388;
  wire [0:0] v_5389;
  wire [0:0] v_5390;
  reg [0:0] v_5391 = 1'h0;
  wire [0:0] v_5392;
  wire [0:0] v_5393;
  wire [0:0] act_5394;
  wire [0:0] v_5395;
  wire [0:0] v_5396;
  wire [0:0] v_5397;
  reg [0:0] v_5398 = 1'h0;
  wire [0:0] v_5399;
  wire [0:0] v_5400;
  wire [0:0] act_5401;
  wire [0:0] v_5402;
  wire [0:0] v_5403;
  wire [0:0] v_5404;
  reg [0:0] v_5405 = 1'h0;
  wire [0:0] v_5406;
  wire [0:0] v_5407;
  wire [0:0] act_5408;
  wire [0:0] v_5409;
  wire [0:0] v_5410;
  wire [0:0] v_5411;
  reg [0:0] v_5412 = 1'h0;
  wire [0:0] v_5413;
  wire [0:0] v_5414;
  wire [0:0] act_5415;
  wire [0:0] v_5416;
  wire [0:0] v_5417;
  wire [0:0] v_5418;
  reg [0:0] v_5419 = 1'h0;
  wire [0:0] v_5420;
  wire [0:0] v_5421;
  wire [0:0] act_5422;
  wire [0:0] v_5423;
  wire [0:0] v_5424;
  wire [0:0] v_5425;
  reg [0:0] v_5426 = 1'h0;
  wire [0:0] v_5427;
  wire [0:0] v_5428;
  wire [0:0] act_5429;
  wire [0:0] v_5430;
  wire [0:0] v_5431;
  wire [0:0] v_5432;
  reg [0:0] v_5433 = 1'h0;
  wire [0:0] v_5434;
  wire [0:0] v_5435;
  wire [0:0] act_5436;
  wire [0:0] v_5437;
  wire [0:0] v_5438;
  wire [0:0] v_5439;
  wire [0:0] v_5440;
  wire [0:0] v_5441;
  wire [0:0] v_5442;
  function [0:0] mux_5442(input [0:0] sel);
    case (sel) 0: mux_5442 = 1'h0; 1: mux_5442 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5443;
  wire [0:0] v_5444;
  function [0:0] mux_5444(input [0:0] sel);
    case (sel) 0: mux_5444 = 1'h0; 1: mux_5444 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5445;
  wire [0:0] v_5446;
  wire [0:0] v_5447;
  wire [0:0] v_5448;
  function [0:0] mux_5448(input [0:0] sel);
    case (sel) 0: mux_5448 = 1'h0; 1: mux_5448 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5449;
  function [0:0] mux_5449(input [0:0] sel);
    case (sel) 0: mux_5449 = 1'h0; 1: mux_5449 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5450 = 1'h0;
  wire [0:0] v_5451;
  wire [0:0] v_5452;
  wire [0:0] act_5453;
  wire [0:0] v_5454;
  wire [0:0] v_5455;
  wire [0:0] v_5456;
  wire [0:0] v_5457;
  wire [0:0] v_5458;
  wire [0:0] v_5459;
  function [0:0] mux_5459(input [0:0] sel);
    case (sel) 0: mux_5459 = 1'h0; 1: mux_5459 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5460;
  function [0:0] mux_5460(input [0:0] sel);
    case (sel) 0: mux_5460 = 1'h0; 1: mux_5460 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5461;
  wire [0:0] v_5462;
  wire [0:0] v_5463;
  wire [0:0] v_5464;
  function [0:0] mux_5464(input [0:0] sel);
    case (sel) 0: mux_5464 = 1'h0; 1: mux_5464 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5465;
  function [0:0] mux_5465(input [0:0] sel);
    case (sel) 0: mux_5465 = 1'h0; 1: mux_5465 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5466;
  wire [0:0] v_5467;
  wire [0:0] v_5468;
  wire [0:0] v_5469;
  wire [0:0] v_5470;
  wire [0:0] v_5471;
  function [0:0] mux_5471(input [0:0] sel);
    case (sel) 0: mux_5471 = 1'h0; 1: mux_5471 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5472;
  wire [0:0] v_5473;
  function [0:0] mux_5473(input [0:0] sel);
    case (sel) 0: mux_5473 = 1'h0; 1: mux_5473 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5474;
  wire [0:0] v_5475;
  wire [0:0] v_5476;
  wire [0:0] v_5477;
  function [0:0] mux_5477(input [0:0] sel);
    case (sel) 0: mux_5477 = 1'h0; 1: mux_5477 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5478;
  function [0:0] mux_5478(input [0:0] sel);
    case (sel) 0: mux_5478 = 1'h0; 1: mux_5478 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5479 = 1'h0;
  wire [0:0] v_5480;
  wire [0:0] v_5481;
  wire [0:0] act_5482;
  wire [0:0] v_5483;
  wire [0:0] v_5484;
  wire [0:0] v_5485;
  reg [0:0] v_5486 = 1'h0;
  wire [0:0] v_5487;
  wire [0:0] v_5488;
  wire [0:0] act_5489;
  wire [0:0] v_5490;
  wire [0:0] v_5491;
  wire [0:0] v_5492;
  wire [0:0] v_5493;
  wire [0:0] v_5494;
  wire [0:0] v_5495;
  function [0:0] mux_5495(input [0:0] sel);
    case (sel) 0: mux_5495 = 1'h0; 1: mux_5495 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5496;
  wire [0:0] v_5497;
  function [0:0] mux_5497(input [0:0] sel);
    case (sel) 0: mux_5497 = 1'h0; 1: mux_5497 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5498;
  wire [0:0] v_5499;
  wire [0:0] v_5500;
  wire [0:0] v_5501;
  function [0:0] mux_5501(input [0:0] sel);
    case (sel) 0: mux_5501 = 1'h0; 1: mux_5501 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5502;
  function [0:0] mux_5502(input [0:0] sel);
    case (sel) 0: mux_5502 = 1'h0; 1: mux_5502 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5503 = 1'h0;
  wire [0:0] v_5504;
  wire [0:0] v_5505;
  wire [0:0] act_5506;
  wire [0:0] v_5507;
  wire [0:0] v_5508;
  wire [0:0] v_5509;
  wire [0:0] v_5510;
  wire [0:0] v_5511;
  wire [0:0] v_5512;
  function [0:0] mux_5512(input [0:0] sel);
    case (sel) 0: mux_5512 = 1'h0; 1: mux_5512 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5513;
  function [0:0] mux_5513(input [0:0] sel);
    case (sel) 0: mux_5513 = 1'h0; 1: mux_5513 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5514;
  wire [0:0] v_5515;
  wire [0:0] v_5516;
  wire [0:0] v_5517;
  function [0:0] mux_5517(input [0:0] sel);
    case (sel) 0: mux_5517 = 1'h0; 1: mux_5517 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5518;
  function [0:0] mux_5518(input [0:0] sel);
    case (sel) 0: mux_5518 = 1'h0; 1: mux_5518 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5519;
  wire [0:0] v_5520;
  wire [0:0] v_5521;
  wire [0:0] v_5522;
  wire [0:0] v_5523;
  wire [0:0] v_5524;
  function [0:0] mux_5524(input [0:0] sel);
    case (sel) 0: mux_5524 = 1'h0; 1: mux_5524 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5525;
  function [0:0] mux_5525(input [0:0] sel);
    case (sel) 0: mux_5525 = 1'h0; 1: mux_5525 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5526;
  wire [0:0] v_5527;
  wire [0:0] v_5528;
  wire [0:0] v_5529;
  function [0:0] mux_5529(input [0:0] sel);
    case (sel) 0: mux_5529 = 1'h0; 1: mux_5529 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5530;
  function [0:0] mux_5530(input [0:0] sel);
    case (sel) 0: mux_5530 = 1'h0; 1: mux_5530 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5531;
  wire [0:0] v_5532;
  wire [0:0] v_5533;
  wire [0:0] v_5534;
  wire [0:0] v_5535;
  wire [0:0] v_5536;
  function [0:0] mux_5536(input [0:0] sel);
    case (sel) 0: mux_5536 = 1'h0; 1: mux_5536 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5537;
  wire [0:0] v_5538;
  function [0:0] mux_5538(input [0:0] sel);
    case (sel) 0: mux_5538 = 1'h0; 1: mux_5538 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5539;
  wire [0:0] v_5540;
  wire [0:0] v_5541;
  wire [0:0] v_5542;
  function [0:0] mux_5542(input [0:0] sel);
    case (sel) 0: mux_5542 = 1'h0; 1: mux_5542 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5543;
  function [0:0] mux_5543(input [0:0] sel);
    case (sel) 0: mux_5543 = 1'h0; 1: mux_5543 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5544 = 1'h0;
  wire [0:0] v_5545;
  wire [0:0] v_5546;
  wire [0:0] act_5547;
  wire [0:0] v_5548;
  wire [0:0] v_5549;
  wire [0:0] v_5550;
  reg [0:0] v_5551 = 1'h0;
  wire [0:0] v_5552;
  wire [0:0] v_5553;
  wire [0:0] act_5554;
  wire [0:0] v_5555;
  wire [0:0] v_5556;
  wire [0:0] v_5557;
  reg [0:0] v_5558 = 1'h0;
  wire [0:0] v_5559;
  wire [0:0] v_5560;
  wire [0:0] act_5561;
  wire [0:0] v_5562;
  wire [0:0] v_5563;
  wire [0:0] v_5564;
  wire [0:0] v_5565;
  wire [0:0] v_5566;
  wire [0:0] v_5567;
  function [0:0] mux_5567(input [0:0] sel);
    case (sel) 0: mux_5567 = 1'h0; 1: mux_5567 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5568;
  wire [0:0] v_5569;
  function [0:0] mux_5569(input [0:0] sel);
    case (sel) 0: mux_5569 = 1'h0; 1: mux_5569 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5570;
  wire [0:0] v_5571;
  wire [0:0] v_5572;
  wire [0:0] v_5573;
  function [0:0] mux_5573(input [0:0] sel);
    case (sel) 0: mux_5573 = 1'h0; 1: mux_5573 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5574;
  function [0:0] mux_5574(input [0:0] sel);
    case (sel) 0: mux_5574 = 1'h0; 1: mux_5574 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5575 = 1'h0;
  wire [0:0] v_5576;
  wire [0:0] v_5577;
  wire [0:0] act_5578;
  wire [0:0] v_5579;
  wire [0:0] v_5580;
  wire [0:0] v_5581;
  wire [0:0] v_5582;
  wire [0:0] v_5583;
  wire [0:0] v_5584;
  function [0:0] mux_5584(input [0:0] sel);
    case (sel) 0: mux_5584 = 1'h0; 1: mux_5584 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5585;
  function [0:0] mux_5585(input [0:0] sel);
    case (sel) 0: mux_5585 = 1'h0; 1: mux_5585 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5586;
  wire [0:0] v_5587;
  wire [0:0] v_5588;
  wire [0:0] v_5589;
  function [0:0] mux_5589(input [0:0] sel);
    case (sel) 0: mux_5589 = 1'h0; 1: mux_5589 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5590;
  function [0:0] mux_5590(input [0:0] sel);
    case (sel) 0: mux_5590 = 1'h0; 1: mux_5590 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5591;
  wire [0:0] v_5592;
  wire [0:0] v_5593;
  wire [0:0] v_5594;
  wire [0:0] v_5595;
  wire [0:0] v_5596;
  function [0:0] mux_5596(input [0:0] sel);
    case (sel) 0: mux_5596 = 1'h0; 1: mux_5596 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5597;
  wire [0:0] v_5598;
  function [0:0] mux_5598(input [0:0] sel);
    case (sel) 0: mux_5598 = 1'h0; 1: mux_5598 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5599;
  wire [0:0] v_5600;
  wire [0:0] v_5601;
  wire [0:0] v_5602;
  function [0:0] mux_5602(input [0:0] sel);
    case (sel) 0: mux_5602 = 1'h0; 1: mux_5602 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5603;
  function [0:0] mux_5603(input [0:0] sel);
    case (sel) 0: mux_5603 = 1'h0; 1: mux_5603 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5604 = 1'h0;
  wire [0:0] v_5605;
  wire [0:0] v_5606;
  wire [0:0] act_5607;
  wire [0:0] v_5608;
  wire [0:0] v_5609;
  wire [0:0] v_5610;
  reg [0:0] v_5611 = 1'h0;
  wire [0:0] v_5612;
  wire [0:0] v_5613;
  wire [0:0] act_5614;
  wire [0:0] v_5615;
  wire [0:0] v_5616;
  wire [0:0] v_5617;
  wire [0:0] v_5618;
  wire [0:0] v_5619;
  wire [0:0] v_5620;
  function [0:0] mux_5620(input [0:0] sel);
    case (sel) 0: mux_5620 = 1'h0; 1: mux_5620 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5621;
  wire [0:0] v_5622;
  function [0:0] mux_5622(input [0:0] sel);
    case (sel) 0: mux_5622 = 1'h0; 1: mux_5622 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5623;
  wire [0:0] v_5624;
  wire [0:0] v_5625;
  wire [0:0] v_5626;
  function [0:0] mux_5626(input [0:0] sel);
    case (sel) 0: mux_5626 = 1'h0; 1: mux_5626 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5627;
  function [0:0] mux_5627(input [0:0] sel);
    case (sel) 0: mux_5627 = 1'h0; 1: mux_5627 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5628 = 1'h0;
  wire [0:0] v_5629;
  wire [0:0] v_5630;
  wire [0:0] act_5631;
  wire [0:0] v_5632;
  wire [0:0] v_5633;
  wire [0:0] v_5634;
  wire [0:0] v_5635;
  wire [0:0] v_5636;
  wire [0:0] v_5637;
  function [0:0] mux_5637(input [0:0] sel);
    case (sel) 0: mux_5637 = 1'h0; 1: mux_5637 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5638;
  function [0:0] mux_5638(input [0:0] sel);
    case (sel) 0: mux_5638 = 1'h0; 1: mux_5638 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5639;
  wire [0:0] v_5640;
  wire [0:0] v_5641;
  wire [0:0] v_5642;
  function [0:0] mux_5642(input [0:0] sel);
    case (sel) 0: mux_5642 = 1'h0; 1: mux_5642 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5643;
  function [0:0] mux_5643(input [0:0] sel);
    case (sel) 0: mux_5643 = 1'h0; 1: mux_5643 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5644;
  wire [0:0] v_5645;
  wire [0:0] v_5646;
  wire [0:0] v_5647;
  wire [0:0] v_5648;
  wire [0:0] v_5649;
  function [0:0] mux_5649(input [0:0] sel);
    case (sel) 0: mux_5649 = 1'h0; 1: mux_5649 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5650;
  function [0:0] mux_5650(input [0:0] sel);
    case (sel) 0: mux_5650 = 1'h0; 1: mux_5650 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5651;
  wire [0:0] v_5652;
  wire [0:0] v_5653;
  wire [0:0] v_5654;
  function [0:0] mux_5654(input [0:0] sel);
    case (sel) 0: mux_5654 = 1'h0; 1: mux_5654 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5655;
  function [0:0] mux_5655(input [0:0] sel);
    case (sel) 0: mux_5655 = 1'h0; 1: mux_5655 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5656;
  wire [0:0] v_5657;
  wire [0:0] v_5658;
  wire [0:0] v_5659;
  wire [0:0] v_5660;
  wire [0:0] v_5661;
  function [0:0] mux_5661(input [0:0] sel);
    case (sel) 0: mux_5661 = 1'h0; 1: mux_5661 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5662;
  function [0:0] mux_5662(input [0:0] sel);
    case (sel) 0: mux_5662 = 1'h0; 1: mux_5662 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5663;
  wire [0:0] v_5664;
  wire [0:0] v_5665;
  wire [0:0] v_5666;
  function [0:0] mux_5666(input [0:0] sel);
    case (sel) 0: mux_5666 = 1'h0; 1: mux_5666 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5667;
  function [0:0] mux_5667(input [0:0] sel);
    case (sel) 0: mux_5667 = 1'h0; 1: mux_5667 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5668;
  wire [0:0] v_5669;
  wire [0:0] v_5670;
  wire [0:0] v_5671;
  wire [0:0] v_5672;
  wire [0:0] v_5673;
  function [0:0] mux_5673(input [0:0] sel);
    case (sel) 0: mux_5673 = 1'h0; 1: mux_5673 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5674;
  wire [0:0] v_5675;
  function [0:0] mux_5675(input [0:0] sel);
    case (sel) 0: mux_5675 = 1'h0; 1: mux_5675 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5676;
  wire [0:0] v_5677;
  wire [0:0] v_5678;
  wire [0:0] v_5679;
  function [0:0] mux_5679(input [0:0] sel);
    case (sel) 0: mux_5679 = 1'h0; 1: mux_5679 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5680;
  function [0:0] mux_5680(input [0:0] sel);
    case (sel) 0: mux_5680 = 1'h0; 1: mux_5680 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5681 = 1'h0;
  wire [0:0] v_5682;
  wire [0:0] v_5683;
  wire [0:0] act_5684;
  wire [0:0] v_5685;
  wire [0:0] v_5686;
  wire [0:0] v_5687;
  reg [0:0] v_5688 = 1'h0;
  wire [0:0] v_5689;
  wire [0:0] v_5690;
  wire [0:0] act_5691;
  wire [0:0] v_5692;
  wire [0:0] v_5693;
  wire [0:0] v_5694;
  reg [0:0] v_5695 = 1'h0;
  wire [0:0] v_5696;
  wire [0:0] v_5697;
  wire [0:0] act_5698;
  wire [0:0] v_5699;
  wire [0:0] v_5700;
  wire [0:0] v_5701;
  reg [0:0] v_5702 = 1'h0;
  wire [0:0] v_5703;
  wire [0:0] v_5704;
  wire [0:0] act_5705;
  wire [0:0] v_5706;
  wire [0:0] v_5707;
  wire [0:0] v_5708;
  wire [0:0] v_5709;
  wire [0:0] v_5710;
  wire [0:0] v_5711;
  function [0:0] mux_5711(input [0:0] sel);
    case (sel) 0: mux_5711 = 1'h0; 1: mux_5711 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5712;
  wire [0:0] v_5713;
  function [0:0] mux_5713(input [0:0] sel);
    case (sel) 0: mux_5713 = 1'h0; 1: mux_5713 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5714;
  wire [0:0] v_5715;
  wire [0:0] v_5716;
  wire [0:0] v_5717;
  function [0:0] mux_5717(input [0:0] sel);
    case (sel) 0: mux_5717 = 1'h0; 1: mux_5717 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5718;
  function [0:0] mux_5718(input [0:0] sel);
    case (sel) 0: mux_5718 = 1'h0; 1: mux_5718 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5719 = 1'h0;
  wire [0:0] v_5720;
  wire [0:0] v_5721;
  wire [0:0] act_5722;
  wire [0:0] v_5723;
  wire [0:0] v_5724;
  wire [0:0] v_5725;
  wire [0:0] v_5726;
  wire [0:0] v_5727;
  wire [0:0] v_5728;
  function [0:0] mux_5728(input [0:0] sel);
    case (sel) 0: mux_5728 = 1'h0; 1: mux_5728 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5729;
  function [0:0] mux_5729(input [0:0] sel);
    case (sel) 0: mux_5729 = 1'h0; 1: mux_5729 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5730;
  wire [0:0] v_5731;
  wire [0:0] v_5732;
  wire [0:0] v_5733;
  function [0:0] mux_5733(input [0:0] sel);
    case (sel) 0: mux_5733 = 1'h0; 1: mux_5733 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5734;
  function [0:0] mux_5734(input [0:0] sel);
    case (sel) 0: mux_5734 = 1'h0; 1: mux_5734 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5735;
  wire [0:0] v_5736;
  wire [0:0] v_5737;
  wire [0:0] v_5738;
  wire [0:0] v_5739;
  wire [0:0] v_5740;
  function [0:0] mux_5740(input [0:0] sel);
    case (sel) 0: mux_5740 = 1'h0; 1: mux_5740 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5741;
  wire [0:0] v_5742;
  function [0:0] mux_5742(input [0:0] sel);
    case (sel) 0: mux_5742 = 1'h0; 1: mux_5742 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5743;
  wire [0:0] v_5744;
  wire [0:0] v_5745;
  wire [0:0] v_5746;
  function [0:0] mux_5746(input [0:0] sel);
    case (sel) 0: mux_5746 = 1'h0; 1: mux_5746 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5747;
  function [0:0] mux_5747(input [0:0] sel);
    case (sel) 0: mux_5747 = 1'h0; 1: mux_5747 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5748 = 1'h0;
  wire [0:0] v_5749;
  wire [0:0] v_5750;
  wire [0:0] act_5751;
  wire [0:0] v_5752;
  wire [0:0] v_5753;
  wire [0:0] v_5754;
  reg [0:0] v_5755 = 1'h0;
  wire [0:0] v_5756;
  wire [0:0] v_5757;
  wire [0:0] act_5758;
  wire [0:0] v_5759;
  wire [0:0] v_5760;
  wire [0:0] v_5761;
  wire [0:0] v_5762;
  wire [0:0] v_5763;
  wire [0:0] v_5764;
  function [0:0] mux_5764(input [0:0] sel);
    case (sel) 0: mux_5764 = 1'h0; 1: mux_5764 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5765;
  wire [0:0] v_5766;
  function [0:0] mux_5766(input [0:0] sel);
    case (sel) 0: mux_5766 = 1'h0; 1: mux_5766 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5767;
  wire [0:0] v_5768;
  wire [0:0] v_5769;
  wire [0:0] v_5770;
  function [0:0] mux_5770(input [0:0] sel);
    case (sel) 0: mux_5770 = 1'h0; 1: mux_5770 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5771;
  function [0:0] mux_5771(input [0:0] sel);
    case (sel) 0: mux_5771 = 1'h0; 1: mux_5771 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5772 = 1'h0;
  wire [0:0] v_5773;
  wire [0:0] v_5774;
  wire [0:0] act_5775;
  wire [0:0] v_5776;
  wire [0:0] v_5777;
  wire [0:0] v_5778;
  wire [0:0] v_5779;
  wire [0:0] v_5780;
  wire [0:0] v_5781;
  function [0:0] mux_5781(input [0:0] sel);
    case (sel) 0: mux_5781 = 1'h0; 1: mux_5781 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5782;
  function [0:0] mux_5782(input [0:0] sel);
    case (sel) 0: mux_5782 = 1'h0; 1: mux_5782 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5783;
  wire [0:0] v_5784;
  wire [0:0] v_5785;
  wire [0:0] v_5786;
  function [0:0] mux_5786(input [0:0] sel);
    case (sel) 0: mux_5786 = 1'h0; 1: mux_5786 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5787;
  function [0:0] mux_5787(input [0:0] sel);
    case (sel) 0: mux_5787 = 1'h0; 1: mux_5787 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5788;
  wire [0:0] v_5789;
  wire [0:0] v_5790;
  wire [0:0] v_5791;
  wire [0:0] v_5792;
  wire [0:0] v_5793;
  function [0:0] mux_5793(input [0:0] sel);
    case (sel) 0: mux_5793 = 1'h0; 1: mux_5793 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5794;
  function [0:0] mux_5794(input [0:0] sel);
    case (sel) 0: mux_5794 = 1'h0; 1: mux_5794 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5795;
  wire [0:0] v_5796;
  wire [0:0] v_5797;
  wire [0:0] v_5798;
  function [0:0] mux_5798(input [0:0] sel);
    case (sel) 0: mux_5798 = 1'h0; 1: mux_5798 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5799;
  function [0:0] mux_5799(input [0:0] sel);
    case (sel) 0: mux_5799 = 1'h0; 1: mux_5799 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5800;
  wire [0:0] v_5801;
  wire [0:0] v_5802;
  wire [0:0] v_5803;
  wire [0:0] v_5804;
  wire [0:0] v_5805;
  function [0:0] mux_5805(input [0:0] sel);
    case (sel) 0: mux_5805 = 1'h0; 1: mux_5805 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5806;
  wire [0:0] v_5807;
  function [0:0] mux_5807(input [0:0] sel);
    case (sel) 0: mux_5807 = 1'h0; 1: mux_5807 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5808;
  wire [0:0] v_5809;
  wire [0:0] v_5810;
  wire [0:0] v_5811;
  function [0:0] mux_5811(input [0:0] sel);
    case (sel) 0: mux_5811 = 1'h0; 1: mux_5811 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5812;
  function [0:0] mux_5812(input [0:0] sel);
    case (sel) 0: mux_5812 = 1'h0; 1: mux_5812 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5813 = 1'h0;
  wire [0:0] v_5814;
  wire [0:0] v_5815;
  wire [0:0] act_5816;
  wire [0:0] v_5817;
  wire [0:0] v_5818;
  wire [0:0] v_5819;
  reg [0:0] v_5820 = 1'h0;
  wire [0:0] v_5821;
  wire [0:0] v_5822;
  wire [0:0] act_5823;
  wire [0:0] v_5824;
  wire [0:0] v_5825;
  wire [0:0] v_5826;
  reg [0:0] v_5827 = 1'h0;
  wire [0:0] v_5828;
  wire [0:0] v_5829;
  wire [0:0] act_5830;
  wire [0:0] v_5831;
  wire [0:0] v_5832;
  wire [0:0] v_5833;
  wire [0:0] v_5834;
  wire [0:0] v_5835;
  wire [0:0] v_5836;
  function [0:0] mux_5836(input [0:0] sel);
    case (sel) 0: mux_5836 = 1'h0; 1: mux_5836 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5837;
  wire [0:0] v_5838;
  function [0:0] mux_5838(input [0:0] sel);
    case (sel) 0: mux_5838 = 1'h0; 1: mux_5838 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5839;
  wire [0:0] v_5840;
  wire [0:0] v_5841;
  wire [0:0] v_5842;
  function [0:0] mux_5842(input [0:0] sel);
    case (sel) 0: mux_5842 = 1'h0; 1: mux_5842 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5843;
  function [0:0] mux_5843(input [0:0] sel);
    case (sel) 0: mux_5843 = 1'h0; 1: mux_5843 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5844 = 1'h0;
  wire [0:0] v_5845;
  wire [0:0] v_5846;
  wire [0:0] act_5847;
  wire [0:0] v_5848;
  wire [0:0] v_5849;
  wire [0:0] v_5850;
  wire [0:0] v_5851;
  wire [0:0] v_5852;
  wire [0:0] v_5853;
  function [0:0] mux_5853(input [0:0] sel);
    case (sel) 0: mux_5853 = 1'h0; 1: mux_5853 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5854;
  function [0:0] mux_5854(input [0:0] sel);
    case (sel) 0: mux_5854 = 1'h0; 1: mux_5854 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5855;
  wire [0:0] v_5856;
  wire [0:0] v_5857;
  wire [0:0] v_5858;
  function [0:0] mux_5858(input [0:0] sel);
    case (sel) 0: mux_5858 = 1'h0; 1: mux_5858 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5859;
  function [0:0] mux_5859(input [0:0] sel);
    case (sel) 0: mux_5859 = 1'h0; 1: mux_5859 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5860;
  wire [0:0] v_5861;
  wire [0:0] v_5862;
  wire [0:0] v_5863;
  wire [0:0] v_5864;
  wire [0:0] v_5865;
  function [0:0] mux_5865(input [0:0] sel);
    case (sel) 0: mux_5865 = 1'h0; 1: mux_5865 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5866;
  wire [0:0] v_5867;
  function [0:0] mux_5867(input [0:0] sel);
    case (sel) 0: mux_5867 = 1'h0; 1: mux_5867 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5868;
  wire [0:0] v_5869;
  wire [0:0] v_5870;
  wire [0:0] v_5871;
  function [0:0] mux_5871(input [0:0] sel);
    case (sel) 0: mux_5871 = 1'h0; 1: mux_5871 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5872;
  function [0:0] mux_5872(input [0:0] sel);
    case (sel) 0: mux_5872 = 1'h0; 1: mux_5872 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5873 = 1'h0;
  wire [0:0] v_5874;
  wire [0:0] v_5875;
  wire [0:0] act_5876;
  wire [0:0] v_5877;
  wire [0:0] v_5878;
  wire [0:0] v_5879;
  reg [0:0] v_5880 = 1'h0;
  wire [0:0] v_5881;
  wire [0:0] v_5882;
  wire [0:0] act_5883;
  wire [0:0] v_5884;
  wire [0:0] v_5885;
  wire [0:0] v_5886;
  wire [0:0] v_5887;
  wire [0:0] v_5888;
  wire [0:0] v_5889;
  function [0:0] mux_5889(input [0:0] sel);
    case (sel) 0: mux_5889 = 1'h0; 1: mux_5889 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5890;
  wire [0:0] v_5891;
  function [0:0] mux_5891(input [0:0] sel);
    case (sel) 0: mux_5891 = 1'h0; 1: mux_5891 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5892;
  wire [0:0] v_5893;
  wire [0:0] v_5894;
  wire [0:0] v_5895;
  function [0:0] mux_5895(input [0:0] sel);
    case (sel) 0: mux_5895 = 1'h0; 1: mux_5895 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5896;
  function [0:0] mux_5896(input [0:0] sel);
    case (sel) 0: mux_5896 = 1'h0; 1: mux_5896 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5897 = 1'h0;
  wire [0:0] v_5898;
  wire [0:0] v_5899;
  wire [0:0] act_5900;
  wire [0:0] v_5901;
  wire [0:0] v_5902;
  wire [0:0] v_5903;
  wire [0:0] v_5904;
  wire [0:0] v_5905;
  wire [0:0] v_5906;
  function [0:0] mux_5906(input [0:0] sel);
    case (sel) 0: mux_5906 = 1'h0; 1: mux_5906 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5907;
  function [0:0] mux_5907(input [0:0] sel);
    case (sel) 0: mux_5907 = 1'h0; 1: mux_5907 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5908;
  wire [0:0] v_5909;
  wire [0:0] v_5910;
  wire [0:0] v_5911;
  function [0:0] mux_5911(input [0:0] sel);
    case (sel) 0: mux_5911 = 1'h0; 1: mux_5911 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5912;
  function [0:0] mux_5912(input [0:0] sel);
    case (sel) 0: mux_5912 = 1'h0; 1: mux_5912 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5913;
  wire [0:0] v_5914;
  wire [0:0] v_5915;
  wire [0:0] v_5916;
  wire [0:0] v_5917;
  wire [0:0] v_5918;
  function [0:0] mux_5918(input [0:0] sel);
    case (sel) 0: mux_5918 = 1'h0; 1: mux_5918 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5919;
  function [0:0] mux_5919(input [0:0] sel);
    case (sel) 0: mux_5919 = 1'h0; 1: mux_5919 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5920;
  wire [0:0] v_5921;
  wire [0:0] v_5922;
  wire [0:0] v_5923;
  function [0:0] mux_5923(input [0:0] sel);
    case (sel) 0: mux_5923 = 1'h0; 1: mux_5923 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5924;
  function [0:0] mux_5924(input [0:0] sel);
    case (sel) 0: mux_5924 = 1'h0; 1: mux_5924 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5925;
  wire [0:0] v_5926;
  wire [0:0] v_5927;
  wire [0:0] v_5928;
  wire [0:0] v_5929;
  wire [0:0] v_5930;
  function [0:0] mux_5930(input [0:0] sel);
    case (sel) 0: mux_5930 = 1'h0; 1: mux_5930 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5931;
  function [0:0] mux_5931(input [0:0] sel);
    case (sel) 0: mux_5931 = 1'h0; 1: mux_5931 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5932;
  wire [0:0] v_5933;
  wire [0:0] v_5934;
  wire [0:0] v_5935;
  function [0:0] mux_5935(input [0:0] sel);
    case (sel) 0: mux_5935 = 1'h0; 1: mux_5935 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5936;
  function [0:0] mux_5936(input [0:0] sel);
    case (sel) 0: mux_5936 = 1'h0; 1: mux_5936 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5937;
  wire [0:0] v_5938;
  wire [0:0] v_5939;
  wire [0:0] v_5940;
  wire [0:0] v_5941;
  wire [0:0] v_5942;
  function [0:0] mux_5942(input [0:0] sel);
    case (sel) 0: mux_5942 = 1'h0; 1: mux_5942 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5943;
  function [0:0] mux_5943(input [0:0] sel);
    case (sel) 0: mux_5943 = 1'h0; 1: mux_5943 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5944;
  wire [0:0] v_5945;
  wire [0:0] v_5946;
  wire [0:0] v_5947;
  function [0:0] mux_5947(input [0:0] sel);
    case (sel) 0: mux_5947 = 1'h0; 1: mux_5947 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5948;
  function [0:0] mux_5948(input [0:0] sel);
    case (sel) 0: mux_5948 = 1'h0; 1: mux_5948 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5949;
  wire [0:0] v_5950;
  wire [0:0] v_5951;
  wire [0:0] v_5952;
  wire [0:0] v_5953;
  wire [0:0] v_5954;
  function [0:0] mux_5954(input [0:0] sel);
    case (sel) 0: mux_5954 = 1'h0; 1: mux_5954 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5955;
  wire [0:0] v_5956;
  function [0:0] mux_5956(input [0:0] sel);
    case (sel) 0: mux_5956 = 1'h0; 1: mux_5956 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_5957;
  wire [0:0] v_5958;
  wire [0:0] v_5959;
  wire [0:0] v_5960;
  function [0:0] mux_5960(input [0:0] sel);
    case (sel) 0: mux_5960 = 1'h0; 1: mux_5960 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_5961;
  function [0:0] mux_5961(input [0:0] sel);
    case (sel) 0: mux_5961 = 1'h0; 1: mux_5961 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_5962 = 1'h0;
  wire [0:0] v_5963;
  wire [0:0] v_5964;
  wire [0:0] act_5965;
  wire [0:0] v_5966;
  wire [0:0] v_5967;
  wire [0:0] v_5968;
  reg [0:0] v_5969 = 1'h0;
  wire [0:0] v_5970;
  wire [0:0] v_5971;
  wire [0:0] act_5972;
  wire [0:0] v_5973;
  wire [0:0] v_5974;
  wire [0:0] v_5975;
  reg [0:0] v_5976 = 1'h0;
  wire [0:0] v_5977;
  wire [0:0] v_5978;
  wire [0:0] act_5979;
  wire [0:0] v_5980;
  wire [0:0] v_5981;
  wire [0:0] v_5982;
  reg [0:0] v_5983 = 1'h0;
  wire [0:0] v_5984;
  wire [0:0] v_5985;
  wire [0:0] act_5986;
  wire [0:0] v_5987;
  wire [0:0] v_5988;
  wire [0:0] v_5989;
  reg [0:0] v_5990 = 1'h0;
  wire [0:0] v_5991;
  wire [0:0] v_5992;
  wire [0:0] act_5993;
  wire [0:0] v_5994;
  wire [0:0] v_5995;
  wire [0:0] v_5996;
  wire [0:0] v_5997;
  wire [0:0] v_5998;
  wire [0:0] v_5999;
  function [0:0] mux_5999(input [0:0] sel);
    case (sel) 0: mux_5999 = 1'h0; 1: mux_5999 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6000;
  wire [0:0] v_6001;
  function [0:0] mux_6001(input [0:0] sel);
    case (sel) 0: mux_6001 = 1'h0; 1: mux_6001 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6002;
  wire [0:0] v_6003;
  wire [0:0] v_6004;
  wire [0:0] v_6005;
  function [0:0] mux_6005(input [0:0] sel);
    case (sel) 0: mux_6005 = 1'h0; 1: mux_6005 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6006;
  function [0:0] mux_6006(input [0:0] sel);
    case (sel) 0: mux_6006 = 1'h0; 1: mux_6006 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6007 = 1'h0;
  wire [0:0] v_6008;
  wire [0:0] v_6009;
  wire [0:0] act_6010;
  wire [0:0] v_6011;
  wire [0:0] v_6012;
  wire [0:0] v_6013;
  wire [0:0] v_6014;
  wire [0:0] v_6015;
  wire [0:0] v_6016;
  function [0:0] mux_6016(input [0:0] sel);
    case (sel) 0: mux_6016 = 1'h0; 1: mux_6016 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6017;
  function [0:0] mux_6017(input [0:0] sel);
    case (sel) 0: mux_6017 = 1'h0; 1: mux_6017 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6018;
  wire [0:0] v_6019;
  wire [0:0] v_6020;
  wire [0:0] v_6021;
  function [0:0] mux_6021(input [0:0] sel);
    case (sel) 0: mux_6021 = 1'h0; 1: mux_6021 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6022;
  function [0:0] mux_6022(input [0:0] sel);
    case (sel) 0: mux_6022 = 1'h0; 1: mux_6022 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6023;
  wire [0:0] v_6024;
  wire [0:0] v_6025;
  wire [0:0] v_6026;
  wire [0:0] v_6027;
  wire [0:0] v_6028;
  function [0:0] mux_6028(input [0:0] sel);
    case (sel) 0: mux_6028 = 1'h0; 1: mux_6028 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6029;
  wire [0:0] v_6030;
  function [0:0] mux_6030(input [0:0] sel);
    case (sel) 0: mux_6030 = 1'h0; 1: mux_6030 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6031;
  wire [0:0] v_6032;
  wire [0:0] v_6033;
  wire [0:0] v_6034;
  function [0:0] mux_6034(input [0:0] sel);
    case (sel) 0: mux_6034 = 1'h0; 1: mux_6034 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6035;
  function [0:0] mux_6035(input [0:0] sel);
    case (sel) 0: mux_6035 = 1'h0; 1: mux_6035 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6036 = 1'h0;
  wire [0:0] v_6037;
  wire [0:0] v_6038;
  wire [0:0] act_6039;
  wire [0:0] v_6040;
  wire [0:0] v_6041;
  wire [0:0] v_6042;
  reg [0:0] v_6043 = 1'h0;
  wire [0:0] v_6044;
  wire [0:0] v_6045;
  wire [0:0] act_6046;
  wire [0:0] v_6047;
  wire [0:0] v_6048;
  wire [0:0] v_6049;
  wire [0:0] v_6050;
  wire [0:0] v_6051;
  wire [0:0] v_6052;
  function [0:0] mux_6052(input [0:0] sel);
    case (sel) 0: mux_6052 = 1'h0; 1: mux_6052 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6053;
  wire [0:0] v_6054;
  function [0:0] mux_6054(input [0:0] sel);
    case (sel) 0: mux_6054 = 1'h0; 1: mux_6054 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6055;
  wire [0:0] v_6056;
  wire [0:0] v_6057;
  wire [0:0] v_6058;
  function [0:0] mux_6058(input [0:0] sel);
    case (sel) 0: mux_6058 = 1'h0; 1: mux_6058 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6059;
  function [0:0] mux_6059(input [0:0] sel);
    case (sel) 0: mux_6059 = 1'h0; 1: mux_6059 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6060 = 1'h0;
  wire [0:0] v_6061;
  wire [0:0] v_6062;
  wire [0:0] act_6063;
  wire [0:0] v_6064;
  wire [0:0] v_6065;
  wire [0:0] v_6066;
  wire [0:0] v_6067;
  wire [0:0] v_6068;
  wire [0:0] v_6069;
  function [0:0] mux_6069(input [0:0] sel);
    case (sel) 0: mux_6069 = 1'h0; 1: mux_6069 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6070;
  function [0:0] mux_6070(input [0:0] sel);
    case (sel) 0: mux_6070 = 1'h0; 1: mux_6070 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6071;
  wire [0:0] v_6072;
  wire [0:0] v_6073;
  wire [0:0] v_6074;
  function [0:0] mux_6074(input [0:0] sel);
    case (sel) 0: mux_6074 = 1'h0; 1: mux_6074 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6075;
  function [0:0] mux_6075(input [0:0] sel);
    case (sel) 0: mux_6075 = 1'h0; 1: mux_6075 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6076;
  wire [0:0] v_6077;
  wire [0:0] v_6078;
  wire [0:0] v_6079;
  wire [0:0] v_6080;
  wire [0:0] v_6081;
  function [0:0] mux_6081(input [0:0] sel);
    case (sel) 0: mux_6081 = 1'h0; 1: mux_6081 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6082;
  function [0:0] mux_6082(input [0:0] sel);
    case (sel) 0: mux_6082 = 1'h0; 1: mux_6082 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6083;
  wire [0:0] v_6084;
  wire [0:0] v_6085;
  wire [0:0] v_6086;
  function [0:0] mux_6086(input [0:0] sel);
    case (sel) 0: mux_6086 = 1'h0; 1: mux_6086 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6087;
  function [0:0] mux_6087(input [0:0] sel);
    case (sel) 0: mux_6087 = 1'h0; 1: mux_6087 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6088;
  wire [0:0] v_6089;
  wire [0:0] v_6090;
  wire [0:0] v_6091;
  wire [0:0] v_6092;
  wire [0:0] v_6093;
  function [0:0] mux_6093(input [0:0] sel);
    case (sel) 0: mux_6093 = 1'h0; 1: mux_6093 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6094;
  wire [0:0] v_6095;
  function [0:0] mux_6095(input [0:0] sel);
    case (sel) 0: mux_6095 = 1'h0; 1: mux_6095 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6096;
  wire [0:0] v_6097;
  wire [0:0] v_6098;
  wire [0:0] v_6099;
  function [0:0] mux_6099(input [0:0] sel);
    case (sel) 0: mux_6099 = 1'h0; 1: mux_6099 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6100;
  function [0:0] mux_6100(input [0:0] sel);
    case (sel) 0: mux_6100 = 1'h0; 1: mux_6100 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6101 = 1'h0;
  wire [0:0] v_6102;
  wire [0:0] v_6103;
  wire [0:0] act_6104;
  wire [0:0] v_6105;
  wire [0:0] v_6106;
  wire [0:0] v_6107;
  reg [0:0] v_6108 = 1'h0;
  wire [0:0] v_6109;
  wire [0:0] v_6110;
  wire [0:0] act_6111;
  wire [0:0] v_6112;
  wire [0:0] v_6113;
  wire [0:0] v_6114;
  reg [0:0] v_6115 = 1'h0;
  wire [0:0] v_6116;
  wire [0:0] v_6117;
  wire [0:0] act_6118;
  wire [0:0] v_6119;
  wire [0:0] v_6120;
  wire [0:0] v_6121;
  wire [0:0] v_6122;
  wire [0:0] v_6123;
  wire [0:0] v_6124;
  function [0:0] mux_6124(input [0:0] sel);
    case (sel) 0: mux_6124 = 1'h0; 1: mux_6124 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6125;
  wire [0:0] v_6126;
  function [0:0] mux_6126(input [0:0] sel);
    case (sel) 0: mux_6126 = 1'h0; 1: mux_6126 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6127;
  wire [0:0] v_6128;
  wire [0:0] v_6129;
  wire [0:0] v_6130;
  function [0:0] mux_6130(input [0:0] sel);
    case (sel) 0: mux_6130 = 1'h0; 1: mux_6130 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6131;
  function [0:0] mux_6131(input [0:0] sel);
    case (sel) 0: mux_6131 = 1'h0; 1: mux_6131 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6132 = 1'h0;
  wire [0:0] v_6133;
  wire [0:0] v_6134;
  wire [0:0] act_6135;
  wire [0:0] v_6136;
  wire [0:0] v_6137;
  wire [0:0] v_6138;
  wire [0:0] v_6139;
  wire [0:0] v_6140;
  wire [0:0] v_6141;
  function [0:0] mux_6141(input [0:0] sel);
    case (sel) 0: mux_6141 = 1'h0; 1: mux_6141 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6142;
  function [0:0] mux_6142(input [0:0] sel);
    case (sel) 0: mux_6142 = 1'h0; 1: mux_6142 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6143;
  wire [0:0] v_6144;
  wire [0:0] v_6145;
  wire [0:0] v_6146;
  function [0:0] mux_6146(input [0:0] sel);
    case (sel) 0: mux_6146 = 1'h0; 1: mux_6146 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6147;
  function [0:0] mux_6147(input [0:0] sel);
    case (sel) 0: mux_6147 = 1'h0; 1: mux_6147 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6148;
  wire [0:0] v_6149;
  wire [0:0] v_6150;
  wire [0:0] v_6151;
  wire [0:0] v_6152;
  wire [0:0] v_6153;
  function [0:0] mux_6153(input [0:0] sel);
    case (sel) 0: mux_6153 = 1'h0; 1: mux_6153 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6154;
  wire [0:0] v_6155;
  function [0:0] mux_6155(input [0:0] sel);
    case (sel) 0: mux_6155 = 1'h0; 1: mux_6155 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6156;
  wire [0:0] v_6157;
  wire [0:0] v_6158;
  wire [0:0] v_6159;
  function [0:0] mux_6159(input [0:0] sel);
    case (sel) 0: mux_6159 = 1'h0; 1: mux_6159 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6160;
  function [0:0] mux_6160(input [0:0] sel);
    case (sel) 0: mux_6160 = 1'h0; 1: mux_6160 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6161 = 1'h0;
  wire [0:0] v_6162;
  wire [0:0] v_6163;
  wire [0:0] act_6164;
  wire [0:0] v_6165;
  wire [0:0] v_6166;
  wire [0:0] v_6167;
  reg [0:0] v_6168 = 1'h0;
  wire [0:0] v_6169;
  wire [0:0] v_6170;
  wire [0:0] act_6171;
  wire [0:0] v_6172;
  wire [0:0] v_6173;
  wire [0:0] v_6174;
  wire [0:0] v_6175;
  wire [0:0] v_6176;
  wire [0:0] v_6177;
  function [0:0] mux_6177(input [0:0] sel);
    case (sel) 0: mux_6177 = 1'h0; 1: mux_6177 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6178;
  wire [0:0] v_6179;
  function [0:0] mux_6179(input [0:0] sel);
    case (sel) 0: mux_6179 = 1'h0; 1: mux_6179 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6180;
  wire [0:0] v_6181;
  wire [0:0] v_6182;
  wire [0:0] v_6183;
  function [0:0] mux_6183(input [0:0] sel);
    case (sel) 0: mux_6183 = 1'h0; 1: mux_6183 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6184;
  function [0:0] mux_6184(input [0:0] sel);
    case (sel) 0: mux_6184 = 1'h0; 1: mux_6184 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6185 = 1'h0;
  wire [0:0] v_6186;
  wire [0:0] v_6187;
  wire [0:0] act_6188;
  wire [0:0] v_6189;
  wire [0:0] v_6190;
  wire [0:0] v_6191;
  wire [0:0] v_6192;
  wire [0:0] v_6193;
  wire [0:0] v_6194;
  function [0:0] mux_6194(input [0:0] sel);
    case (sel) 0: mux_6194 = 1'h0; 1: mux_6194 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6195;
  function [0:0] mux_6195(input [0:0] sel);
    case (sel) 0: mux_6195 = 1'h0; 1: mux_6195 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6196;
  wire [0:0] v_6197;
  wire [0:0] v_6198;
  wire [0:0] v_6199;
  function [0:0] mux_6199(input [0:0] sel);
    case (sel) 0: mux_6199 = 1'h0; 1: mux_6199 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6200;
  function [0:0] mux_6200(input [0:0] sel);
    case (sel) 0: mux_6200 = 1'h0; 1: mux_6200 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6201;
  wire [0:0] v_6202;
  wire [0:0] v_6203;
  wire [0:0] v_6204;
  wire [0:0] v_6205;
  wire [0:0] v_6206;
  function [0:0] mux_6206(input [0:0] sel);
    case (sel) 0: mux_6206 = 1'h0; 1: mux_6206 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6207;
  function [0:0] mux_6207(input [0:0] sel);
    case (sel) 0: mux_6207 = 1'h0; 1: mux_6207 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6208;
  wire [0:0] v_6209;
  wire [0:0] v_6210;
  wire [0:0] v_6211;
  function [0:0] mux_6211(input [0:0] sel);
    case (sel) 0: mux_6211 = 1'h0; 1: mux_6211 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6212;
  function [0:0] mux_6212(input [0:0] sel);
    case (sel) 0: mux_6212 = 1'h0; 1: mux_6212 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6213;
  wire [0:0] v_6214;
  wire [0:0] v_6215;
  wire [0:0] v_6216;
  wire [0:0] v_6217;
  wire [0:0] v_6218;
  function [0:0] mux_6218(input [0:0] sel);
    case (sel) 0: mux_6218 = 1'h0; 1: mux_6218 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6219;
  function [0:0] mux_6219(input [0:0] sel);
    case (sel) 0: mux_6219 = 1'h0; 1: mux_6219 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6220;
  wire [0:0] v_6221;
  wire [0:0] v_6222;
  wire [0:0] v_6223;
  function [0:0] mux_6223(input [0:0] sel);
    case (sel) 0: mux_6223 = 1'h0; 1: mux_6223 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6224;
  function [0:0] mux_6224(input [0:0] sel);
    case (sel) 0: mux_6224 = 1'h0; 1: mux_6224 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6225;
  wire [0:0] v_6226;
  wire [0:0] v_6227;
  wire [0:0] v_6228;
  wire [0:0] v_6229;
  wire [0:0] v_6230;
  function [0:0] mux_6230(input [0:0] sel);
    case (sel) 0: mux_6230 = 1'h0; 1: mux_6230 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6231;
  wire [0:0] v_6232;
  function [0:0] mux_6232(input [0:0] sel);
    case (sel) 0: mux_6232 = 1'h0; 1: mux_6232 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6233;
  wire [0:0] v_6234;
  wire [0:0] v_6235;
  wire [0:0] v_6236;
  function [0:0] mux_6236(input [0:0] sel);
    case (sel) 0: mux_6236 = 1'h0; 1: mux_6236 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6237;
  function [0:0] mux_6237(input [0:0] sel);
    case (sel) 0: mux_6237 = 1'h0; 1: mux_6237 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6238 = 1'h0;
  wire [0:0] v_6239;
  wire [0:0] v_6240;
  wire [0:0] act_6241;
  wire [0:0] v_6242;
  wire [0:0] v_6243;
  wire [0:0] v_6244;
  reg [0:0] v_6245 = 1'h0;
  wire [0:0] v_6246;
  wire [0:0] v_6247;
  wire [0:0] act_6248;
  wire [0:0] v_6249;
  wire [0:0] v_6250;
  wire [0:0] v_6251;
  reg [0:0] v_6252 = 1'h0;
  wire [0:0] v_6253;
  wire [0:0] v_6254;
  wire [0:0] act_6255;
  wire [0:0] v_6256;
  wire [0:0] v_6257;
  wire [0:0] v_6258;
  reg [0:0] v_6259 = 1'h0;
  wire [0:0] v_6260;
  wire [0:0] v_6261;
  wire [0:0] act_6262;
  wire [0:0] v_6263;
  wire [0:0] v_6264;
  wire [0:0] v_6265;
  wire [0:0] v_6266;
  wire [0:0] v_6267;
  wire [0:0] v_6268;
  function [0:0] mux_6268(input [0:0] sel);
    case (sel) 0: mux_6268 = 1'h0; 1: mux_6268 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6269;
  wire [0:0] v_6270;
  function [0:0] mux_6270(input [0:0] sel);
    case (sel) 0: mux_6270 = 1'h0; 1: mux_6270 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6271;
  wire [0:0] v_6272;
  wire [0:0] v_6273;
  wire [0:0] v_6274;
  function [0:0] mux_6274(input [0:0] sel);
    case (sel) 0: mux_6274 = 1'h0; 1: mux_6274 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6275;
  function [0:0] mux_6275(input [0:0] sel);
    case (sel) 0: mux_6275 = 1'h0; 1: mux_6275 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6276 = 1'h0;
  wire [0:0] v_6277;
  wire [0:0] v_6278;
  wire [0:0] act_6279;
  wire [0:0] v_6280;
  wire [0:0] v_6281;
  wire [0:0] v_6282;
  wire [0:0] v_6283;
  wire [0:0] v_6284;
  wire [0:0] v_6285;
  function [0:0] mux_6285(input [0:0] sel);
    case (sel) 0: mux_6285 = 1'h0; 1: mux_6285 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6286;
  function [0:0] mux_6286(input [0:0] sel);
    case (sel) 0: mux_6286 = 1'h0; 1: mux_6286 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6287;
  wire [0:0] v_6288;
  wire [0:0] v_6289;
  wire [0:0] v_6290;
  function [0:0] mux_6290(input [0:0] sel);
    case (sel) 0: mux_6290 = 1'h0; 1: mux_6290 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6291;
  function [0:0] mux_6291(input [0:0] sel);
    case (sel) 0: mux_6291 = 1'h0; 1: mux_6291 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6292;
  wire [0:0] v_6293;
  wire [0:0] v_6294;
  wire [0:0] v_6295;
  wire [0:0] v_6296;
  wire [0:0] v_6297;
  function [0:0] mux_6297(input [0:0] sel);
    case (sel) 0: mux_6297 = 1'h0; 1: mux_6297 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6298;
  wire [0:0] v_6299;
  function [0:0] mux_6299(input [0:0] sel);
    case (sel) 0: mux_6299 = 1'h0; 1: mux_6299 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6300;
  wire [0:0] v_6301;
  wire [0:0] v_6302;
  wire [0:0] v_6303;
  function [0:0] mux_6303(input [0:0] sel);
    case (sel) 0: mux_6303 = 1'h0; 1: mux_6303 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6304;
  function [0:0] mux_6304(input [0:0] sel);
    case (sel) 0: mux_6304 = 1'h0; 1: mux_6304 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6305 = 1'h0;
  wire [0:0] v_6306;
  wire [0:0] v_6307;
  wire [0:0] act_6308;
  wire [0:0] v_6309;
  wire [0:0] v_6310;
  wire [0:0] v_6311;
  reg [0:0] v_6312 = 1'h0;
  wire [0:0] v_6313;
  wire [0:0] v_6314;
  wire [0:0] act_6315;
  wire [0:0] v_6316;
  wire [0:0] v_6317;
  wire [0:0] v_6318;
  wire [0:0] v_6319;
  wire [0:0] v_6320;
  wire [0:0] v_6321;
  function [0:0] mux_6321(input [0:0] sel);
    case (sel) 0: mux_6321 = 1'h0; 1: mux_6321 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6322;
  wire [0:0] v_6323;
  function [0:0] mux_6323(input [0:0] sel);
    case (sel) 0: mux_6323 = 1'h0; 1: mux_6323 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6324;
  wire [0:0] v_6325;
  wire [0:0] v_6326;
  wire [0:0] v_6327;
  function [0:0] mux_6327(input [0:0] sel);
    case (sel) 0: mux_6327 = 1'h0; 1: mux_6327 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6328;
  function [0:0] mux_6328(input [0:0] sel);
    case (sel) 0: mux_6328 = 1'h0; 1: mux_6328 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6329 = 1'h0;
  wire [0:0] v_6330;
  wire [0:0] v_6331;
  wire [0:0] act_6332;
  wire [0:0] v_6333;
  wire [0:0] v_6334;
  wire [0:0] v_6335;
  wire [0:0] v_6336;
  wire [0:0] v_6337;
  wire [0:0] v_6338;
  function [0:0] mux_6338(input [0:0] sel);
    case (sel) 0: mux_6338 = 1'h0; 1: mux_6338 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6339;
  function [0:0] mux_6339(input [0:0] sel);
    case (sel) 0: mux_6339 = 1'h0; 1: mux_6339 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6340;
  wire [0:0] v_6341;
  wire [0:0] v_6342;
  wire [0:0] v_6343;
  function [0:0] mux_6343(input [0:0] sel);
    case (sel) 0: mux_6343 = 1'h0; 1: mux_6343 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6344;
  function [0:0] mux_6344(input [0:0] sel);
    case (sel) 0: mux_6344 = 1'h0; 1: mux_6344 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6345;
  wire [0:0] v_6346;
  wire [0:0] v_6347;
  wire [0:0] v_6348;
  wire [0:0] v_6349;
  wire [0:0] v_6350;
  function [0:0] mux_6350(input [0:0] sel);
    case (sel) 0: mux_6350 = 1'h0; 1: mux_6350 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6351;
  function [0:0] mux_6351(input [0:0] sel);
    case (sel) 0: mux_6351 = 1'h0; 1: mux_6351 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6352;
  wire [0:0] v_6353;
  wire [0:0] v_6354;
  wire [0:0] v_6355;
  function [0:0] mux_6355(input [0:0] sel);
    case (sel) 0: mux_6355 = 1'h0; 1: mux_6355 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6356;
  function [0:0] mux_6356(input [0:0] sel);
    case (sel) 0: mux_6356 = 1'h0; 1: mux_6356 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6357;
  wire [0:0] v_6358;
  wire [0:0] v_6359;
  wire [0:0] v_6360;
  wire [0:0] v_6361;
  wire [0:0] v_6362;
  function [0:0] mux_6362(input [0:0] sel);
    case (sel) 0: mux_6362 = 1'h0; 1: mux_6362 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6363;
  wire [0:0] v_6364;
  function [0:0] mux_6364(input [0:0] sel);
    case (sel) 0: mux_6364 = 1'h0; 1: mux_6364 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6365;
  wire [0:0] v_6366;
  wire [0:0] v_6367;
  wire [0:0] v_6368;
  function [0:0] mux_6368(input [0:0] sel);
    case (sel) 0: mux_6368 = 1'h0; 1: mux_6368 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6369;
  function [0:0] mux_6369(input [0:0] sel);
    case (sel) 0: mux_6369 = 1'h0; 1: mux_6369 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6370 = 1'h0;
  wire [0:0] v_6371;
  wire [0:0] v_6372;
  wire [0:0] act_6373;
  wire [0:0] v_6374;
  wire [0:0] v_6375;
  wire [0:0] v_6376;
  reg [0:0] v_6377 = 1'h0;
  wire [0:0] v_6378;
  wire [0:0] v_6379;
  wire [0:0] act_6380;
  wire [0:0] v_6381;
  wire [0:0] v_6382;
  wire [0:0] v_6383;
  reg [0:0] v_6384 = 1'h0;
  wire [0:0] v_6385;
  wire [0:0] v_6386;
  wire [0:0] act_6387;
  wire [0:0] v_6388;
  wire [0:0] v_6389;
  wire [0:0] v_6390;
  wire [0:0] v_6391;
  wire [0:0] v_6392;
  wire [0:0] v_6393;
  function [0:0] mux_6393(input [0:0] sel);
    case (sel) 0: mux_6393 = 1'h0; 1: mux_6393 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6394;
  wire [0:0] v_6395;
  function [0:0] mux_6395(input [0:0] sel);
    case (sel) 0: mux_6395 = 1'h0; 1: mux_6395 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6396;
  wire [0:0] v_6397;
  wire [0:0] v_6398;
  wire [0:0] v_6399;
  function [0:0] mux_6399(input [0:0] sel);
    case (sel) 0: mux_6399 = 1'h0; 1: mux_6399 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6400;
  function [0:0] mux_6400(input [0:0] sel);
    case (sel) 0: mux_6400 = 1'h0; 1: mux_6400 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6401 = 1'h0;
  wire [0:0] v_6402;
  wire [0:0] v_6403;
  wire [0:0] act_6404;
  wire [0:0] v_6405;
  wire [0:0] v_6406;
  wire [0:0] v_6407;
  wire [0:0] v_6408;
  wire [0:0] v_6409;
  wire [0:0] v_6410;
  function [0:0] mux_6410(input [0:0] sel);
    case (sel) 0: mux_6410 = 1'h0; 1: mux_6410 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6411;
  function [0:0] mux_6411(input [0:0] sel);
    case (sel) 0: mux_6411 = 1'h0; 1: mux_6411 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6412;
  wire [0:0] v_6413;
  wire [0:0] v_6414;
  wire [0:0] v_6415;
  function [0:0] mux_6415(input [0:0] sel);
    case (sel) 0: mux_6415 = 1'h0; 1: mux_6415 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6416;
  function [0:0] mux_6416(input [0:0] sel);
    case (sel) 0: mux_6416 = 1'h0; 1: mux_6416 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6417;
  wire [0:0] v_6418;
  wire [0:0] v_6419;
  wire [0:0] v_6420;
  wire [0:0] v_6421;
  wire [0:0] v_6422;
  function [0:0] mux_6422(input [0:0] sel);
    case (sel) 0: mux_6422 = 1'h0; 1: mux_6422 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6423;
  wire [0:0] v_6424;
  function [0:0] mux_6424(input [0:0] sel);
    case (sel) 0: mux_6424 = 1'h0; 1: mux_6424 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6425;
  wire [0:0] v_6426;
  wire [0:0] v_6427;
  wire [0:0] v_6428;
  function [0:0] mux_6428(input [0:0] sel);
    case (sel) 0: mux_6428 = 1'h0; 1: mux_6428 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6429;
  function [0:0] mux_6429(input [0:0] sel);
    case (sel) 0: mux_6429 = 1'h0; 1: mux_6429 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6430 = 1'h0;
  wire [0:0] v_6431;
  wire [0:0] v_6432;
  wire [0:0] act_6433;
  wire [0:0] v_6434;
  wire [0:0] v_6435;
  wire [0:0] v_6436;
  reg [0:0] v_6437 = 1'h0;
  wire [0:0] v_6438;
  wire [0:0] v_6439;
  wire [0:0] act_6440;
  wire [0:0] v_6441;
  wire [0:0] v_6442;
  wire [0:0] v_6443;
  wire [0:0] v_6444;
  wire [0:0] v_6445;
  wire [0:0] v_6446;
  function [0:0] mux_6446(input [0:0] sel);
    case (sel) 0: mux_6446 = 1'h0; 1: mux_6446 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6447;
  wire [0:0] v_6448;
  function [0:0] mux_6448(input [0:0] sel);
    case (sel) 0: mux_6448 = 1'h0; 1: mux_6448 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6449;
  wire [0:0] v_6450;
  wire [0:0] v_6451;
  wire [0:0] v_6452;
  function [0:0] mux_6452(input [0:0] sel);
    case (sel) 0: mux_6452 = 1'h0; 1: mux_6452 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6453;
  function [0:0] mux_6453(input [0:0] sel);
    case (sel) 0: mux_6453 = 1'h0; 1: mux_6453 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6454 = 1'h0;
  wire [0:0] v_6455;
  wire [0:0] v_6456;
  wire [0:0] act_6457;
  wire [0:0] v_6458;
  wire [0:0] v_6459;
  wire [0:0] v_6460;
  wire [0:0] v_6461;
  wire [0:0] v_6462;
  wire [0:0] v_6463;
  function [0:0] mux_6463(input [0:0] sel);
    case (sel) 0: mux_6463 = 1'h0; 1: mux_6463 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6464;
  function [0:0] mux_6464(input [0:0] sel);
    case (sel) 0: mux_6464 = 1'h0; 1: mux_6464 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6465;
  wire [0:0] v_6466;
  wire [0:0] v_6467;
  wire [0:0] v_6468;
  function [0:0] mux_6468(input [0:0] sel);
    case (sel) 0: mux_6468 = 1'h0; 1: mux_6468 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6469;
  function [0:0] mux_6469(input [0:0] sel);
    case (sel) 0: mux_6469 = 1'h0; 1: mux_6469 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6470;
  wire [0:0] v_6471;
  wire [0:0] v_6472;
  wire [0:0] v_6473;
  wire [0:0] v_6474;
  wire [0:0] v_6475;
  function [0:0] mux_6475(input [0:0] sel);
    case (sel) 0: mux_6475 = 1'h0; 1: mux_6475 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6476;
  function [0:0] mux_6476(input [0:0] sel);
    case (sel) 0: mux_6476 = 1'h0; 1: mux_6476 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6477;
  wire [0:0] v_6478;
  wire [0:0] v_6479;
  wire [0:0] v_6480;
  function [0:0] mux_6480(input [0:0] sel);
    case (sel) 0: mux_6480 = 1'h0; 1: mux_6480 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6481;
  function [0:0] mux_6481(input [0:0] sel);
    case (sel) 0: mux_6481 = 1'h0; 1: mux_6481 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6482;
  wire [0:0] v_6483;
  wire [0:0] v_6484;
  wire [0:0] v_6485;
  wire [0:0] v_6486;
  wire [0:0] v_6487;
  function [0:0] mux_6487(input [0:0] sel);
    case (sel) 0: mux_6487 = 1'h0; 1: mux_6487 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6488;
  function [0:0] mux_6488(input [0:0] sel);
    case (sel) 0: mux_6488 = 1'h0; 1: mux_6488 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6489;
  wire [0:0] v_6490;
  wire [0:0] v_6491;
  wire [0:0] v_6492;
  function [0:0] mux_6492(input [0:0] sel);
    case (sel) 0: mux_6492 = 1'h0; 1: mux_6492 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6493;
  function [0:0] mux_6493(input [0:0] sel);
    case (sel) 0: mux_6493 = 1'h0; 1: mux_6493 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6494;
  wire [0:0] v_6495;
  wire [0:0] v_6496;
  wire [0:0] v_6497;
  wire [0:0] v_6498;
  wire [0:0] v_6499;
  function [0:0] mux_6499(input [0:0] sel);
    case (sel) 0: mux_6499 = 1'h0; 1: mux_6499 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6500;
  function [0:0] mux_6500(input [0:0] sel);
    case (sel) 0: mux_6500 = 1'h0; 1: mux_6500 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6501;
  wire [0:0] v_6502;
  wire [0:0] v_6503;
  wire [0:0] v_6504;
  function [0:0] mux_6504(input [0:0] sel);
    case (sel) 0: mux_6504 = 1'h0; 1: mux_6504 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6505;
  function [0:0] mux_6505(input [0:0] sel);
    case (sel) 0: mux_6505 = 1'h0; 1: mux_6505 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6506;
  wire [0:0] v_6507;
  wire [0:0] v_6508;
  wire [0:0] v_6509;
  wire [0:0] v_6510;
  wire [0:0] v_6511;
  function [0:0] mux_6511(input [0:0] sel);
    case (sel) 0: mux_6511 = 1'h0; 1: mux_6511 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6512;
  function [0:0] mux_6512(input [0:0] sel);
    case (sel) 0: mux_6512 = 1'h0; 1: mux_6512 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6513;
  wire [0:0] v_6514;
  wire [0:0] v_6515;
  wire [0:0] v_6516;
  function [0:0] mux_6516(input [0:0] sel);
    case (sel) 0: mux_6516 = 1'h0; 1: mux_6516 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6517;
  function [0:0] mux_6517(input [0:0] sel);
    case (sel) 0: mux_6517 = 1'h0; 1: mux_6517 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6518;
  wire [0:0] v_6519;
  wire [0:0] v_6520;
  wire [0:0] v_6521;
  wire [0:0] v_6522;
  wire [0:0] v_6523;
  function [0:0] mux_6523(input [0:0] sel);
    case (sel) 0: mux_6523 = 1'h0; 1: mux_6523 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6524;
  wire [0:0] v_6525;
  function [0:0] mux_6525(input [0:0] sel);
    case (sel) 0: mux_6525 = 1'h0; 1: mux_6525 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6526;
  wire [0:0] v_6527;
  wire [0:0] v_6528;
  wire [0:0] v_6529;
  function [0:0] mux_6529(input [0:0] sel);
    case (sel) 0: mux_6529 = 1'h0; 1: mux_6529 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6530;
  function [0:0] mux_6530(input [0:0] sel);
    case (sel) 0: mux_6530 = 1'h0; 1: mux_6530 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6531 = 1'h0;
  wire [0:0] v_6532;
  wire [0:0] v_6533;
  wire [0:0] act_6534;
  wire [0:0] v_6535;
  wire [0:0] v_6536;
  wire [0:0] v_6537;
  reg [0:0] v_6538 = 1'h0;
  wire [0:0] v_6539;
  wire [0:0] v_6540;
  wire [0:0] act_6541;
  wire [0:0] v_6542;
  wire [0:0] v_6543;
  wire [0:0] v_6544;
  reg [0:0] v_6545 = 1'h0;
  wire [0:0] v_6546;
  wire [0:0] v_6547;
  wire [0:0] act_6548;
  wire [0:0] v_6549;
  wire [0:0] v_6550;
  wire [0:0] v_6551;
  reg [0:0] v_6552 = 1'h0;
  wire [0:0] v_6553;
  wire [0:0] v_6554;
  wire [0:0] act_6555;
  wire [0:0] v_6556;
  wire [0:0] v_6557;
  wire [0:0] v_6558;
  reg [0:0] v_6559 = 1'h0;
  wire [0:0] v_6560;
  wire [0:0] v_6561;
  wire [0:0] act_6562;
  wire [0:0] v_6563;
  wire [0:0] v_6564;
  wire [0:0] v_6565;
  reg [0:0] v_6566 = 1'h0;
  wire [0:0] v_6567;
  wire [0:0] v_6568;
  wire [0:0] act_6569;
  wire [0:0] v_6570;
  wire [0:0] v_6571;
  wire [0:0] v_6572;
  wire [0:0] v_6573;
  wire [0:0] v_6574;
  wire [0:0] v_6575;
  function [0:0] mux_6575(input [0:0] sel);
    case (sel) 0: mux_6575 = 1'h0; 1: mux_6575 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6576;
  wire [0:0] v_6577;
  function [0:0] mux_6577(input [0:0] sel);
    case (sel) 0: mux_6577 = 1'h0; 1: mux_6577 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6578;
  wire [0:0] v_6579;
  wire [0:0] v_6580;
  wire [0:0] v_6581;
  function [0:0] mux_6581(input [0:0] sel);
    case (sel) 0: mux_6581 = 1'h0; 1: mux_6581 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6582;
  function [0:0] mux_6582(input [0:0] sel);
    case (sel) 0: mux_6582 = 1'h0; 1: mux_6582 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6583 = 1'h0;
  wire [0:0] v_6584;
  wire [0:0] v_6585;
  wire [0:0] act_6586;
  wire [0:0] v_6587;
  wire [0:0] v_6588;
  wire [0:0] v_6589;
  wire [0:0] v_6590;
  wire [0:0] v_6591;
  wire [0:0] v_6592;
  function [0:0] mux_6592(input [0:0] sel);
    case (sel) 0: mux_6592 = 1'h0; 1: mux_6592 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6593;
  function [0:0] mux_6593(input [0:0] sel);
    case (sel) 0: mux_6593 = 1'h0; 1: mux_6593 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6594;
  wire [0:0] v_6595;
  wire [0:0] v_6596;
  wire [0:0] v_6597;
  function [0:0] mux_6597(input [0:0] sel);
    case (sel) 0: mux_6597 = 1'h0; 1: mux_6597 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6598;
  function [0:0] mux_6598(input [0:0] sel);
    case (sel) 0: mux_6598 = 1'h0; 1: mux_6598 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6599;
  wire [0:0] v_6600;
  wire [0:0] v_6601;
  wire [0:0] v_6602;
  wire [0:0] v_6603;
  wire [0:0] v_6604;
  function [0:0] mux_6604(input [0:0] sel);
    case (sel) 0: mux_6604 = 1'h0; 1: mux_6604 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6605;
  wire [0:0] v_6606;
  function [0:0] mux_6606(input [0:0] sel);
    case (sel) 0: mux_6606 = 1'h0; 1: mux_6606 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6607;
  wire [0:0] v_6608;
  wire [0:0] v_6609;
  wire [0:0] v_6610;
  function [0:0] mux_6610(input [0:0] sel);
    case (sel) 0: mux_6610 = 1'h0; 1: mux_6610 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6611;
  function [0:0] mux_6611(input [0:0] sel);
    case (sel) 0: mux_6611 = 1'h0; 1: mux_6611 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6612 = 1'h0;
  wire [0:0] v_6613;
  wire [0:0] v_6614;
  wire [0:0] act_6615;
  wire [0:0] v_6616;
  wire [0:0] v_6617;
  wire [0:0] v_6618;
  reg [0:0] v_6619 = 1'h0;
  wire [0:0] v_6620;
  wire [0:0] v_6621;
  wire [0:0] act_6622;
  wire [0:0] v_6623;
  wire [0:0] v_6624;
  wire [0:0] v_6625;
  wire [0:0] v_6626;
  wire [0:0] v_6627;
  wire [0:0] v_6628;
  function [0:0] mux_6628(input [0:0] sel);
    case (sel) 0: mux_6628 = 1'h0; 1: mux_6628 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6629;
  wire [0:0] v_6630;
  function [0:0] mux_6630(input [0:0] sel);
    case (sel) 0: mux_6630 = 1'h0; 1: mux_6630 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6631;
  wire [0:0] v_6632;
  wire [0:0] v_6633;
  wire [0:0] v_6634;
  function [0:0] mux_6634(input [0:0] sel);
    case (sel) 0: mux_6634 = 1'h0; 1: mux_6634 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6635;
  function [0:0] mux_6635(input [0:0] sel);
    case (sel) 0: mux_6635 = 1'h0; 1: mux_6635 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6636 = 1'h0;
  wire [0:0] v_6637;
  wire [0:0] v_6638;
  wire [0:0] act_6639;
  wire [0:0] v_6640;
  wire [0:0] v_6641;
  wire [0:0] v_6642;
  wire [0:0] v_6643;
  wire [0:0] v_6644;
  wire [0:0] v_6645;
  function [0:0] mux_6645(input [0:0] sel);
    case (sel) 0: mux_6645 = 1'h0; 1: mux_6645 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6646;
  function [0:0] mux_6646(input [0:0] sel);
    case (sel) 0: mux_6646 = 1'h0; 1: mux_6646 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6647;
  wire [0:0] v_6648;
  wire [0:0] v_6649;
  wire [0:0] v_6650;
  function [0:0] mux_6650(input [0:0] sel);
    case (sel) 0: mux_6650 = 1'h0; 1: mux_6650 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6651;
  function [0:0] mux_6651(input [0:0] sel);
    case (sel) 0: mux_6651 = 1'h0; 1: mux_6651 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6652;
  wire [0:0] v_6653;
  wire [0:0] v_6654;
  wire [0:0] v_6655;
  wire [0:0] v_6656;
  wire [0:0] v_6657;
  function [0:0] mux_6657(input [0:0] sel);
    case (sel) 0: mux_6657 = 1'h0; 1: mux_6657 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6658;
  function [0:0] mux_6658(input [0:0] sel);
    case (sel) 0: mux_6658 = 1'h0; 1: mux_6658 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6659;
  wire [0:0] v_6660;
  wire [0:0] v_6661;
  wire [0:0] v_6662;
  function [0:0] mux_6662(input [0:0] sel);
    case (sel) 0: mux_6662 = 1'h0; 1: mux_6662 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6663;
  function [0:0] mux_6663(input [0:0] sel);
    case (sel) 0: mux_6663 = 1'h0; 1: mux_6663 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6664;
  wire [0:0] v_6665;
  wire [0:0] v_6666;
  wire [0:0] v_6667;
  wire [0:0] v_6668;
  wire [0:0] v_6669;
  function [0:0] mux_6669(input [0:0] sel);
    case (sel) 0: mux_6669 = 1'h0; 1: mux_6669 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6670;
  wire [0:0] v_6671;
  function [0:0] mux_6671(input [0:0] sel);
    case (sel) 0: mux_6671 = 1'h0; 1: mux_6671 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6672;
  wire [0:0] v_6673;
  wire [0:0] v_6674;
  wire [0:0] v_6675;
  function [0:0] mux_6675(input [0:0] sel);
    case (sel) 0: mux_6675 = 1'h0; 1: mux_6675 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6676;
  function [0:0] mux_6676(input [0:0] sel);
    case (sel) 0: mux_6676 = 1'h0; 1: mux_6676 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6677 = 1'h0;
  wire [0:0] v_6678;
  wire [0:0] v_6679;
  wire [0:0] act_6680;
  wire [0:0] v_6681;
  wire [0:0] v_6682;
  wire [0:0] v_6683;
  reg [0:0] v_6684 = 1'h0;
  wire [0:0] v_6685;
  wire [0:0] v_6686;
  wire [0:0] act_6687;
  wire [0:0] v_6688;
  wire [0:0] v_6689;
  wire [0:0] v_6690;
  reg [0:0] v_6691 = 1'h0;
  wire [0:0] v_6692;
  wire [0:0] v_6693;
  wire [0:0] act_6694;
  wire [0:0] v_6695;
  wire [0:0] v_6696;
  wire [0:0] v_6697;
  wire [0:0] v_6698;
  wire [0:0] v_6699;
  wire [0:0] v_6700;
  function [0:0] mux_6700(input [0:0] sel);
    case (sel) 0: mux_6700 = 1'h0; 1: mux_6700 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6701;
  wire [0:0] v_6702;
  function [0:0] mux_6702(input [0:0] sel);
    case (sel) 0: mux_6702 = 1'h0; 1: mux_6702 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6703;
  wire [0:0] v_6704;
  wire [0:0] v_6705;
  wire [0:0] v_6706;
  function [0:0] mux_6706(input [0:0] sel);
    case (sel) 0: mux_6706 = 1'h0; 1: mux_6706 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6707;
  function [0:0] mux_6707(input [0:0] sel);
    case (sel) 0: mux_6707 = 1'h0; 1: mux_6707 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6708 = 1'h0;
  wire [0:0] v_6709;
  wire [0:0] v_6710;
  wire [0:0] act_6711;
  wire [0:0] v_6712;
  wire [0:0] v_6713;
  wire [0:0] v_6714;
  wire [0:0] v_6715;
  wire [0:0] v_6716;
  wire [0:0] v_6717;
  function [0:0] mux_6717(input [0:0] sel);
    case (sel) 0: mux_6717 = 1'h0; 1: mux_6717 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6718;
  function [0:0] mux_6718(input [0:0] sel);
    case (sel) 0: mux_6718 = 1'h0; 1: mux_6718 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6719;
  wire [0:0] v_6720;
  wire [0:0] v_6721;
  wire [0:0] v_6722;
  function [0:0] mux_6722(input [0:0] sel);
    case (sel) 0: mux_6722 = 1'h0; 1: mux_6722 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6723;
  function [0:0] mux_6723(input [0:0] sel);
    case (sel) 0: mux_6723 = 1'h0; 1: mux_6723 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6724;
  wire [0:0] v_6725;
  wire [0:0] v_6726;
  wire [0:0] v_6727;
  wire [0:0] v_6728;
  wire [0:0] v_6729;
  function [0:0] mux_6729(input [0:0] sel);
    case (sel) 0: mux_6729 = 1'h0; 1: mux_6729 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6730;
  wire [0:0] v_6731;
  function [0:0] mux_6731(input [0:0] sel);
    case (sel) 0: mux_6731 = 1'h0; 1: mux_6731 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6732;
  wire [0:0] v_6733;
  wire [0:0] v_6734;
  wire [0:0] v_6735;
  function [0:0] mux_6735(input [0:0] sel);
    case (sel) 0: mux_6735 = 1'h0; 1: mux_6735 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6736;
  function [0:0] mux_6736(input [0:0] sel);
    case (sel) 0: mux_6736 = 1'h0; 1: mux_6736 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6737 = 1'h0;
  wire [0:0] v_6738;
  wire [0:0] v_6739;
  wire [0:0] act_6740;
  wire [0:0] v_6741;
  wire [0:0] v_6742;
  wire [0:0] v_6743;
  reg [0:0] v_6744 = 1'h0;
  wire [0:0] v_6745;
  wire [0:0] v_6746;
  wire [0:0] act_6747;
  wire [0:0] v_6748;
  wire [0:0] v_6749;
  wire [0:0] v_6750;
  wire [0:0] v_6751;
  wire [0:0] v_6752;
  wire [0:0] v_6753;
  function [0:0] mux_6753(input [0:0] sel);
    case (sel) 0: mux_6753 = 1'h0; 1: mux_6753 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6754;
  wire [0:0] v_6755;
  function [0:0] mux_6755(input [0:0] sel);
    case (sel) 0: mux_6755 = 1'h0; 1: mux_6755 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6756;
  wire [0:0] v_6757;
  wire [0:0] v_6758;
  wire [0:0] v_6759;
  function [0:0] mux_6759(input [0:0] sel);
    case (sel) 0: mux_6759 = 1'h0; 1: mux_6759 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6760;
  function [0:0] mux_6760(input [0:0] sel);
    case (sel) 0: mux_6760 = 1'h0; 1: mux_6760 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6761 = 1'h0;
  wire [0:0] v_6762;
  wire [0:0] v_6763;
  wire [0:0] act_6764;
  wire [0:0] v_6765;
  wire [0:0] v_6766;
  wire [0:0] v_6767;
  wire [0:0] v_6768;
  wire [0:0] v_6769;
  wire [0:0] v_6770;
  function [0:0] mux_6770(input [0:0] sel);
    case (sel) 0: mux_6770 = 1'h0; 1: mux_6770 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6771;
  function [0:0] mux_6771(input [0:0] sel);
    case (sel) 0: mux_6771 = 1'h0; 1: mux_6771 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6772;
  wire [0:0] v_6773;
  wire [0:0] v_6774;
  wire [0:0] v_6775;
  function [0:0] mux_6775(input [0:0] sel);
    case (sel) 0: mux_6775 = 1'h0; 1: mux_6775 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6776;
  function [0:0] mux_6776(input [0:0] sel);
    case (sel) 0: mux_6776 = 1'h0; 1: mux_6776 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6777;
  wire [0:0] v_6778;
  wire [0:0] v_6779;
  wire [0:0] v_6780;
  wire [0:0] v_6781;
  wire [0:0] v_6782;
  function [0:0] mux_6782(input [0:0] sel);
    case (sel) 0: mux_6782 = 1'h0; 1: mux_6782 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6783;
  function [0:0] mux_6783(input [0:0] sel);
    case (sel) 0: mux_6783 = 1'h0; 1: mux_6783 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6784;
  wire [0:0] v_6785;
  wire [0:0] v_6786;
  wire [0:0] v_6787;
  function [0:0] mux_6787(input [0:0] sel);
    case (sel) 0: mux_6787 = 1'h0; 1: mux_6787 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6788;
  function [0:0] mux_6788(input [0:0] sel);
    case (sel) 0: mux_6788 = 1'h0; 1: mux_6788 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6789;
  wire [0:0] v_6790;
  wire [0:0] v_6791;
  wire [0:0] v_6792;
  wire [0:0] v_6793;
  wire [0:0] v_6794;
  function [0:0] mux_6794(input [0:0] sel);
    case (sel) 0: mux_6794 = 1'h0; 1: mux_6794 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6795;
  function [0:0] mux_6795(input [0:0] sel);
    case (sel) 0: mux_6795 = 1'h0; 1: mux_6795 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6796;
  wire [0:0] v_6797;
  wire [0:0] v_6798;
  wire [0:0] v_6799;
  function [0:0] mux_6799(input [0:0] sel);
    case (sel) 0: mux_6799 = 1'h0; 1: mux_6799 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6800;
  function [0:0] mux_6800(input [0:0] sel);
    case (sel) 0: mux_6800 = 1'h0; 1: mux_6800 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6801;
  wire [0:0] v_6802;
  wire [0:0] v_6803;
  wire [0:0] v_6804;
  wire [0:0] v_6805;
  wire [0:0] v_6806;
  function [0:0] mux_6806(input [0:0] sel);
    case (sel) 0: mux_6806 = 1'h0; 1: mux_6806 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6807;
  wire [0:0] v_6808;
  function [0:0] mux_6808(input [0:0] sel);
    case (sel) 0: mux_6808 = 1'h0; 1: mux_6808 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6809;
  wire [0:0] v_6810;
  wire [0:0] v_6811;
  wire [0:0] v_6812;
  function [0:0] mux_6812(input [0:0] sel);
    case (sel) 0: mux_6812 = 1'h0; 1: mux_6812 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6813;
  function [0:0] mux_6813(input [0:0] sel);
    case (sel) 0: mux_6813 = 1'h0; 1: mux_6813 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6814 = 1'h0;
  wire [0:0] v_6815;
  wire [0:0] v_6816;
  wire [0:0] act_6817;
  wire [0:0] v_6818;
  wire [0:0] v_6819;
  wire [0:0] v_6820;
  reg [0:0] v_6821 = 1'h0;
  wire [0:0] v_6822;
  wire [0:0] v_6823;
  wire [0:0] act_6824;
  wire [0:0] v_6825;
  wire [0:0] v_6826;
  wire [0:0] v_6827;
  reg [0:0] v_6828 = 1'h0;
  wire [0:0] v_6829;
  wire [0:0] v_6830;
  wire [0:0] act_6831;
  wire [0:0] v_6832;
  wire [0:0] v_6833;
  wire [0:0] v_6834;
  reg [0:0] v_6835 = 1'h0;
  wire [0:0] v_6836;
  wire [0:0] v_6837;
  wire [0:0] act_6838;
  wire [0:0] v_6839;
  wire [0:0] v_6840;
  wire [0:0] v_6841;
  wire [0:0] v_6842;
  wire [0:0] v_6843;
  wire [0:0] v_6844;
  function [0:0] mux_6844(input [0:0] sel);
    case (sel) 0: mux_6844 = 1'h0; 1: mux_6844 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6845;
  wire [0:0] v_6846;
  function [0:0] mux_6846(input [0:0] sel);
    case (sel) 0: mux_6846 = 1'h0; 1: mux_6846 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6847;
  wire [0:0] v_6848;
  wire [0:0] v_6849;
  wire [0:0] v_6850;
  function [0:0] mux_6850(input [0:0] sel);
    case (sel) 0: mux_6850 = 1'h0; 1: mux_6850 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6851;
  function [0:0] mux_6851(input [0:0] sel);
    case (sel) 0: mux_6851 = 1'h0; 1: mux_6851 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6852 = 1'h0;
  wire [0:0] v_6853;
  wire [0:0] v_6854;
  wire [0:0] act_6855;
  wire [0:0] v_6856;
  wire [0:0] v_6857;
  wire [0:0] v_6858;
  wire [0:0] v_6859;
  wire [0:0] v_6860;
  wire [0:0] v_6861;
  function [0:0] mux_6861(input [0:0] sel);
    case (sel) 0: mux_6861 = 1'h0; 1: mux_6861 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6862;
  function [0:0] mux_6862(input [0:0] sel);
    case (sel) 0: mux_6862 = 1'h0; 1: mux_6862 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6863;
  wire [0:0] v_6864;
  wire [0:0] v_6865;
  wire [0:0] v_6866;
  function [0:0] mux_6866(input [0:0] sel);
    case (sel) 0: mux_6866 = 1'h0; 1: mux_6866 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6867;
  function [0:0] mux_6867(input [0:0] sel);
    case (sel) 0: mux_6867 = 1'h0; 1: mux_6867 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6868;
  wire [0:0] v_6869;
  wire [0:0] v_6870;
  wire [0:0] v_6871;
  wire [0:0] v_6872;
  wire [0:0] v_6873;
  function [0:0] mux_6873(input [0:0] sel);
    case (sel) 0: mux_6873 = 1'h0; 1: mux_6873 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6874;
  wire [0:0] v_6875;
  function [0:0] mux_6875(input [0:0] sel);
    case (sel) 0: mux_6875 = 1'h0; 1: mux_6875 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6876;
  wire [0:0] v_6877;
  wire [0:0] v_6878;
  wire [0:0] v_6879;
  function [0:0] mux_6879(input [0:0] sel);
    case (sel) 0: mux_6879 = 1'h0; 1: mux_6879 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6880;
  function [0:0] mux_6880(input [0:0] sel);
    case (sel) 0: mux_6880 = 1'h0; 1: mux_6880 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6881 = 1'h0;
  wire [0:0] v_6882;
  wire [0:0] v_6883;
  wire [0:0] act_6884;
  wire [0:0] v_6885;
  wire [0:0] v_6886;
  wire [0:0] v_6887;
  reg [0:0] v_6888 = 1'h0;
  wire [0:0] v_6889;
  wire [0:0] v_6890;
  wire [0:0] act_6891;
  wire [0:0] v_6892;
  wire [0:0] v_6893;
  wire [0:0] v_6894;
  wire [0:0] v_6895;
  wire [0:0] v_6896;
  wire [0:0] v_6897;
  function [0:0] mux_6897(input [0:0] sel);
    case (sel) 0: mux_6897 = 1'h0; 1: mux_6897 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6898;
  wire [0:0] v_6899;
  function [0:0] mux_6899(input [0:0] sel);
    case (sel) 0: mux_6899 = 1'h0; 1: mux_6899 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6900;
  wire [0:0] v_6901;
  wire [0:0] v_6902;
  wire [0:0] v_6903;
  function [0:0] mux_6903(input [0:0] sel);
    case (sel) 0: mux_6903 = 1'h0; 1: mux_6903 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6904;
  function [0:0] mux_6904(input [0:0] sel);
    case (sel) 0: mux_6904 = 1'h0; 1: mux_6904 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6905 = 1'h0;
  wire [0:0] v_6906;
  wire [0:0] v_6907;
  wire [0:0] act_6908;
  wire [0:0] v_6909;
  wire [0:0] v_6910;
  wire [0:0] v_6911;
  wire [0:0] v_6912;
  wire [0:0] v_6913;
  wire [0:0] v_6914;
  function [0:0] mux_6914(input [0:0] sel);
    case (sel) 0: mux_6914 = 1'h0; 1: mux_6914 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6915;
  function [0:0] mux_6915(input [0:0] sel);
    case (sel) 0: mux_6915 = 1'h0; 1: mux_6915 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6916;
  wire [0:0] v_6917;
  wire [0:0] v_6918;
  wire [0:0] v_6919;
  function [0:0] mux_6919(input [0:0] sel);
    case (sel) 0: mux_6919 = 1'h0; 1: mux_6919 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6920;
  function [0:0] mux_6920(input [0:0] sel);
    case (sel) 0: mux_6920 = 1'h0; 1: mux_6920 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6921;
  wire [0:0] v_6922;
  wire [0:0] v_6923;
  wire [0:0] v_6924;
  wire [0:0] v_6925;
  wire [0:0] v_6926;
  function [0:0] mux_6926(input [0:0] sel);
    case (sel) 0: mux_6926 = 1'h0; 1: mux_6926 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6927;
  function [0:0] mux_6927(input [0:0] sel);
    case (sel) 0: mux_6927 = 1'h0; 1: mux_6927 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6928;
  wire [0:0] v_6929;
  wire [0:0] v_6930;
  wire [0:0] v_6931;
  function [0:0] mux_6931(input [0:0] sel);
    case (sel) 0: mux_6931 = 1'h0; 1: mux_6931 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6932;
  function [0:0] mux_6932(input [0:0] sel);
    case (sel) 0: mux_6932 = 1'h0; 1: mux_6932 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6933;
  wire [0:0] v_6934;
  wire [0:0] v_6935;
  wire [0:0] v_6936;
  wire [0:0] v_6937;
  wire [0:0] v_6938;
  function [0:0] mux_6938(input [0:0] sel);
    case (sel) 0: mux_6938 = 1'h0; 1: mux_6938 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6939;
  wire [0:0] v_6940;
  function [0:0] mux_6940(input [0:0] sel);
    case (sel) 0: mux_6940 = 1'h0; 1: mux_6940 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6941;
  wire [0:0] v_6942;
  wire [0:0] v_6943;
  wire [0:0] v_6944;
  function [0:0] mux_6944(input [0:0] sel);
    case (sel) 0: mux_6944 = 1'h0; 1: mux_6944 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6945;
  function [0:0] mux_6945(input [0:0] sel);
    case (sel) 0: mux_6945 = 1'h0; 1: mux_6945 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6946 = 1'h0;
  wire [0:0] v_6947;
  wire [0:0] v_6948;
  wire [0:0] act_6949;
  wire [0:0] v_6950;
  wire [0:0] v_6951;
  wire [0:0] v_6952;
  reg [0:0] v_6953 = 1'h0;
  wire [0:0] v_6954;
  wire [0:0] v_6955;
  wire [0:0] act_6956;
  wire [0:0] v_6957;
  wire [0:0] v_6958;
  wire [0:0] v_6959;
  reg [0:0] v_6960 = 1'h0;
  wire [0:0] v_6961;
  wire [0:0] v_6962;
  wire [0:0] act_6963;
  wire [0:0] v_6964;
  wire [0:0] v_6965;
  wire [0:0] v_6966;
  wire [0:0] v_6967;
  wire [0:0] v_6968;
  wire [0:0] v_6969;
  function [0:0] mux_6969(input [0:0] sel);
    case (sel) 0: mux_6969 = 1'h0; 1: mux_6969 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6970;
  wire [0:0] v_6971;
  function [0:0] mux_6971(input [0:0] sel);
    case (sel) 0: mux_6971 = 1'h0; 1: mux_6971 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6972;
  wire [0:0] v_6973;
  wire [0:0] v_6974;
  wire [0:0] v_6975;
  function [0:0] mux_6975(input [0:0] sel);
    case (sel) 0: mux_6975 = 1'h0; 1: mux_6975 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6976;
  function [0:0] mux_6976(input [0:0] sel);
    case (sel) 0: mux_6976 = 1'h0; 1: mux_6976 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_6977 = 1'h0;
  wire [0:0] v_6978;
  wire [0:0] v_6979;
  wire [0:0] act_6980;
  wire [0:0] v_6981;
  wire [0:0] v_6982;
  wire [0:0] v_6983;
  wire [0:0] v_6984;
  wire [0:0] v_6985;
  wire [0:0] v_6986;
  function [0:0] mux_6986(input [0:0] sel);
    case (sel) 0: mux_6986 = 1'h0; 1: mux_6986 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6987;
  function [0:0] mux_6987(input [0:0] sel);
    case (sel) 0: mux_6987 = 1'h0; 1: mux_6987 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6988;
  wire [0:0] v_6989;
  wire [0:0] v_6990;
  wire [0:0] v_6991;
  function [0:0] mux_6991(input [0:0] sel);
    case (sel) 0: mux_6991 = 1'h0; 1: mux_6991 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6992;
  function [0:0] mux_6992(input [0:0] sel);
    case (sel) 0: mux_6992 = 1'h0; 1: mux_6992 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_6993;
  wire [0:0] v_6994;
  wire [0:0] v_6995;
  wire [0:0] v_6996;
  wire [0:0] v_6997;
  wire [0:0] v_6998;
  function [0:0] mux_6998(input [0:0] sel);
    case (sel) 0: mux_6998 = 1'h0; 1: mux_6998 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_6999;
  wire [0:0] v_7000;
  function [0:0] mux_7000(input [0:0] sel);
    case (sel) 0: mux_7000 = 1'h0; 1: mux_7000 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7001;
  wire [0:0] v_7002;
  wire [0:0] v_7003;
  wire [0:0] v_7004;
  function [0:0] mux_7004(input [0:0] sel);
    case (sel) 0: mux_7004 = 1'h0; 1: mux_7004 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7005;
  function [0:0] mux_7005(input [0:0] sel);
    case (sel) 0: mux_7005 = 1'h0; 1: mux_7005 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7006 = 1'h0;
  wire [0:0] v_7007;
  wire [0:0] v_7008;
  wire [0:0] act_7009;
  wire [0:0] v_7010;
  wire [0:0] v_7011;
  wire [0:0] v_7012;
  reg [0:0] v_7013 = 1'h0;
  wire [0:0] v_7014;
  wire [0:0] v_7015;
  wire [0:0] act_7016;
  wire [0:0] v_7017;
  wire [0:0] v_7018;
  wire [0:0] v_7019;
  wire [0:0] v_7020;
  wire [0:0] v_7021;
  wire [0:0] v_7022;
  function [0:0] mux_7022(input [0:0] sel);
    case (sel) 0: mux_7022 = 1'h0; 1: mux_7022 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7023;
  wire [0:0] v_7024;
  function [0:0] mux_7024(input [0:0] sel);
    case (sel) 0: mux_7024 = 1'h0; 1: mux_7024 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7025;
  wire [0:0] v_7026;
  wire [0:0] v_7027;
  wire [0:0] v_7028;
  function [0:0] mux_7028(input [0:0] sel);
    case (sel) 0: mux_7028 = 1'h0; 1: mux_7028 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7029;
  function [0:0] mux_7029(input [0:0] sel);
    case (sel) 0: mux_7029 = 1'h0; 1: mux_7029 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7030 = 1'h0;
  wire [0:0] v_7031;
  wire [0:0] v_7032;
  wire [0:0] act_7033;
  wire [0:0] v_7034;
  wire [0:0] v_7035;
  wire [0:0] v_7036;
  wire [0:0] v_7037;
  wire [0:0] v_7038;
  wire [0:0] v_7039;
  function [0:0] mux_7039(input [0:0] sel);
    case (sel) 0: mux_7039 = 1'h0; 1: mux_7039 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7040;
  function [0:0] mux_7040(input [0:0] sel);
    case (sel) 0: mux_7040 = 1'h0; 1: mux_7040 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7041;
  wire [0:0] v_7042;
  wire [0:0] v_7043;
  wire [0:0] v_7044;
  function [0:0] mux_7044(input [0:0] sel);
    case (sel) 0: mux_7044 = 1'h0; 1: mux_7044 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7045;
  function [0:0] mux_7045(input [0:0] sel);
    case (sel) 0: mux_7045 = 1'h0; 1: mux_7045 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7046;
  wire [0:0] v_7047;
  wire [0:0] v_7048;
  wire [0:0] v_7049;
  wire [0:0] v_7050;
  wire [0:0] v_7051;
  function [0:0] mux_7051(input [0:0] sel);
    case (sel) 0: mux_7051 = 1'h0; 1: mux_7051 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7052;
  function [0:0] mux_7052(input [0:0] sel);
    case (sel) 0: mux_7052 = 1'h0; 1: mux_7052 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7053;
  wire [0:0] v_7054;
  wire [0:0] v_7055;
  wire [0:0] v_7056;
  function [0:0] mux_7056(input [0:0] sel);
    case (sel) 0: mux_7056 = 1'h0; 1: mux_7056 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7057;
  function [0:0] mux_7057(input [0:0] sel);
    case (sel) 0: mux_7057 = 1'h0; 1: mux_7057 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7058;
  wire [0:0] v_7059;
  wire [0:0] v_7060;
  wire [0:0] v_7061;
  wire [0:0] v_7062;
  wire [0:0] v_7063;
  function [0:0] mux_7063(input [0:0] sel);
    case (sel) 0: mux_7063 = 1'h0; 1: mux_7063 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7064;
  function [0:0] mux_7064(input [0:0] sel);
    case (sel) 0: mux_7064 = 1'h0; 1: mux_7064 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7065;
  wire [0:0] v_7066;
  wire [0:0] v_7067;
  wire [0:0] v_7068;
  function [0:0] mux_7068(input [0:0] sel);
    case (sel) 0: mux_7068 = 1'h0; 1: mux_7068 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7069;
  function [0:0] mux_7069(input [0:0] sel);
    case (sel) 0: mux_7069 = 1'h0; 1: mux_7069 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7070;
  wire [0:0] v_7071;
  wire [0:0] v_7072;
  wire [0:0] v_7073;
  wire [0:0] v_7074;
  wire [0:0] v_7075;
  function [0:0] mux_7075(input [0:0] sel);
    case (sel) 0: mux_7075 = 1'h0; 1: mux_7075 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7076;
  function [0:0] mux_7076(input [0:0] sel);
    case (sel) 0: mux_7076 = 1'h0; 1: mux_7076 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7077;
  wire [0:0] v_7078;
  wire [0:0] v_7079;
  wire [0:0] v_7080;
  function [0:0] mux_7080(input [0:0] sel);
    case (sel) 0: mux_7080 = 1'h0; 1: mux_7080 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7081;
  function [0:0] mux_7081(input [0:0] sel);
    case (sel) 0: mux_7081 = 1'h0; 1: mux_7081 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7082;
  wire [0:0] v_7083;
  wire [0:0] v_7084;
  wire [0:0] v_7085;
  wire [0:0] v_7086;
  wire [0:0] v_7087;
  function [0:0] mux_7087(input [0:0] sel);
    case (sel) 0: mux_7087 = 1'h0; 1: mux_7087 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7088;
  wire [0:0] v_7089;
  function [0:0] mux_7089(input [0:0] sel);
    case (sel) 0: mux_7089 = 1'h0; 1: mux_7089 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7090;
  wire [0:0] v_7091;
  wire [0:0] v_7092;
  wire [0:0] v_7093;
  function [0:0] mux_7093(input [0:0] sel);
    case (sel) 0: mux_7093 = 1'h0; 1: mux_7093 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7094;
  function [0:0] mux_7094(input [0:0] sel);
    case (sel) 0: mux_7094 = 1'h0; 1: mux_7094 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7095 = 1'h0;
  wire [0:0] v_7096;
  wire [0:0] v_7097;
  wire [0:0] act_7098;
  wire [0:0] v_7099;
  wire [0:0] v_7100;
  wire [0:0] v_7101;
  reg [0:0] v_7102 = 1'h0;
  wire [0:0] v_7103;
  wire [0:0] v_7104;
  wire [0:0] act_7105;
  wire [0:0] v_7106;
  wire [0:0] v_7107;
  wire [0:0] v_7108;
  reg [0:0] v_7109 = 1'h0;
  wire [0:0] v_7110;
  wire [0:0] v_7111;
  wire [0:0] act_7112;
  wire [0:0] v_7113;
  wire [0:0] v_7114;
  wire [0:0] v_7115;
  reg [0:0] v_7116 = 1'h0;
  wire [0:0] v_7117;
  wire [0:0] v_7118;
  wire [0:0] act_7119;
  wire [0:0] v_7120;
  wire [0:0] v_7121;
  wire [0:0] v_7122;
  reg [0:0] v_7123 = 1'h0;
  wire [0:0] v_7124;
  wire [0:0] v_7125;
  wire [0:0] act_7126;
  wire [0:0] v_7127;
  wire [0:0] v_7128;
  wire [0:0] v_7129;
  wire [0:0] v_7130;
  wire [0:0] v_7131;
  wire [0:0] v_7132;
  function [0:0] mux_7132(input [0:0] sel);
    case (sel) 0: mux_7132 = 1'h0; 1: mux_7132 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7133;
  wire [0:0] v_7134;
  function [0:0] mux_7134(input [0:0] sel);
    case (sel) 0: mux_7134 = 1'h0; 1: mux_7134 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7135;
  wire [0:0] v_7136;
  wire [0:0] v_7137;
  wire [0:0] v_7138;
  function [0:0] mux_7138(input [0:0] sel);
    case (sel) 0: mux_7138 = 1'h0; 1: mux_7138 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7139;
  function [0:0] mux_7139(input [0:0] sel);
    case (sel) 0: mux_7139 = 1'h0; 1: mux_7139 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7140 = 1'h0;
  wire [0:0] v_7141;
  wire [0:0] v_7142;
  wire [0:0] act_7143;
  wire [0:0] v_7144;
  wire [0:0] v_7145;
  wire [0:0] v_7146;
  wire [0:0] v_7147;
  wire [0:0] v_7148;
  wire [0:0] v_7149;
  function [0:0] mux_7149(input [0:0] sel);
    case (sel) 0: mux_7149 = 1'h0; 1: mux_7149 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7150;
  function [0:0] mux_7150(input [0:0] sel);
    case (sel) 0: mux_7150 = 1'h0; 1: mux_7150 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7151;
  wire [0:0] v_7152;
  wire [0:0] v_7153;
  wire [0:0] v_7154;
  function [0:0] mux_7154(input [0:0] sel);
    case (sel) 0: mux_7154 = 1'h0; 1: mux_7154 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7155;
  function [0:0] mux_7155(input [0:0] sel);
    case (sel) 0: mux_7155 = 1'h0; 1: mux_7155 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7156;
  wire [0:0] v_7157;
  wire [0:0] v_7158;
  wire [0:0] v_7159;
  wire [0:0] v_7160;
  wire [0:0] v_7161;
  function [0:0] mux_7161(input [0:0] sel);
    case (sel) 0: mux_7161 = 1'h0; 1: mux_7161 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7162;
  wire [0:0] v_7163;
  function [0:0] mux_7163(input [0:0] sel);
    case (sel) 0: mux_7163 = 1'h0; 1: mux_7163 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7164;
  wire [0:0] v_7165;
  wire [0:0] v_7166;
  wire [0:0] v_7167;
  function [0:0] mux_7167(input [0:0] sel);
    case (sel) 0: mux_7167 = 1'h0; 1: mux_7167 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7168;
  function [0:0] mux_7168(input [0:0] sel);
    case (sel) 0: mux_7168 = 1'h0; 1: mux_7168 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7169 = 1'h0;
  wire [0:0] v_7170;
  wire [0:0] v_7171;
  wire [0:0] act_7172;
  wire [0:0] v_7173;
  wire [0:0] v_7174;
  wire [0:0] v_7175;
  reg [0:0] v_7176 = 1'h0;
  wire [0:0] v_7177;
  wire [0:0] v_7178;
  wire [0:0] act_7179;
  wire [0:0] v_7180;
  wire [0:0] v_7181;
  wire [0:0] v_7182;
  wire [0:0] v_7183;
  wire [0:0] v_7184;
  wire [0:0] v_7185;
  function [0:0] mux_7185(input [0:0] sel);
    case (sel) 0: mux_7185 = 1'h0; 1: mux_7185 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7186;
  wire [0:0] v_7187;
  function [0:0] mux_7187(input [0:0] sel);
    case (sel) 0: mux_7187 = 1'h0; 1: mux_7187 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7188;
  wire [0:0] v_7189;
  wire [0:0] v_7190;
  wire [0:0] v_7191;
  function [0:0] mux_7191(input [0:0] sel);
    case (sel) 0: mux_7191 = 1'h0; 1: mux_7191 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7192;
  function [0:0] mux_7192(input [0:0] sel);
    case (sel) 0: mux_7192 = 1'h0; 1: mux_7192 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7193 = 1'h0;
  wire [0:0] v_7194;
  wire [0:0] v_7195;
  wire [0:0] act_7196;
  wire [0:0] v_7197;
  wire [0:0] v_7198;
  wire [0:0] v_7199;
  wire [0:0] v_7200;
  wire [0:0] v_7201;
  wire [0:0] v_7202;
  function [0:0] mux_7202(input [0:0] sel);
    case (sel) 0: mux_7202 = 1'h0; 1: mux_7202 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7203;
  function [0:0] mux_7203(input [0:0] sel);
    case (sel) 0: mux_7203 = 1'h0; 1: mux_7203 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7204;
  wire [0:0] v_7205;
  wire [0:0] v_7206;
  wire [0:0] v_7207;
  function [0:0] mux_7207(input [0:0] sel);
    case (sel) 0: mux_7207 = 1'h0; 1: mux_7207 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7208;
  function [0:0] mux_7208(input [0:0] sel);
    case (sel) 0: mux_7208 = 1'h0; 1: mux_7208 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7209;
  wire [0:0] v_7210;
  wire [0:0] v_7211;
  wire [0:0] v_7212;
  wire [0:0] v_7213;
  wire [0:0] v_7214;
  function [0:0] mux_7214(input [0:0] sel);
    case (sel) 0: mux_7214 = 1'h0; 1: mux_7214 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7215;
  function [0:0] mux_7215(input [0:0] sel);
    case (sel) 0: mux_7215 = 1'h0; 1: mux_7215 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7216;
  wire [0:0] v_7217;
  wire [0:0] v_7218;
  wire [0:0] v_7219;
  function [0:0] mux_7219(input [0:0] sel);
    case (sel) 0: mux_7219 = 1'h0; 1: mux_7219 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7220;
  function [0:0] mux_7220(input [0:0] sel);
    case (sel) 0: mux_7220 = 1'h0; 1: mux_7220 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7221;
  wire [0:0] v_7222;
  wire [0:0] v_7223;
  wire [0:0] v_7224;
  wire [0:0] v_7225;
  wire [0:0] v_7226;
  function [0:0] mux_7226(input [0:0] sel);
    case (sel) 0: mux_7226 = 1'h0; 1: mux_7226 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7227;
  wire [0:0] v_7228;
  function [0:0] mux_7228(input [0:0] sel);
    case (sel) 0: mux_7228 = 1'h0; 1: mux_7228 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7229;
  wire [0:0] v_7230;
  wire [0:0] v_7231;
  wire [0:0] v_7232;
  function [0:0] mux_7232(input [0:0] sel);
    case (sel) 0: mux_7232 = 1'h0; 1: mux_7232 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7233;
  function [0:0] mux_7233(input [0:0] sel);
    case (sel) 0: mux_7233 = 1'h0; 1: mux_7233 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7234 = 1'h0;
  wire [0:0] v_7235;
  wire [0:0] v_7236;
  wire [0:0] act_7237;
  wire [0:0] v_7238;
  wire [0:0] v_7239;
  wire [0:0] v_7240;
  reg [0:0] v_7241 = 1'h0;
  wire [0:0] v_7242;
  wire [0:0] v_7243;
  wire [0:0] act_7244;
  wire [0:0] v_7245;
  wire [0:0] v_7246;
  wire [0:0] v_7247;
  reg [0:0] v_7248 = 1'h0;
  wire [0:0] v_7249;
  wire [0:0] v_7250;
  wire [0:0] act_7251;
  wire [0:0] v_7252;
  wire [0:0] v_7253;
  wire [0:0] v_7254;
  wire [0:0] v_7255;
  wire [0:0] v_7256;
  wire [0:0] v_7257;
  function [0:0] mux_7257(input [0:0] sel);
    case (sel) 0: mux_7257 = 1'h0; 1: mux_7257 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7258;
  wire [0:0] v_7259;
  function [0:0] mux_7259(input [0:0] sel);
    case (sel) 0: mux_7259 = 1'h0; 1: mux_7259 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7260;
  wire [0:0] v_7261;
  wire [0:0] v_7262;
  wire [0:0] v_7263;
  function [0:0] mux_7263(input [0:0] sel);
    case (sel) 0: mux_7263 = 1'h0; 1: mux_7263 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7264;
  function [0:0] mux_7264(input [0:0] sel);
    case (sel) 0: mux_7264 = 1'h0; 1: mux_7264 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7265 = 1'h0;
  wire [0:0] v_7266;
  wire [0:0] v_7267;
  wire [0:0] act_7268;
  wire [0:0] v_7269;
  wire [0:0] v_7270;
  wire [0:0] v_7271;
  wire [0:0] v_7272;
  wire [0:0] v_7273;
  wire [0:0] v_7274;
  function [0:0] mux_7274(input [0:0] sel);
    case (sel) 0: mux_7274 = 1'h0; 1: mux_7274 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7275;
  function [0:0] mux_7275(input [0:0] sel);
    case (sel) 0: mux_7275 = 1'h0; 1: mux_7275 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7276;
  wire [0:0] v_7277;
  wire [0:0] v_7278;
  wire [0:0] v_7279;
  function [0:0] mux_7279(input [0:0] sel);
    case (sel) 0: mux_7279 = 1'h0; 1: mux_7279 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7280;
  function [0:0] mux_7280(input [0:0] sel);
    case (sel) 0: mux_7280 = 1'h0; 1: mux_7280 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7281;
  wire [0:0] v_7282;
  wire [0:0] v_7283;
  wire [0:0] v_7284;
  wire [0:0] v_7285;
  wire [0:0] v_7286;
  function [0:0] mux_7286(input [0:0] sel);
    case (sel) 0: mux_7286 = 1'h0; 1: mux_7286 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7287;
  wire [0:0] v_7288;
  function [0:0] mux_7288(input [0:0] sel);
    case (sel) 0: mux_7288 = 1'h0; 1: mux_7288 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7289;
  wire [0:0] v_7290;
  wire [0:0] v_7291;
  wire [0:0] v_7292;
  function [0:0] mux_7292(input [0:0] sel);
    case (sel) 0: mux_7292 = 1'h0; 1: mux_7292 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7293;
  function [0:0] mux_7293(input [0:0] sel);
    case (sel) 0: mux_7293 = 1'h0; 1: mux_7293 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7294 = 1'h0;
  wire [0:0] v_7295;
  wire [0:0] v_7296;
  wire [0:0] act_7297;
  wire [0:0] v_7298;
  wire [0:0] v_7299;
  wire [0:0] v_7300;
  reg [0:0] v_7301 = 1'h0;
  wire [0:0] v_7302;
  wire [0:0] v_7303;
  wire [0:0] act_7304;
  wire [0:0] v_7305;
  wire [0:0] v_7306;
  wire [0:0] v_7307;
  wire [0:0] v_7308;
  wire [0:0] v_7309;
  wire [0:0] v_7310;
  function [0:0] mux_7310(input [0:0] sel);
    case (sel) 0: mux_7310 = 1'h0; 1: mux_7310 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7311;
  wire [0:0] v_7312;
  function [0:0] mux_7312(input [0:0] sel);
    case (sel) 0: mux_7312 = 1'h0; 1: mux_7312 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7313;
  wire [0:0] v_7314;
  wire [0:0] v_7315;
  wire [0:0] v_7316;
  function [0:0] mux_7316(input [0:0] sel);
    case (sel) 0: mux_7316 = 1'h0; 1: mux_7316 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7317;
  function [0:0] mux_7317(input [0:0] sel);
    case (sel) 0: mux_7317 = 1'h0; 1: mux_7317 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7318 = 1'h0;
  wire [0:0] v_7319;
  wire [0:0] v_7320;
  wire [0:0] act_7321;
  wire [0:0] v_7322;
  wire [0:0] v_7323;
  wire [0:0] v_7324;
  wire [0:0] v_7325;
  wire [0:0] v_7326;
  wire [0:0] v_7327;
  function [0:0] mux_7327(input [0:0] sel);
    case (sel) 0: mux_7327 = 1'h0; 1: mux_7327 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7328;
  function [0:0] mux_7328(input [0:0] sel);
    case (sel) 0: mux_7328 = 1'h0; 1: mux_7328 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7329;
  wire [0:0] v_7330;
  wire [0:0] v_7331;
  wire [0:0] v_7332;
  function [0:0] mux_7332(input [0:0] sel);
    case (sel) 0: mux_7332 = 1'h0; 1: mux_7332 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7333;
  function [0:0] mux_7333(input [0:0] sel);
    case (sel) 0: mux_7333 = 1'h0; 1: mux_7333 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7334;
  wire [0:0] v_7335;
  wire [0:0] v_7336;
  wire [0:0] v_7337;
  wire [0:0] v_7338;
  wire [0:0] v_7339;
  function [0:0] mux_7339(input [0:0] sel);
    case (sel) 0: mux_7339 = 1'h0; 1: mux_7339 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7340;
  function [0:0] mux_7340(input [0:0] sel);
    case (sel) 0: mux_7340 = 1'h0; 1: mux_7340 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7341;
  wire [0:0] v_7342;
  wire [0:0] v_7343;
  wire [0:0] v_7344;
  function [0:0] mux_7344(input [0:0] sel);
    case (sel) 0: mux_7344 = 1'h0; 1: mux_7344 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7345;
  function [0:0] mux_7345(input [0:0] sel);
    case (sel) 0: mux_7345 = 1'h0; 1: mux_7345 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7346;
  wire [0:0] v_7347;
  wire [0:0] v_7348;
  wire [0:0] v_7349;
  wire [0:0] v_7350;
  wire [0:0] v_7351;
  function [0:0] mux_7351(input [0:0] sel);
    case (sel) 0: mux_7351 = 1'h0; 1: mux_7351 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7352;
  function [0:0] mux_7352(input [0:0] sel);
    case (sel) 0: mux_7352 = 1'h0; 1: mux_7352 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7353;
  wire [0:0] v_7354;
  wire [0:0] v_7355;
  wire [0:0] v_7356;
  function [0:0] mux_7356(input [0:0] sel);
    case (sel) 0: mux_7356 = 1'h0; 1: mux_7356 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7357;
  function [0:0] mux_7357(input [0:0] sel);
    case (sel) 0: mux_7357 = 1'h0; 1: mux_7357 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7358;
  wire [0:0] v_7359;
  wire [0:0] v_7360;
  wire [0:0] v_7361;
  wire [0:0] v_7362;
  wire [0:0] v_7363;
  function [0:0] mux_7363(input [0:0] sel);
    case (sel) 0: mux_7363 = 1'h0; 1: mux_7363 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7364;
  wire [0:0] v_7365;
  function [0:0] mux_7365(input [0:0] sel);
    case (sel) 0: mux_7365 = 1'h0; 1: mux_7365 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7366;
  wire [0:0] v_7367;
  wire [0:0] v_7368;
  wire [0:0] v_7369;
  function [0:0] mux_7369(input [0:0] sel);
    case (sel) 0: mux_7369 = 1'h0; 1: mux_7369 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7370;
  function [0:0] mux_7370(input [0:0] sel);
    case (sel) 0: mux_7370 = 1'h0; 1: mux_7370 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7371 = 1'h0;
  wire [0:0] v_7372;
  wire [0:0] v_7373;
  wire [0:0] act_7374;
  wire [0:0] v_7375;
  wire [0:0] v_7376;
  wire [0:0] v_7377;
  reg [0:0] v_7378 = 1'h0;
  wire [0:0] v_7379;
  wire [0:0] v_7380;
  wire [0:0] act_7381;
  wire [0:0] v_7382;
  wire [0:0] v_7383;
  wire [0:0] v_7384;
  reg [0:0] v_7385 = 1'h0;
  wire [0:0] v_7386;
  wire [0:0] v_7387;
  wire [0:0] act_7388;
  wire [0:0] v_7389;
  wire [0:0] v_7390;
  wire [0:0] v_7391;
  reg [0:0] v_7392 = 1'h0;
  wire [0:0] v_7393;
  wire [0:0] v_7394;
  wire [0:0] act_7395;
  wire [0:0] v_7396;
  wire [0:0] v_7397;
  wire [0:0] v_7398;
  wire [0:0] v_7399;
  wire [0:0] v_7400;
  wire [0:0] v_7401;
  function [0:0] mux_7401(input [0:0] sel);
    case (sel) 0: mux_7401 = 1'h0; 1: mux_7401 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7402;
  wire [0:0] v_7403;
  function [0:0] mux_7403(input [0:0] sel);
    case (sel) 0: mux_7403 = 1'h0; 1: mux_7403 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7404;
  wire [0:0] v_7405;
  wire [0:0] v_7406;
  wire [0:0] v_7407;
  function [0:0] mux_7407(input [0:0] sel);
    case (sel) 0: mux_7407 = 1'h0; 1: mux_7407 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7408;
  function [0:0] mux_7408(input [0:0] sel);
    case (sel) 0: mux_7408 = 1'h0; 1: mux_7408 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7409 = 1'h0;
  wire [0:0] v_7410;
  wire [0:0] v_7411;
  wire [0:0] act_7412;
  wire [0:0] v_7413;
  wire [0:0] v_7414;
  wire [0:0] v_7415;
  wire [0:0] v_7416;
  wire [0:0] v_7417;
  wire [0:0] v_7418;
  function [0:0] mux_7418(input [0:0] sel);
    case (sel) 0: mux_7418 = 1'h0; 1: mux_7418 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7419;
  function [0:0] mux_7419(input [0:0] sel);
    case (sel) 0: mux_7419 = 1'h0; 1: mux_7419 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7420;
  wire [0:0] v_7421;
  wire [0:0] v_7422;
  wire [0:0] v_7423;
  function [0:0] mux_7423(input [0:0] sel);
    case (sel) 0: mux_7423 = 1'h0; 1: mux_7423 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7424;
  function [0:0] mux_7424(input [0:0] sel);
    case (sel) 0: mux_7424 = 1'h0; 1: mux_7424 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7425;
  wire [0:0] v_7426;
  wire [0:0] v_7427;
  wire [0:0] v_7428;
  wire [0:0] v_7429;
  wire [0:0] v_7430;
  function [0:0] mux_7430(input [0:0] sel);
    case (sel) 0: mux_7430 = 1'h0; 1: mux_7430 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7431;
  wire [0:0] v_7432;
  function [0:0] mux_7432(input [0:0] sel);
    case (sel) 0: mux_7432 = 1'h0; 1: mux_7432 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7433;
  wire [0:0] v_7434;
  wire [0:0] v_7435;
  wire [0:0] v_7436;
  function [0:0] mux_7436(input [0:0] sel);
    case (sel) 0: mux_7436 = 1'h0; 1: mux_7436 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7437;
  function [0:0] mux_7437(input [0:0] sel);
    case (sel) 0: mux_7437 = 1'h0; 1: mux_7437 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7438 = 1'h0;
  wire [0:0] v_7439;
  wire [0:0] v_7440;
  wire [0:0] act_7441;
  wire [0:0] v_7442;
  wire [0:0] v_7443;
  wire [0:0] v_7444;
  reg [0:0] v_7445 = 1'h0;
  wire [0:0] v_7446;
  wire [0:0] v_7447;
  wire [0:0] act_7448;
  wire [0:0] v_7449;
  wire [0:0] v_7450;
  wire [0:0] v_7451;
  wire [0:0] v_7452;
  wire [0:0] v_7453;
  wire [0:0] v_7454;
  function [0:0] mux_7454(input [0:0] sel);
    case (sel) 0: mux_7454 = 1'h0; 1: mux_7454 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7455;
  wire [0:0] v_7456;
  function [0:0] mux_7456(input [0:0] sel);
    case (sel) 0: mux_7456 = 1'h0; 1: mux_7456 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7457;
  wire [0:0] v_7458;
  wire [0:0] v_7459;
  wire [0:0] v_7460;
  function [0:0] mux_7460(input [0:0] sel);
    case (sel) 0: mux_7460 = 1'h0; 1: mux_7460 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7461;
  function [0:0] mux_7461(input [0:0] sel);
    case (sel) 0: mux_7461 = 1'h0; 1: mux_7461 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7462 = 1'h0;
  wire [0:0] v_7463;
  wire [0:0] v_7464;
  wire [0:0] act_7465;
  wire [0:0] v_7466;
  wire [0:0] v_7467;
  wire [0:0] v_7468;
  wire [0:0] v_7469;
  wire [0:0] v_7470;
  wire [0:0] v_7471;
  function [0:0] mux_7471(input [0:0] sel);
    case (sel) 0: mux_7471 = 1'h0; 1: mux_7471 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7472;
  function [0:0] mux_7472(input [0:0] sel);
    case (sel) 0: mux_7472 = 1'h0; 1: mux_7472 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7473;
  wire [0:0] v_7474;
  wire [0:0] v_7475;
  wire [0:0] v_7476;
  function [0:0] mux_7476(input [0:0] sel);
    case (sel) 0: mux_7476 = 1'h0; 1: mux_7476 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7477;
  function [0:0] mux_7477(input [0:0] sel);
    case (sel) 0: mux_7477 = 1'h0; 1: mux_7477 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7478;
  wire [0:0] v_7479;
  wire [0:0] v_7480;
  wire [0:0] v_7481;
  wire [0:0] v_7482;
  wire [0:0] v_7483;
  function [0:0] mux_7483(input [0:0] sel);
    case (sel) 0: mux_7483 = 1'h0; 1: mux_7483 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7484;
  function [0:0] mux_7484(input [0:0] sel);
    case (sel) 0: mux_7484 = 1'h0; 1: mux_7484 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7485;
  wire [0:0] v_7486;
  wire [0:0] v_7487;
  wire [0:0] v_7488;
  function [0:0] mux_7488(input [0:0] sel);
    case (sel) 0: mux_7488 = 1'h0; 1: mux_7488 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7489;
  function [0:0] mux_7489(input [0:0] sel);
    case (sel) 0: mux_7489 = 1'h0; 1: mux_7489 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7490;
  wire [0:0] v_7491;
  wire [0:0] v_7492;
  wire [0:0] v_7493;
  wire [0:0] v_7494;
  wire [0:0] v_7495;
  function [0:0] mux_7495(input [0:0] sel);
    case (sel) 0: mux_7495 = 1'h0; 1: mux_7495 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7496;
  wire [0:0] v_7497;
  function [0:0] mux_7497(input [0:0] sel);
    case (sel) 0: mux_7497 = 1'h0; 1: mux_7497 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7498;
  wire [0:0] v_7499;
  wire [0:0] v_7500;
  wire [0:0] v_7501;
  function [0:0] mux_7501(input [0:0] sel);
    case (sel) 0: mux_7501 = 1'h0; 1: mux_7501 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7502;
  function [0:0] mux_7502(input [0:0] sel);
    case (sel) 0: mux_7502 = 1'h0; 1: mux_7502 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7503 = 1'h0;
  wire [0:0] v_7504;
  wire [0:0] v_7505;
  wire [0:0] act_7506;
  wire [0:0] v_7507;
  wire [0:0] v_7508;
  wire [0:0] v_7509;
  reg [0:0] v_7510 = 1'h0;
  wire [0:0] v_7511;
  wire [0:0] v_7512;
  wire [0:0] act_7513;
  wire [0:0] v_7514;
  wire [0:0] v_7515;
  wire [0:0] v_7516;
  reg [0:0] v_7517 = 1'h0;
  wire [0:0] v_7518;
  wire [0:0] v_7519;
  wire [0:0] act_7520;
  wire [0:0] v_7521;
  wire [0:0] v_7522;
  wire [0:0] v_7523;
  wire [0:0] v_7524;
  wire [0:0] v_7525;
  wire [0:0] v_7526;
  function [0:0] mux_7526(input [0:0] sel);
    case (sel) 0: mux_7526 = 1'h0; 1: mux_7526 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7527;
  wire [0:0] v_7528;
  function [0:0] mux_7528(input [0:0] sel);
    case (sel) 0: mux_7528 = 1'h0; 1: mux_7528 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7529;
  wire [0:0] v_7530;
  wire [0:0] v_7531;
  wire [0:0] v_7532;
  function [0:0] mux_7532(input [0:0] sel);
    case (sel) 0: mux_7532 = 1'h0; 1: mux_7532 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7533;
  function [0:0] mux_7533(input [0:0] sel);
    case (sel) 0: mux_7533 = 1'h0; 1: mux_7533 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7534 = 1'h0;
  wire [0:0] v_7535;
  wire [0:0] v_7536;
  wire [0:0] act_7537;
  wire [0:0] v_7538;
  wire [0:0] v_7539;
  wire [0:0] v_7540;
  wire [0:0] v_7541;
  wire [0:0] v_7542;
  wire [0:0] v_7543;
  function [0:0] mux_7543(input [0:0] sel);
    case (sel) 0: mux_7543 = 1'h0; 1: mux_7543 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7544;
  function [0:0] mux_7544(input [0:0] sel);
    case (sel) 0: mux_7544 = 1'h0; 1: mux_7544 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7545;
  wire [0:0] v_7546;
  wire [0:0] v_7547;
  wire [0:0] v_7548;
  function [0:0] mux_7548(input [0:0] sel);
    case (sel) 0: mux_7548 = 1'h0; 1: mux_7548 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7549;
  function [0:0] mux_7549(input [0:0] sel);
    case (sel) 0: mux_7549 = 1'h0; 1: mux_7549 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7550;
  wire [0:0] v_7551;
  wire [0:0] v_7552;
  wire [0:0] v_7553;
  wire [0:0] v_7554;
  wire [0:0] v_7555;
  function [0:0] mux_7555(input [0:0] sel);
    case (sel) 0: mux_7555 = 1'h0; 1: mux_7555 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7556;
  wire [0:0] v_7557;
  function [0:0] mux_7557(input [0:0] sel);
    case (sel) 0: mux_7557 = 1'h0; 1: mux_7557 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7558;
  wire [0:0] v_7559;
  wire [0:0] v_7560;
  wire [0:0] v_7561;
  function [0:0] mux_7561(input [0:0] sel);
    case (sel) 0: mux_7561 = 1'h0; 1: mux_7561 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7562;
  function [0:0] mux_7562(input [0:0] sel);
    case (sel) 0: mux_7562 = 1'h0; 1: mux_7562 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7563 = 1'h0;
  wire [0:0] v_7564;
  wire [0:0] v_7565;
  wire [0:0] act_7566;
  wire [0:0] v_7567;
  wire [0:0] v_7568;
  wire [0:0] v_7569;
  reg [0:0] v_7570 = 1'h0;
  wire [0:0] v_7571;
  wire [0:0] v_7572;
  wire [0:0] act_7573;
  wire [0:0] v_7574;
  wire [0:0] v_7575;
  wire [0:0] v_7576;
  wire [0:0] v_7577;
  wire [0:0] v_7578;
  wire [0:0] v_7579;
  function [0:0] mux_7579(input [0:0] sel);
    case (sel) 0: mux_7579 = 1'h0; 1: mux_7579 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7580;
  wire [0:0] v_7581;
  function [0:0] mux_7581(input [0:0] sel);
    case (sel) 0: mux_7581 = 1'h0; 1: mux_7581 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7582;
  wire [0:0] v_7583;
  wire [0:0] v_7584;
  wire [0:0] v_7585;
  function [0:0] mux_7585(input [0:0] sel);
    case (sel) 0: mux_7585 = 1'h0; 1: mux_7585 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7586;
  function [0:0] mux_7586(input [0:0] sel);
    case (sel) 0: mux_7586 = 1'h0; 1: mux_7586 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7587 = 1'h0;
  wire [0:0] v_7588;
  wire [0:0] v_7589;
  wire [0:0] act_7590;
  wire [0:0] v_7591;
  wire [0:0] v_7592;
  wire [0:0] v_7593;
  wire [0:0] v_7594;
  wire [0:0] v_7595;
  wire [0:0] v_7596;
  function [0:0] mux_7596(input [0:0] sel);
    case (sel) 0: mux_7596 = 1'h0; 1: mux_7596 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7597;
  function [0:0] mux_7597(input [0:0] sel);
    case (sel) 0: mux_7597 = 1'h0; 1: mux_7597 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7598;
  wire [0:0] v_7599;
  wire [0:0] v_7600;
  wire [0:0] v_7601;
  function [0:0] mux_7601(input [0:0] sel);
    case (sel) 0: mux_7601 = 1'h0; 1: mux_7601 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7602;
  function [0:0] mux_7602(input [0:0] sel);
    case (sel) 0: mux_7602 = 1'h0; 1: mux_7602 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7603;
  wire [0:0] v_7604;
  wire [0:0] v_7605;
  wire [0:0] v_7606;
  wire [0:0] v_7607;
  wire [0:0] v_7608;
  function [0:0] mux_7608(input [0:0] sel);
    case (sel) 0: mux_7608 = 1'h0; 1: mux_7608 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7609;
  function [0:0] mux_7609(input [0:0] sel);
    case (sel) 0: mux_7609 = 1'h0; 1: mux_7609 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7610;
  wire [0:0] v_7611;
  wire [0:0] v_7612;
  wire [0:0] v_7613;
  function [0:0] mux_7613(input [0:0] sel);
    case (sel) 0: mux_7613 = 1'h0; 1: mux_7613 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7614;
  function [0:0] mux_7614(input [0:0] sel);
    case (sel) 0: mux_7614 = 1'h0; 1: mux_7614 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7615;
  wire [0:0] v_7616;
  wire [0:0] v_7617;
  wire [0:0] v_7618;
  wire [0:0] v_7619;
  wire [0:0] v_7620;
  function [0:0] mux_7620(input [0:0] sel);
    case (sel) 0: mux_7620 = 1'h0; 1: mux_7620 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7621;
  function [0:0] mux_7621(input [0:0] sel);
    case (sel) 0: mux_7621 = 1'h0; 1: mux_7621 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7622;
  wire [0:0] v_7623;
  wire [0:0] v_7624;
  wire [0:0] v_7625;
  function [0:0] mux_7625(input [0:0] sel);
    case (sel) 0: mux_7625 = 1'h0; 1: mux_7625 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7626;
  function [0:0] mux_7626(input [0:0] sel);
    case (sel) 0: mux_7626 = 1'h0; 1: mux_7626 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7627;
  wire [0:0] v_7628;
  wire [0:0] v_7629;
  wire [0:0] v_7630;
  wire [0:0] v_7631;
  wire [0:0] v_7632;
  function [0:0] mux_7632(input [0:0] sel);
    case (sel) 0: mux_7632 = 1'h0; 1: mux_7632 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7633;
  function [0:0] mux_7633(input [0:0] sel);
    case (sel) 0: mux_7633 = 1'h0; 1: mux_7633 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7634;
  wire [0:0] v_7635;
  wire [0:0] v_7636;
  wire [0:0] v_7637;
  function [0:0] mux_7637(input [0:0] sel);
    case (sel) 0: mux_7637 = 1'h0; 1: mux_7637 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7638;
  function [0:0] mux_7638(input [0:0] sel);
    case (sel) 0: mux_7638 = 1'h0; 1: mux_7638 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7639;
  wire [0:0] v_7640;
  wire [0:0] v_7641;
  wire [0:0] v_7642;
  wire [0:0] v_7643;
  wire [0:0] v_7644;
  function [0:0] mux_7644(input [0:0] sel);
    case (sel) 0: mux_7644 = 1'h0; 1: mux_7644 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7645;
  function [0:0] mux_7645(input [0:0] sel);
    case (sel) 0: mux_7645 = 1'h0; 1: mux_7645 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7646;
  wire [0:0] v_7647;
  wire [0:0] v_7648;
  wire [0:0] v_7649;
  function [0:0] mux_7649(input [0:0] sel);
    case (sel) 0: mux_7649 = 1'h0; 1: mux_7649 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7650;
  function [0:0] mux_7650(input [0:0] sel);
    case (sel) 0: mux_7650 = 1'h0; 1: mux_7650 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7651;
  wire [0:0] v_7652;
  wire [0:0] v_7653;
  wire [0:0] v_7654;
  wire [0:0] v_7655;
  wire [0:0] v_7656;
  function [0:0] mux_7656(input [0:0] sel);
    case (sel) 0: mux_7656 = 1'h0; 1: mux_7656 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7657;
  function [0:0] mux_7657(input [0:0] sel);
    case (sel) 0: mux_7657 = 1'h0; 1: mux_7657 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7658;
  wire [0:0] v_7659;
  wire [0:0] v_7660;
  wire [0:0] v_7661;
  function [0:0] mux_7661(input [0:0] sel);
    case (sel) 0: mux_7661 = 1'h0; 1: mux_7661 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7662;
  function [0:0] mux_7662(input [0:0] sel);
    case (sel) 0: mux_7662 = 1'h0; 1: mux_7662 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7663;
  wire [0:0] v_7664;
  wire [0:0] v_7665;
  wire [0:0] v_7666;
  wire [0:0] v_7667;
  wire [0:0] v_7668;
  function [0:0] mux_7668(input [0:0] sel);
    case (sel) 0: mux_7668 = 1'h0; 1: mux_7668 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7669;
  wire [0:0] v_7670;
  function [0:0] mux_7670(input [0:0] sel);
    case (sel) 0: mux_7670 = 1'h0; 1: mux_7670 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7671;
  wire [0:0] v_7672;
  wire [0:0] v_7673;
  wire [0:0] v_7674;
  function [0:0] mux_7674(input [0:0] sel);
    case (sel) 0: mux_7674 = 1'h0; 1: mux_7674 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7675;
  function [0:0] mux_7675(input [0:0] sel);
    case (sel) 0: mux_7675 = 1'h0; 1: mux_7675 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7676 = 1'h0;
  wire [0:0] v_7677;
  wire [0:0] v_7678;
  wire [0:0] act_7679;
  wire [0:0] v_7680;
  wire [0:0] v_7681;
  wire [0:0] v_7682;
  reg [0:0] v_7683 = 1'h0;
  wire [0:0] v_7684;
  wire [0:0] v_7685;
  wire [0:0] act_7686;
  wire [0:0] v_7687;
  wire [0:0] v_7688;
  wire [0:0] v_7689;
  reg [0:0] v_7690 = 1'h0;
  wire [0:0] v_7691;
  wire [0:0] v_7692;
  wire [0:0] act_7693;
  wire [0:0] v_7694;
  wire [0:0] v_7695;
  wire [0:0] v_7696;
  reg [0:0] v_7697 = 1'h0;
  wire [0:0] v_7698;
  wire [0:0] v_7699;
  wire [0:0] act_7700;
  wire [0:0] v_7701;
  wire [0:0] v_7702;
  wire [0:0] v_7703;
  reg [0:0] v_7704 = 1'h0;
  wire [0:0] v_7705;
  wire [0:0] v_7706;
  wire [0:0] act_7707;
  wire [0:0] v_7708;
  wire [0:0] v_7709;
  wire [0:0] v_7710;
  reg [0:0] v_7711 = 1'h0;
  wire [0:0] v_7712;
  wire [0:0] v_7713;
  wire [0:0] act_7714;
  wire [0:0] v_7715;
  wire [0:0] v_7716;
  wire [0:0] v_7717;
  reg [0:0] v_7718 = 1'h0;
  wire [0:0] v_7719;
  wire [0:0] v_7720;
  wire [0:0] act_7721;
  wire [0:0] v_7722;
  wire [0:0] v_7723;
  wire [0:0] v_7724;
  wire [0:0] v_7725;
  wire [0:0] v_7726;
  wire [0:0] v_7727;
  function [0:0] mux_7727(input [0:0] sel);
    case (sel) 0: mux_7727 = 1'h0; 1: mux_7727 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7728;
  wire [0:0] v_7729;
  function [0:0] mux_7729(input [0:0] sel);
    case (sel) 0: mux_7729 = 1'h0; 1: mux_7729 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7730;
  wire [0:0] v_7731;
  wire [0:0] v_7732;
  wire [0:0] v_7733;
  function [0:0] mux_7733(input [0:0] sel);
    case (sel) 0: mux_7733 = 1'h0; 1: mux_7733 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7734;
  function [0:0] mux_7734(input [0:0] sel);
    case (sel) 0: mux_7734 = 1'h0; 1: mux_7734 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7735 = 1'h0;
  wire [0:0] v_7736;
  wire [0:0] v_7737;
  wire [0:0] act_7738;
  wire [0:0] v_7739;
  wire [0:0] v_7740;
  wire [0:0] v_7741;
  wire [0:0] v_7742;
  wire [0:0] v_7743;
  wire [0:0] v_7744;
  function [0:0] mux_7744(input [0:0] sel);
    case (sel) 0: mux_7744 = 1'h0; 1: mux_7744 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7745;
  function [0:0] mux_7745(input [0:0] sel);
    case (sel) 0: mux_7745 = 1'h0; 1: mux_7745 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7746;
  wire [0:0] v_7747;
  wire [0:0] v_7748;
  wire [0:0] v_7749;
  function [0:0] mux_7749(input [0:0] sel);
    case (sel) 0: mux_7749 = 1'h0; 1: mux_7749 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7750;
  function [0:0] mux_7750(input [0:0] sel);
    case (sel) 0: mux_7750 = 1'h0; 1: mux_7750 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7751;
  wire [0:0] v_7752;
  wire [0:0] v_7753;
  wire [0:0] v_7754;
  wire [0:0] v_7755;
  wire [0:0] v_7756;
  function [0:0] mux_7756(input [0:0] sel);
    case (sel) 0: mux_7756 = 1'h0; 1: mux_7756 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7757;
  wire [0:0] v_7758;
  function [0:0] mux_7758(input [0:0] sel);
    case (sel) 0: mux_7758 = 1'h0; 1: mux_7758 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7759;
  wire [0:0] v_7760;
  wire [0:0] v_7761;
  wire [0:0] v_7762;
  function [0:0] mux_7762(input [0:0] sel);
    case (sel) 0: mux_7762 = 1'h0; 1: mux_7762 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7763;
  function [0:0] mux_7763(input [0:0] sel);
    case (sel) 0: mux_7763 = 1'h0; 1: mux_7763 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7764 = 1'h0;
  wire [0:0] v_7765;
  wire [0:0] v_7766;
  wire [0:0] act_7767;
  wire [0:0] v_7768;
  wire [0:0] v_7769;
  wire [0:0] v_7770;
  reg [0:0] v_7771 = 1'h0;
  wire [0:0] v_7772;
  wire [0:0] v_7773;
  wire [0:0] act_7774;
  wire [0:0] v_7775;
  wire [0:0] v_7776;
  wire [0:0] v_7777;
  wire [0:0] v_7778;
  wire [0:0] v_7779;
  wire [0:0] v_7780;
  function [0:0] mux_7780(input [0:0] sel);
    case (sel) 0: mux_7780 = 1'h0; 1: mux_7780 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7781;
  wire [0:0] v_7782;
  function [0:0] mux_7782(input [0:0] sel);
    case (sel) 0: mux_7782 = 1'h0; 1: mux_7782 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7783;
  wire [0:0] v_7784;
  wire [0:0] v_7785;
  wire [0:0] v_7786;
  function [0:0] mux_7786(input [0:0] sel);
    case (sel) 0: mux_7786 = 1'h0; 1: mux_7786 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7787;
  function [0:0] mux_7787(input [0:0] sel);
    case (sel) 0: mux_7787 = 1'h0; 1: mux_7787 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7788 = 1'h0;
  wire [0:0] v_7789;
  wire [0:0] v_7790;
  wire [0:0] act_7791;
  wire [0:0] v_7792;
  wire [0:0] v_7793;
  wire [0:0] v_7794;
  wire [0:0] v_7795;
  wire [0:0] v_7796;
  wire [0:0] v_7797;
  function [0:0] mux_7797(input [0:0] sel);
    case (sel) 0: mux_7797 = 1'h0; 1: mux_7797 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7798;
  function [0:0] mux_7798(input [0:0] sel);
    case (sel) 0: mux_7798 = 1'h0; 1: mux_7798 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7799;
  wire [0:0] v_7800;
  wire [0:0] v_7801;
  wire [0:0] v_7802;
  function [0:0] mux_7802(input [0:0] sel);
    case (sel) 0: mux_7802 = 1'h0; 1: mux_7802 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7803;
  function [0:0] mux_7803(input [0:0] sel);
    case (sel) 0: mux_7803 = 1'h0; 1: mux_7803 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7804;
  wire [0:0] v_7805;
  wire [0:0] v_7806;
  wire [0:0] v_7807;
  wire [0:0] v_7808;
  wire [0:0] v_7809;
  function [0:0] mux_7809(input [0:0] sel);
    case (sel) 0: mux_7809 = 1'h0; 1: mux_7809 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7810;
  function [0:0] mux_7810(input [0:0] sel);
    case (sel) 0: mux_7810 = 1'h0; 1: mux_7810 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7811;
  wire [0:0] v_7812;
  wire [0:0] v_7813;
  wire [0:0] v_7814;
  function [0:0] mux_7814(input [0:0] sel);
    case (sel) 0: mux_7814 = 1'h0; 1: mux_7814 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7815;
  function [0:0] mux_7815(input [0:0] sel);
    case (sel) 0: mux_7815 = 1'h0; 1: mux_7815 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7816;
  wire [0:0] v_7817;
  wire [0:0] v_7818;
  wire [0:0] v_7819;
  wire [0:0] v_7820;
  wire [0:0] v_7821;
  function [0:0] mux_7821(input [0:0] sel);
    case (sel) 0: mux_7821 = 1'h0; 1: mux_7821 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7822;
  wire [0:0] v_7823;
  function [0:0] mux_7823(input [0:0] sel);
    case (sel) 0: mux_7823 = 1'h0; 1: mux_7823 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7824;
  wire [0:0] v_7825;
  wire [0:0] v_7826;
  wire [0:0] v_7827;
  function [0:0] mux_7827(input [0:0] sel);
    case (sel) 0: mux_7827 = 1'h0; 1: mux_7827 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7828;
  function [0:0] mux_7828(input [0:0] sel);
    case (sel) 0: mux_7828 = 1'h0; 1: mux_7828 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7829 = 1'h0;
  wire [0:0] v_7830;
  wire [0:0] v_7831;
  wire [0:0] act_7832;
  wire [0:0] v_7833;
  wire [0:0] v_7834;
  wire [0:0] v_7835;
  reg [0:0] v_7836 = 1'h0;
  wire [0:0] v_7837;
  wire [0:0] v_7838;
  wire [0:0] act_7839;
  wire [0:0] v_7840;
  wire [0:0] v_7841;
  wire [0:0] v_7842;
  reg [0:0] v_7843 = 1'h0;
  wire [0:0] v_7844;
  wire [0:0] v_7845;
  wire [0:0] act_7846;
  wire [0:0] v_7847;
  wire [0:0] v_7848;
  wire [0:0] v_7849;
  wire [0:0] v_7850;
  wire [0:0] v_7851;
  wire [0:0] v_7852;
  function [0:0] mux_7852(input [0:0] sel);
    case (sel) 0: mux_7852 = 1'h0; 1: mux_7852 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7853;
  wire [0:0] v_7854;
  function [0:0] mux_7854(input [0:0] sel);
    case (sel) 0: mux_7854 = 1'h0; 1: mux_7854 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7855;
  wire [0:0] v_7856;
  wire [0:0] v_7857;
  wire [0:0] v_7858;
  function [0:0] mux_7858(input [0:0] sel);
    case (sel) 0: mux_7858 = 1'h0; 1: mux_7858 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7859;
  function [0:0] mux_7859(input [0:0] sel);
    case (sel) 0: mux_7859 = 1'h0; 1: mux_7859 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7860 = 1'h0;
  wire [0:0] v_7861;
  wire [0:0] v_7862;
  wire [0:0] act_7863;
  wire [0:0] v_7864;
  wire [0:0] v_7865;
  wire [0:0] v_7866;
  wire [0:0] v_7867;
  wire [0:0] v_7868;
  wire [0:0] v_7869;
  function [0:0] mux_7869(input [0:0] sel);
    case (sel) 0: mux_7869 = 1'h0; 1: mux_7869 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7870;
  function [0:0] mux_7870(input [0:0] sel);
    case (sel) 0: mux_7870 = 1'h0; 1: mux_7870 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7871;
  wire [0:0] v_7872;
  wire [0:0] v_7873;
  wire [0:0] v_7874;
  function [0:0] mux_7874(input [0:0] sel);
    case (sel) 0: mux_7874 = 1'h0; 1: mux_7874 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7875;
  function [0:0] mux_7875(input [0:0] sel);
    case (sel) 0: mux_7875 = 1'h0; 1: mux_7875 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7876;
  wire [0:0] v_7877;
  wire [0:0] v_7878;
  wire [0:0] v_7879;
  wire [0:0] v_7880;
  wire [0:0] v_7881;
  function [0:0] mux_7881(input [0:0] sel);
    case (sel) 0: mux_7881 = 1'h0; 1: mux_7881 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7882;
  wire [0:0] v_7883;
  function [0:0] mux_7883(input [0:0] sel);
    case (sel) 0: mux_7883 = 1'h0; 1: mux_7883 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7884;
  wire [0:0] v_7885;
  wire [0:0] v_7886;
  wire [0:0] v_7887;
  function [0:0] mux_7887(input [0:0] sel);
    case (sel) 0: mux_7887 = 1'h0; 1: mux_7887 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7888;
  function [0:0] mux_7888(input [0:0] sel);
    case (sel) 0: mux_7888 = 1'h0; 1: mux_7888 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7889 = 1'h0;
  wire [0:0] v_7890;
  wire [0:0] v_7891;
  wire [0:0] act_7892;
  wire [0:0] v_7893;
  wire [0:0] v_7894;
  wire [0:0] v_7895;
  reg [0:0] v_7896 = 1'h0;
  wire [0:0] v_7897;
  wire [0:0] v_7898;
  wire [0:0] act_7899;
  wire [0:0] v_7900;
  wire [0:0] v_7901;
  wire [0:0] v_7902;
  wire [0:0] v_7903;
  wire [0:0] v_7904;
  wire [0:0] v_7905;
  function [0:0] mux_7905(input [0:0] sel);
    case (sel) 0: mux_7905 = 1'h0; 1: mux_7905 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7906;
  wire [0:0] v_7907;
  function [0:0] mux_7907(input [0:0] sel);
    case (sel) 0: mux_7907 = 1'h0; 1: mux_7907 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7908;
  wire [0:0] v_7909;
  wire [0:0] v_7910;
  wire [0:0] v_7911;
  function [0:0] mux_7911(input [0:0] sel);
    case (sel) 0: mux_7911 = 1'h0; 1: mux_7911 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7912;
  function [0:0] mux_7912(input [0:0] sel);
    case (sel) 0: mux_7912 = 1'h0; 1: mux_7912 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7913 = 1'h0;
  wire [0:0] v_7914;
  wire [0:0] v_7915;
  wire [0:0] act_7916;
  wire [0:0] v_7917;
  wire [0:0] v_7918;
  wire [0:0] v_7919;
  wire [0:0] v_7920;
  wire [0:0] v_7921;
  wire [0:0] v_7922;
  function [0:0] mux_7922(input [0:0] sel);
    case (sel) 0: mux_7922 = 1'h0; 1: mux_7922 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7923;
  function [0:0] mux_7923(input [0:0] sel);
    case (sel) 0: mux_7923 = 1'h0; 1: mux_7923 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7924;
  wire [0:0] v_7925;
  wire [0:0] v_7926;
  wire [0:0] v_7927;
  function [0:0] mux_7927(input [0:0] sel);
    case (sel) 0: mux_7927 = 1'h0; 1: mux_7927 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7928;
  function [0:0] mux_7928(input [0:0] sel);
    case (sel) 0: mux_7928 = 1'h0; 1: mux_7928 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7929;
  wire [0:0] v_7930;
  wire [0:0] v_7931;
  wire [0:0] v_7932;
  wire [0:0] v_7933;
  wire [0:0] v_7934;
  function [0:0] mux_7934(input [0:0] sel);
    case (sel) 0: mux_7934 = 1'h0; 1: mux_7934 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7935;
  function [0:0] mux_7935(input [0:0] sel);
    case (sel) 0: mux_7935 = 1'h0; 1: mux_7935 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7936;
  wire [0:0] v_7937;
  wire [0:0] v_7938;
  wire [0:0] v_7939;
  function [0:0] mux_7939(input [0:0] sel);
    case (sel) 0: mux_7939 = 1'h0; 1: mux_7939 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7940;
  function [0:0] mux_7940(input [0:0] sel);
    case (sel) 0: mux_7940 = 1'h0; 1: mux_7940 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7941;
  wire [0:0] v_7942;
  wire [0:0] v_7943;
  wire [0:0] v_7944;
  wire [0:0] v_7945;
  wire [0:0] v_7946;
  function [0:0] mux_7946(input [0:0] sel);
    case (sel) 0: mux_7946 = 1'h0; 1: mux_7946 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7947;
  function [0:0] mux_7947(input [0:0] sel);
    case (sel) 0: mux_7947 = 1'h0; 1: mux_7947 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7948;
  wire [0:0] v_7949;
  wire [0:0] v_7950;
  wire [0:0] v_7951;
  function [0:0] mux_7951(input [0:0] sel);
    case (sel) 0: mux_7951 = 1'h0; 1: mux_7951 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7952;
  function [0:0] mux_7952(input [0:0] sel);
    case (sel) 0: mux_7952 = 1'h0; 1: mux_7952 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7953;
  wire [0:0] v_7954;
  wire [0:0] v_7955;
  wire [0:0] v_7956;
  wire [0:0] v_7957;
  wire [0:0] v_7958;
  function [0:0] mux_7958(input [0:0] sel);
    case (sel) 0: mux_7958 = 1'h0; 1: mux_7958 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7959;
  wire [0:0] v_7960;
  function [0:0] mux_7960(input [0:0] sel);
    case (sel) 0: mux_7960 = 1'h0; 1: mux_7960 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7961;
  wire [0:0] v_7962;
  wire [0:0] v_7963;
  wire [0:0] v_7964;
  function [0:0] mux_7964(input [0:0] sel);
    case (sel) 0: mux_7964 = 1'h0; 1: mux_7964 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7965;
  function [0:0] mux_7965(input [0:0] sel);
    case (sel) 0: mux_7965 = 1'h0; 1: mux_7965 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_7966 = 1'h0;
  wire [0:0] v_7967;
  wire [0:0] v_7968;
  wire [0:0] act_7969;
  wire [0:0] v_7970;
  wire [0:0] v_7971;
  wire [0:0] v_7972;
  reg [0:0] v_7973 = 1'h0;
  wire [0:0] v_7974;
  wire [0:0] v_7975;
  wire [0:0] act_7976;
  wire [0:0] v_7977;
  wire [0:0] v_7978;
  wire [0:0] v_7979;
  reg [0:0] v_7980 = 1'h0;
  wire [0:0] v_7981;
  wire [0:0] v_7982;
  wire [0:0] act_7983;
  wire [0:0] v_7984;
  wire [0:0] v_7985;
  wire [0:0] v_7986;
  reg [0:0] v_7987 = 1'h0;
  wire [0:0] v_7988;
  wire [0:0] v_7989;
  wire [0:0] act_7990;
  wire [0:0] v_7991;
  wire [0:0] v_7992;
  wire [0:0] v_7993;
  wire [0:0] v_7994;
  wire [0:0] v_7995;
  wire [0:0] v_7996;
  function [0:0] mux_7996(input [0:0] sel);
    case (sel) 0: mux_7996 = 1'h0; 1: mux_7996 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_7997;
  wire [0:0] v_7998;
  function [0:0] mux_7998(input [0:0] sel);
    case (sel) 0: mux_7998 = 1'h0; 1: mux_7998 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_7999;
  wire [0:0] v_8000;
  wire [0:0] v_8001;
  wire [0:0] v_8002;
  function [0:0] mux_8002(input [0:0] sel);
    case (sel) 0: mux_8002 = 1'h0; 1: mux_8002 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8003;
  function [0:0] mux_8003(input [0:0] sel);
    case (sel) 0: mux_8003 = 1'h0; 1: mux_8003 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8004 = 1'h0;
  wire [0:0] v_8005;
  wire [0:0] v_8006;
  wire [0:0] act_8007;
  wire [0:0] v_8008;
  wire [0:0] v_8009;
  wire [0:0] v_8010;
  wire [0:0] v_8011;
  wire [0:0] v_8012;
  wire [0:0] v_8013;
  function [0:0] mux_8013(input [0:0] sel);
    case (sel) 0: mux_8013 = 1'h0; 1: mux_8013 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8014;
  function [0:0] mux_8014(input [0:0] sel);
    case (sel) 0: mux_8014 = 1'h0; 1: mux_8014 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8015;
  wire [0:0] v_8016;
  wire [0:0] v_8017;
  wire [0:0] v_8018;
  function [0:0] mux_8018(input [0:0] sel);
    case (sel) 0: mux_8018 = 1'h0; 1: mux_8018 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8019;
  function [0:0] mux_8019(input [0:0] sel);
    case (sel) 0: mux_8019 = 1'h0; 1: mux_8019 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8020;
  wire [0:0] v_8021;
  wire [0:0] v_8022;
  wire [0:0] v_8023;
  wire [0:0] v_8024;
  wire [0:0] v_8025;
  function [0:0] mux_8025(input [0:0] sel);
    case (sel) 0: mux_8025 = 1'h0; 1: mux_8025 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8026;
  wire [0:0] v_8027;
  function [0:0] mux_8027(input [0:0] sel);
    case (sel) 0: mux_8027 = 1'h0; 1: mux_8027 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8028;
  wire [0:0] v_8029;
  wire [0:0] v_8030;
  wire [0:0] v_8031;
  function [0:0] mux_8031(input [0:0] sel);
    case (sel) 0: mux_8031 = 1'h0; 1: mux_8031 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8032;
  function [0:0] mux_8032(input [0:0] sel);
    case (sel) 0: mux_8032 = 1'h0; 1: mux_8032 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8033 = 1'h0;
  wire [0:0] v_8034;
  wire [0:0] v_8035;
  wire [0:0] act_8036;
  wire [0:0] v_8037;
  wire [0:0] v_8038;
  wire [0:0] v_8039;
  reg [0:0] v_8040 = 1'h0;
  wire [0:0] v_8041;
  wire [0:0] v_8042;
  wire [0:0] act_8043;
  wire [0:0] v_8044;
  wire [0:0] v_8045;
  wire [0:0] v_8046;
  wire [0:0] v_8047;
  wire [0:0] v_8048;
  wire [0:0] v_8049;
  function [0:0] mux_8049(input [0:0] sel);
    case (sel) 0: mux_8049 = 1'h0; 1: mux_8049 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8050;
  wire [0:0] v_8051;
  function [0:0] mux_8051(input [0:0] sel);
    case (sel) 0: mux_8051 = 1'h0; 1: mux_8051 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8052;
  wire [0:0] v_8053;
  wire [0:0] v_8054;
  wire [0:0] v_8055;
  function [0:0] mux_8055(input [0:0] sel);
    case (sel) 0: mux_8055 = 1'h0; 1: mux_8055 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8056;
  function [0:0] mux_8056(input [0:0] sel);
    case (sel) 0: mux_8056 = 1'h0; 1: mux_8056 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8057 = 1'h0;
  wire [0:0] v_8058;
  wire [0:0] v_8059;
  wire [0:0] act_8060;
  wire [0:0] v_8061;
  wire [0:0] v_8062;
  wire [0:0] v_8063;
  wire [0:0] v_8064;
  wire [0:0] v_8065;
  wire [0:0] v_8066;
  function [0:0] mux_8066(input [0:0] sel);
    case (sel) 0: mux_8066 = 1'h0; 1: mux_8066 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8067;
  function [0:0] mux_8067(input [0:0] sel);
    case (sel) 0: mux_8067 = 1'h0; 1: mux_8067 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8068;
  wire [0:0] v_8069;
  wire [0:0] v_8070;
  wire [0:0] v_8071;
  function [0:0] mux_8071(input [0:0] sel);
    case (sel) 0: mux_8071 = 1'h0; 1: mux_8071 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8072;
  function [0:0] mux_8072(input [0:0] sel);
    case (sel) 0: mux_8072 = 1'h0; 1: mux_8072 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8073;
  wire [0:0] v_8074;
  wire [0:0] v_8075;
  wire [0:0] v_8076;
  wire [0:0] v_8077;
  wire [0:0] v_8078;
  function [0:0] mux_8078(input [0:0] sel);
    case (sel) 0: mux_8078 = 1'h0; 1: mux_8078 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8079;
  function [0:0] mux_8079(input [0:0] sel);
    case (sel) 0: mux_8079 = 1'h0; 1: mux_8079 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8080;
  wire [0:0] v_8081;
  wire [0:0] v_8082;
  wire [0:0] v_8083;
  function [0:0] mux_8083(input [0:0] sel);
    case (sel) 0: mux_8083 = 1'h0; 1: mux_8083 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8084;
  function [0:0] mux_8084(input [0:0] sel);
    case (sel) 0: mux_8084 = 1'h0; 1: mux_8084 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8085;
  wire [0:0] v_8086;
  wire [0:0] v_8087;
  wire [0:0] v_8088;
  wire [0:0] v_8089;
  wire [0:0] v_8090;
  function [0:0] mux_8090(input [0:0] sel);
    case (sel) 0: mux_8090 = 1'h0; 1: mux_8090 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8091;
  wire [0:0] v_8092;
  function [0:0] mux_8092(input [0:0] sel);
    case (sel) 0: mux_8092 = 1'h0; 1: mux_8092 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8093;
  wire [0:0] v_8094;
  wire [0:0] v_8095;
  wire [0:0] v_8096;
  function [0:0] mux_8096(input [0:0] sel);
    case (sel) 0: mux_8096 = 1'h0; 1: mux_8096 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8097;
  function [0:0] mux_8097(input [0:0] sel);
    case (sel) 0: mux_8097 = 1'h0; 1: mux_8097 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8098 = 1'h0;
  wire [0:0] v_8099;
  wire [0:0] v_8100;
  wire [0:0] act_8101;
  wire [0:0] v_8102;
  wire [0:0] v_8103;
  wire [0:0] v_8104;
  reg [0:0] v_8105 = 1'h0;
  wire [0:0] v_8106;
  wire [0:0] v_8107;
  wire [0:0] act_8108;
  wire [0:0] v_8109;
  wire [0:0] v_8110;
  wire [0:0] v_8111;
  reg [0:0] v_8112 = 1'h0;
  wire [0:0] v_8113;
  wire [0:0] v_8114;
  wire [0:0] act_8115;
  wire [0:0] v_8116;
  wire [0:0] v_8117;
  wire [0:0] v_8118;
  wire [0:0] v_8119;
  wire [0:0] v_8120;
  wire [0:0] v_8121;
  function [0:0] mux_8121(input [0:0] sel);
    case (sel) 0: mux_8121 = 1'h0; 1: mux_8121 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8122;
  wire [0:0] v_8123;
  function [0:0] mux_8123(input [0:0] sel);
    case (sel) 0: mux_8123 = 1'h0; 1: mux_8123 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8124;
  wire [0:0] v_8125;
  wire [0:0] v_8126;
  wire [0:0] v_8127;
  function [0:0] mux_8127(input [0:0] sel);
    case (sel) 0: mux_8127 = 1'h0; 1: mux_8127 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8128;
  function [0:0] mux_8128(input [0:0] sel);
    case (sel) 0: mux_8128 = 1'h0; 1: mux_8128 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8129 = 1'h0;
  wire [0:0] v_8130;
  wire [0:0] v_8131;
  wire [0:0] act_8132;
  wire [0:0] v_8133;
  wire [0:0] v_8134;
  wire [0:0] v_8135;
  wire [0:0] v_8136;
  wire [0:0] v_8137;
  wire [0:0] v_8138;
  function [0:0] mux_8138(input [0:0] sel);
    case (sel) 0: mux_8138 = 1'h0; 1: mux_8138 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8139;
  function [0:0] mux_8139(input [0:0] sel);
    case (sel) 0: mux_8139 = 1'h0; 1: mux_8139 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8140;
  wire [0:0] v_8141;
  wire [0:0] v_8142;
  wire [0:0] v_8143;
  function [0:0] mux_8143(input [0:0] sel);
    case (sel) 0: mux_8143 = 1'h0; 1: mux_8143 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8144;
  function [0:0] mux_8144(input [0:0] sel);
    case (sel) 0: mux_8144 = 1'h0; 1: mux_8144 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8145;
  wire [0:0] v_8146;
  wire [0:0] v_8147;
  wire [0:0] v_8148;
  wire [0:0] v_8149;
  wire [0:0] v_8150;
  function [0:0] mux_8150(input [0:0] sel);
    case (sel) 0: mux_8150 = 1'h0; 1: mux_8150 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8151;
  wire [0:0] v_8152;
  function [0:0] mux_8152(input [0:0] sel);
    case (sel) 0: mux_8152 = 1'h0; 1: mux_8152 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8153;
  wire [0:0] v_8154;
  wire [0:0] v_8155;
  wire [0:0] v_8156;
  function [0:0] mux_8156(input [0:0] sel);
    case (sel) 0: mux_8156 = 1'h0; 1: mux_8156 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8157;
  function [0:0] mux_8157(input [0:0] sel);
    case (sel) 0: mux_8157 = 1'h0; 1: mux_8157 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8158 = 1'h0;
  wire [0:0] v_8159;
  wire [0:0] v_8160;
  wire [0:0] act_8161;
  wire [0:0] v_8162;
  wire [0:0] v_8163;
  wire [0:0] v_8164;
  reg [0:0] v_8165 = 1'h0;
  wire [0:0] v_8166;
  wire [0:0] v_8167;
  wire [0:0] act_8168;
  wire [0:0] v_8169;
  wire [0:0] v_8170;
  wire [0:0] v_8171;
  wire [0:0] v_8172;
  wire [0:0] v_8173;
  wire [0:0] v_8174;
  function [0:0] mux_8174(input [0:0] sel);
    case (sel) 0: mux_8174 = 1'h0; 1: mux_8174 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8175;
  wire [0:0] v_8176;
  function [0:0] mux_8176(input [0:0] sel);
    case (sel) 0: mux_8176 = 1'h0; 1: mux_8176 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8177;
  wire [0:0] v_8178;
  wire [0:0] v_8179;
  wire [0:0] v_8180;
  function [0:0] mux_8180(input [0:0] sel);
    case (sel) 0: mux_8180 = 1'h0; 1: mux_8180 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8181;
  function [0:0] mux_8181(input [0:0] sel);
    case (sel) 0: mux_8181 = 1'h0; 1: mux_8181 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8182 = 1'h0;
  wire [0:0] v_8183;
  wire [0:0] v_8184;
  wire [0:0] act_8185;
  wire [0:0] v_8186;
  wire [0:0] v_8187;
  wire [0:0] v_8188;
  wire [0:0] v_8189;
  wire [0:0] v_8190;
  wire [0:0] v_8191;
  function [0:0] mux_8191(input [0:0] sel);
    case (sel) 0: mux_8191 = 1'h0; 1: mux_8191 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8192;
  function [0:0] mux_8192(input [0:0] sel);
    case (sel) 0: mux_8192 = 1'h0; 1: mux_8192 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8193;
  wire [0:0] v_8194;
  wire [0:0] v_8195;
  wire [0:0] v_8196;
  function [0:0] mux_8196(input [0:0] sel);
    case (sel) 0: mux_8196 = 1'h0; 1: mux_8196 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8197;
  function [0:0] mux_8197(input [0:0] sel);
    case (sel) 0: mux_8197 = 1'h0; 1: mux_8197 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8198;
  wire [0:0] v_8199;
  wire [0:0] v_8200;
  wire [0:0] v_8201;
  wire [0:0] v_8202;
  wire [0:0] v_8203;
  function [0:0] mux_8203(input [0:0] sel);
    case (sel) 0: mux_8203 = 1'h0; 1: mux_8203 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8204;
  function [0:0] mux_8204(input [0:0] sel);
    case (sel) 0: mux_8204 = 1'h0; 1: mux_8204 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8205;
  wire [0:0] v_8206;
  wire [0:0] v_8207;
  wire [0:0] v_8208;
  function [0:0] mux_8208(input [0:0] sel);
    case (sel) 0: mux_8208 = 1'h0; 1: mux_8208 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8209;
  function [0:0] mux_8209(input [0:0] sel);
    case (sel) 0: mux_8209 = 1'h0; 1: mux_8209 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8210;
  wire [0:0] v_8211;
  wire [0:0] v_8212;
  wire [0:0] v_8213;
  wire [0:0] v_8214;
  wire [0:0] v_8215;
  function [0:0] mux_8215(input [0:0] sel);
    case (sel) 0: mux_8215 = 1'h0; 1: mux_8215 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8216;
  function [0:0] mux_8216(input [0:0] sel);
    case (sel) 0: mux_8216 = 1'h0; 1: mux_8216 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8217;
  wire [0:0] v_8218;
  wire [0:0] v_8219;
  wire [0:0] v_8220;
  function [0:0] mux_8220(input [0:0] sel);
    case (sel) 0: mux_8220 = 1'h0; 1: mux_8220 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8221;
  function [0:0] mux_8221(input [0:0] sel);
    case (sel) 0: mux_8221 = 1'h0; 1: mux_8221 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8222;
  wire [0:0] v_8223;
  wire [0:0] v_8224;
  wire [0:0] v_8225;
  wire [0:0] v_8226;
  wire [0:0] v_8227;
  function [0:0] mux_8227(input [0:0] sel);
    case (sel) 0: mux_8227 = 1'h0; 1: mux_8227 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8228;
  function [0:0] mux_8228(input [0:0] sel);
    case (sel) 0: mux_8228 = 1'h0; 1: mux_8228 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8229;
  wire [0:0] v_8230;
  wire [0:0] v_8231;
  wire [0:0] v_8232;
  function [0:0] mux_8232(input [0:0] sel);
    case (sel) 0: mux_8232 = 1'h0; 1: mux_8232 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8233;
  function [0:0] mux_8233(input [0:0] sel);
    case (sel) 0: mux_8233 = 1'h0; 1: mux_8233 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8234;
  wire [0:0] v_8235;
  wire [0:0] v_8236;
  wire [0:0] v_8237;
  wire [0:0] v_8238;
  wire [0:0] v_8239;
  function [0:0] mux_8239(input [0:0] sel);
    case (sel) 0: mux_8239 = 1'h0; 1: mux_8239 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8240;
  wire [0:0] v_8241;
  function [0:0] mux_8241(input [0:0] sel);
    case (sel) 0: mux_8241 = 1'h0; 1: mux_8241 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8242;
  wire [0:0] v_8243;
  wire [0:0] v_8244;
  wire [0:0] v_8245;
  function [0:0] mux_8245(input [0:0] sel);
    case (sel) 0: mux_8245 = 1'h0; 1: mux_8245 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8246;
  function [0:0] mux_8246(input [0:0] sel);
    case (sel) 0: mux_8246 = 1'h0; 1: mux_8246 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8247 = 1'h0;
  wire [0:0] v_8248;
  wire [0:0] v_8249;
  wire [0:0] act_8250;
  wire [0:0] v_8251;
  wire [0:0] v_8252;
  wire [0:0] v_8253;
  reg [0:0] v_8254 = 1'h0;
  wire [0:0] v_8255;
  wire [0:0] v_8256;
  wire [0:0] act_8257;
  wire [0:0] v_8258;
  wire [0:0] v_8259;
  wire [0:0] v_8260;
  reg [0:0] v_8261 = 1'h0;
  wire [0:0] v_8262;
  wire [0:0] v_8263;
  wire [0:0] act_8264;
  wire [0:0] v_8265;
  wire [0:0] v_8266;
  wire [0:0] v_8267;
  reg [0:0] v_8268 = 1'h0;
  wire [0:0] v_8269;
  wire [0:0] v_8270;
  wire [0:0] act_8271;
  wire [0:0] v_8272;
  wire [0:0] v_8273;
  wire [0:0] v_8274;
  reg [0:0] v_8275 = 1'h0;
  wire [0:0] v_8276;
  wire [0:0] v_8277;
  wire [0:0] act_8278;
  wire [0:0] v_8279;
  wire [0:0] v_8280;
  wire [0:0] v_8281;
  wire [0:0] v_8282;
  wire [0:0] v_8283;
  wire [0:0] v_8284;
  function [0:0] mux_8284(input [0:0] sel);
    case (sel) 0: mux_8284 = 1'h0; 1: mux_8284 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8285;
  wire [0:0] v_8286;
  function [0:0] mux_8286(input [0:0] sel);
    case (sel) 0: mux_8286 = 1'h0; 1: mux_8286 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8287;
  wire [0:0] v_8288;
  wire [0:0] v_8289;
  wire [0:0] v_8290;
  function [0:0] mux_8290(input [0:0] sel);
    case (sel) 0: mux_8290 = 1'h0; 1: mux_8290 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8291;
  function [0:0] mux_8291(input [0:0] sel);
    case (sel) 0: mux_8291 = 1'h0; 1: mux_8291 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8292 = 1'h0;
  wire [0:0] v_8293;
  wire [0:0] v_8294;
  wire [0:0] act_8295;
  wire [0:0] v_8296;
  wire [0:0] v_8297;
  wire [0:0] v_8298;
  wire [0:0] v_8299;
  wire [0:0] v_8300;
  wire [0:0] v_8301;
  function [0:0] mux_8301(input [0:0] sel);
    case (sel) 0: mux_8301 = 1'h0; 1: mux_8301 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8302;
  function [0:0] mux_8302(input [0:0] sel);
    case (sel) 0: mux_8302 = 1'h0; 1: mux_8302 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8303;
  wire [0:0] v_8304;
  wire [0:0] v_8305;
  wire [0:0] v_8306;
  function [0:0] mux_8306(input [0:0] sel);
    case (sel) 0: mux_8306 = 1'h0; 1: mux_8306 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8307;
  function [0:0] mux_8307(input [0:0] sel);
    case (sel) 0: mux_8307 = 1'h0; 1: mux_8307 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8308;
  wire [0:0] v_8309;
  wire [0:0] v_8310;
  wire [0:0] v_8311;
  wire [0:0] v_8312;
  wire [0:0] v_8313;
  function [0:0] mux_8313(input [0:0] sel);
    case (sel) 0: mux_8313 = 1'h0; 1: mux_8313 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8314;
  wire [0:0] v_8315;
  function [0:0] mux_8315(input [0:0] sel);
    case (sel) 0: mux_8315 = 1'h0; 1: mux_8315 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8316;
  wire [0:0] v_8317;
  wire [0:0] v_8318;
  wire [0:0] v_8319;
  function [0:0] mux_8319(input [0:0] sel);
    case (sel) 0: mux_8319 = 1'h0; 1: mux_8319 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8320;
  function [0:0] mux_8320(input [0:0] sel);
    case (sel) 0: mux_8320 = 1'h0; 1: mux_8320 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8321 = 1'h0;
  wire [0:0] v_8322;
  wire [0:0] v_8323;
  wire [0:0] act_8324;
  wire [0:0] v_8325;
  wire [0:0] v_8326;
  wire [0:0] v_8327;
  reg [0:0] v_8328 = 1'h0;
  wire [0:0] v_8329;
  wire [0:0] v_8330;
  wire [0:0] act_8331;
  wire [0:0] v_8332;
  wire [0:0] v_8333;
  wire [0:0] v_8334;
  wire [0:0] v_8335;
  wire [0:0] v_8336;
  wire [0:0] v_8337;
  function [0:0] mux_8337(input [0:0] sel);
    case (sel) 0: mux_8337 = 1'h0; 1: mux_8337 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8338;
  wire [0:0] v_8339;
  function [0:0] mux_8339(input [0:0] sel);
    case (sel) 0: mux_8339 = 1'h0; 1: mux_8339 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8340;
  wire [0:0] v_8341;
  wire [0:0] v_8342;
  wire [0:0] v_8343;
  function [0:0] mux_8343(input [0:0] sel);
    case (sel) 0: mux_8343 = 1'h0; 1: mux_8343 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8344;
  function [0:0] mux_8344(input [0:0] sel);
    case (sel) 0: mux_8344 = 1'h0; 1: mux_8344 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8345 = 1'h0;
  wire [0:0] v_8346;
  wire [0:0] v_8347;
  wire [0:0] act_8348;
  wire [0:0] v_8349;
  wire [0:0] v_8350;
  wire [0:0] v_8351;
  wire [0:0] v_8352;
  wire [0:0] v_8353;
  wire [0:0] v_8354;
  function [0:0] mux_8354(input [0:0] sel);
    case (sel) 0: mux_8354 = 1'h0; 1: mux_8354 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8355;
  function [0:0] mux_8355(input [0:0] sel);
    case (sel) 0: mux_8355 = 1'h0; 1: mux_8355 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8356;
  wire [0:0] v_8357;
  wire [0:0] v_8358;
  wire [0:0] v_8359;
  function [0:0] mux_8359(input [0:0] sel);
    case (sel) 0: mux_8359 = 1'h0; 1: mux_8359 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8360;
  function [0:0] mux_8360(input [0:0] sel);
    case (sel) 0: mux_8360 = 1'h0; 1: mux_8360 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8361;
  wire [0:0] v_8362;
  wire [0:0] v_8363;
  wire [0:0] v_8364;
  wire [0:0] v_8365;
  wire [0:0] v_8366;
  function [0:0] mux_8366(input [0:0] sel);
    case (sel) 0: mux_8366 = 1'h0; 1: mux_8366 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8367;
  function [0:0] mux_8367(input [0:0] sel);
    case (sel) 0: mux_8367 = 1'h0; 1: mux_8367 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8368;
  wire [0:0] v_8369;
  wire [0:0] v_8370;
  wire [0:0] v_8371;
  function [0:0] mux_8371(input [0:0] sel);
    case (sel) 0: mux_8371 = 1'h0; 1: mux_8371 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8372;
  function [0:0] mux_8372(input [0:0] sel);
    case (sel) 0: mux_8372 = 1'h0; 1: mux_8372 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8373;
  wire [0:0] v_8374;
  wire [0:0] v_8375;
  wire [0:0] v_8376;
  wire [0:0] v_8377;
  wire [0:0] v_8378;
  function [0:0] mux_8378(input [0:0] sel);
    case (sel) 0: mux_8378 = 1'h0; 1: mux_8378 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8379;
  wire [0:0] v_8380;
  function [0:0] mux_8380(input [0:0] sel);
    case (sel) 0: mux_8380 = 1'h0; 1: mux_8380 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8381;
  wire [0:0] v_8382;
  wire [0:0] v_8383;
  wire [0:0] v_8384;
  function [0:0] mux_8384(input [0:0] sel);
    case (sel) 0: mux_8384 = 1'h0; 1: mux_8384 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8385;
  function [0:0] mux_8385(input [0:0] sel);
    case (sel) 0: mux_8385 = 1'h0; 1: mux_8385 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8386 = 1'h0;
  wire [0:0] v_8387;
  wire [0:0] v_8388;
  wire [0:0] act_8389;
  wire [0:0] v_8390;
  wire [0:0] v_8391;
  wire [0:0] v_8392;
  reg [0:0] v_8393 = 1'h0;
  wire [0:0] v_8394;
  wire [0:0] v_8395;
  wire [0:0] act_8396;
  wire [0:0] v_8397;
  wire [0:0] v_8398;
  wire [0:0] v_8399;
  reg [0:0] v_8400 = 1'h0;
  wire [0:0] v_8401;
  wire [0:0] v_8402;
  wire [0:0] act_8403;
  wire [0:0] v_8404;
  wire [0:0] v_8405;
  wire [0:0] v_8406;
  wire [0:0] v_8407;
  wire [0:0] v_8408;
  wire [0:0] v_8409;
  function [0:0] mux_8409(input [0:0] sel);
    case (sel) 0: mux_8409 = 1'h0; 1: mux_8409 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8410;
  wire [0:0] v_8411;
  function [0:0] mux_8411(input [0:0] sel);
    case (sel) 0: mux_8411 = 1'h0; 1: mux_8411 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8412;
  wire [0:0] v_8413;
  wire [0:0] v_8414;
  wire [0:0] v_8415;
  function [0:0] mux_8415(input [0:0] sel);
    case (sel) 0: mux_8415 = 1'h0; 1: mux_8415 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8416;
  function [0:0] mux_8416(input [0:0] sel);
    case (sel) 0: mux_8416 = 1'h0; 1: mux_8416 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8417 = 1'h0;
  wire [0:0] v_8418;
  wire [0:0] v_8419;
  wire [0:0] act_8420;
  wire [0:0] v_8421;
  wire [0:0] v_8422;
  wire [0:0] v_8423;
  wire [0:0] v_8424;
  wire [0:0] v_8425;
  wire [0:0] v_8426;
  function [0:0] mux_8426(input [0:0] sel);
    case (sel) 0: mux_8426 = 1'h0; 1: mux_8426 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8427;
  function [0:0] mux_8427(input [0:0] sel);
    case (sel) 0: mux_8427 = 1'h0; 1: mux_8427 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8428;
  wire [0:0] v_8429;
  wire [0:0] v_8430;
  wire [0:0] v_8431;
  function [0:0] mux_8431(input [0:0] sel);
    case (sel) 0: mux_8431 = 1'h0; 1: mux_8431 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8432;
  function [0:0] mux_8432(input [0:0] sel);
    case (sel) 0: mux_8432 = 1'h0; 1: mux_8432 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8433;
  wire [0:0] v_8434;
  wire [0:0] v_8435;
  wire [0:0] v_8436;
  wire [0:0] v_8437;
  wire [0:0] v_8438;
  function [0:0] mux_8438(input [0:0] sel);
    case (sel) 0: mux_8438 = 1'h0; 1: mux_8438 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8439;
  wire [0:0] v_8440;
  function [0:0] mux_8440(input [0:0] sel);
    case (sel) 0: mux_8440 = 1'h0; 1: mux_8440 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8441;
  wire [0:0] v_8442;
  wire [0:0] v_8443;
  wire [0:0] v_8444;
  function [0:0] mux_8444(input [0:0] sel);
    case (sel) 0: mux_8444 = 1'h0; 1: mux_8444 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8445;
  function [0:0] mux_8445(input [0:0] sel);
    case (sel) 0: mux_8445 = 1'h0; 1: mux_8445 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8446 = 1'h0;
  wire [0:0] v_8447;
  wire [0:0] v_8448;
  wire [0:0] act_8449;
  wire [0:0] v_8450;
  wire [0:0] v_8451;
  wire [0:0] v_8452;
  reg [0:0] v_8453 = 1'h0;
  wire [0:0] v_8454;
  wire [0:0] v_8455;
  wire [0:0] act_8456;
  wire [0:0] v_8457;
  wire [0:0] v_8458;
  wire [0:0] v_8459;
  wire [0:0] v_8460;
  wire [0:0] v_8461;
  wire [0:0] v_8462;
  function [0:0] mux_8462(input [0:0] sel);
    case (sel) 0: mux_8462 = 1'h0; 1: mux_8462 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8463;
  wire [0:0] v_8464;
  function [0:0] mux_8464(input [0:0] sel);
    case (sel) 0: mux_8464 = 1'h0; 1: mux_8464 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8465;
  wire [0:0] v_8466;
  wire [0:0] v_8467;
  wire [0:0] v_8468;
  function [0:0] mux_8468(input [0:0] sel);
    case (sel) 0: mux_8468 = 1'h0; 1: mux_8468 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8469;
  function [0:0] mux_8469(input [0:0] sel);
    case (sel) 0: mux_8469 = 1'h0; 1: mux_8469 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8470 = 1'h0;
  wire [0:0] v_8471;
  wire [0:0] v_8472;
  wire [0:0] act_8473;
  wire [0:0] v_8474;
  wire [0:0] v_8475;
  wire [0:0] v_8476;
  wire [0:0] v_8477;
  wire [0:0] v_8478;
  wire [0:0] v_8479;
  function [0:0] mux_8479(input [0:0] sel);
    case (sel) 0: mux_8479 = 1'h0; 1: mux_8479 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8480;
  function [0:0] mux_8480(input [0:0] sel);
    case (sel) 0: mux_8480 = 1'h0; 1: mux_8480 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8481;
  wire [0:0] v_8482;
  wire [0:0] v_8483;
  wire [0:0] v_8484;
  function [0:0] mux_8484(input [0:0] sel);
    case (sel) 0: mux_8484 = 1'h0; 1: mux_8484 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8485;
  function [0:0] mux_8485(input [0:0] sel);
    case (sel) 0: mux_8485 = 1'h0; 1: mux_8485 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8486;
  wire [0:0] v_8487;
  wire [0:0] v_8488;
  wire [0:0] v_8489;
  wire [0:0] v_8490;
  wire [0:0] v_8491;
  function [0:0] mux_8491(input [0:0] sel);
    case (sel) 0: mux_8491 = 1'h0; 1: mux_8491 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8492;
  function [0:0] mux_8492(input [0:0] sel);
    case (sel) 0: mux_8492 = 1'h0; 1: mux_8492 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8493;
  wire [0:0] v_8494;
  wire [0:0] v_8495;
  wire [0:0] v_8496;
  function [0:0] mux_8496(input [0:0] sel);
    case (sel) 0: mux_8496 = 1'h0; 1: mux_8496 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8497;
  function [0:0] mux_8497(input [0:0] sel);
    case (sel) 0: mux_8497 = 1'h0; 1: mux_8497 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8498;
  wire [0:0] v_8499;
  wire [0:0] v_8500;
  wire [0:0] v_8501;
  wire [0:0] v_8502;
  wire [0:0] v_8503;
  function [0:0] mux_8503(input [0:0] sel);
    case (sel) 0: mux_8503 = 1'h0; 1: mux_8503 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8504;
  function [0:0] mux_8504(input [0:0] sel);
    case (sel) 0: mux_8504 = 1'h0; 1: mux_8504 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8505;
  wire [0:0] v_8506;
  wire [0:0] v_8507;
  wire [0:0] v_8508;
  function [0:0] mux_8508(input [0:0] sel);
    case (sel) 0: mux_8508 = 1'h0; 1: mux_8508 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8509;
  function [0:0] mux_8509(input [0:0] sel);
    case (sel) 0: mux_8509 = 1'h0; 1: mux_8509 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8510;
  wire [0:0] v_8511;
  wire [0:0] v_8512;
  wire [0:0] v_8513;
  wire [0:0] v_8514;
  wire [0:0] v_8515;
  function [0:0] mux_8515(input [0:0] sel);
    case (sel) 0: mux_8515 = 1'h0; 1: mux_8515 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8516;
  wire [0:0] v_8517;
  function [0:0] mux_8517(input [0:0] sel);
    case (sel) 0: mux_8517 = 1'h0; 1: mux_8517 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8518;
  wire [0:0] v_8519;
  wire [0:0] v_8520;
  wire [0:0] v_8521;
  function [0:0] mux_8521(input [0:0] sel);
    case (sel) 0: mux_8521 = 1'h0; 1: mux_8521 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8522;
  function [0:0] mux_8522(input [0:0] sel);
    case (sel) 0: mux_8522 = 1'h0; 1: mux_8522 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8523 = 1'h0;
  wire [0:0] v_8524;
  wire [0:0] v_8525;
  wire [0:0] act_8526;
  wire [0:0] v_8527;
  wire [0:0] v_8528;
  wire [0:0] v_8529;
  reg [0:0] v_8530 = 1'h0;
  wire [0:0] v_8531;
  wire [0:0] v_8532;
  wire [0:0] act_8533;
  wire [0:0] v_8534;
  wire [0:0] v_8535;
  wire [0:0] v_8536;
  reg [0:0] v_8537 = 1'h0;
  wire [0:0] v_8538;
  wire [0:0] v_8539;
  wire [0:0] act_8540;
  wire [0:0] v_8541;
  wire [0:0] v_8542;
  wire [0:0] v_8543;
  reg [0:0] v_8544 = 1'h0;
  wire [0:0] v_8545;
  wire [0:0] v_8546;
  wire [0:0] act_8547;
  wire [0:0] v_8548;
  wire [0:0] v_8549;
  wire [0:0] v_8550;
  wire [0:0] v_8551;
  wire [0:0] v_8552;
  wire [0:0] v_8553;
  function [0:0] mux_8553(input [0:0] sel);
    case (sel) 0: mux_8553 = 1'h0; 1: mux_8553 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8554;
  wire [0:0] v_8555;
  function [0:0] mux_8555(input [0:0] sel);
    case (sel) 0: mux_8555 = 1'h0; 1: mux_8555 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8556;
  wire [0:0] v_8557;
  wire [0:0] v_8558;
  wire [0:0] v_8559;
  function [0:0] mux_8559(input [0:0] sel);
    case (sel) 0: mux_8559 = 1'h0; 1: mux_8559 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8560;
  function [0:0] mux_8560(input [0:0] sel);
    case (sel) 0: mux_8560 = 1'h0; 1: mux_8560 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8561 = 1'h0;
  wire [0:0] v_8562;
  wire [0:0] v_8563;
  wire [0:0] act_8564;
  wire [0:0] v_8565;
  wire [0:0] v_8566;
  wire [0:0] v_8567;
  wire [0:0] v_8568;
  wire [0:0] v_8569;
  wire [0:0] v_8570;
  function [0:0] mux_8570(input [0:0] sel);
    case (sel) 0: mux_8570 = 1'h0; 1: mux_8570 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8571;
  function [0:0] mux_8571(input [0:0] sel);
    case (sel) 0: mux_8571 = 1'h0; 1: mux_8571 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8572;
  wire [0:0] v_8573;
  wire [0:0] v_8574;
  wire [0:0] v_8575;
  function [0:0] mux_8575(input [0:0] sel);
    case (sel) 0: mux_8575 = 1'h0; 1: mux_8575 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8576;
  function [0:0] mux_8576(input [0:0] sel);
    case (sel) 0: mux_8576 = 1'h0; 1: mux_8576 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8577;
  wire [0:0] v_8578;
  wire [0:0] v_8579;
  wire [0:0] v_8580;
  wire [0:0] v_8581;
  wire [0:0] v_8582;
  function [0:0] mux_8582(input [0:0] sel);
    case (sel) 0: mux_8582 = 1'h0; 1: mux_8582 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8583;
  wire [0:0] v_8584;
  function [0:0] mux_8584(input [0:0] sel);
    case (sel) 0: mux_8584 = 1'h0; 1: mux_8584 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8585;
  wire [0:0] v_8586;
  wire [0:0] v_8587;
  wire [0:0] v_8588;
  function [0:0] mux_8588(input [0:0] sel);
    case (sel) 0: mux_8588 = 1'h0; 1: mux_8588 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8589;
  function [0:0] mux_8589(input [0:0] sel);
    case (sel) 0: mux_8589 = 1'h0; 1: mux_8589 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8590 = 1'h0;
  wire [0:0] v_8591;
  wire [0:0] v_8592;
  wire [0:0] act_8593;
  wire [0:0] v_8594;
  wire [0:0] v_8595;
  wire [0:0] v_8596;
  reg [0:0] v_8597 = 1'h0;
  wire [0:0] v_8598;
  wire [0:0] v_8599;
  wire [0:0] act_8600;
  wire [0:0] v_8601;
  wire [0:0] v_8602;
  wire [0:0] v_8603;
  wire [0:0] v_8604;
  wire [0:0] v_8605;
  wire [0:0] v_8606;
  function [0:0] mux_8606(input [0:0] sel);
    case (sel) 0: mux_8606 = 1'h0; 1: mux_8606 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8607;
  wire [0:0] v_8608;
  function [0:0] mux_8608(input [0:0] sel);
    case (sel) 0: mux_8608 = 1'h0; 1: mux_8608 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8609;
  wire [0:0] v_8610;
  wire [0:0] v_8611;
  wire [0:0] v_8612;
  function [0:0] mux_8612(input [0:0] sel);
    case (sel) 0: mux_8612 = 1'h0; 1: mux_8612 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8613;
  function [0:0] mux_8613(input [0:0] sel);
    case (sel) 0: mux_8613 = 1'h0; 1: mux_8613 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8614 = 1'h0;
  wire [0:0] v_8615;
  wire [0:0] v_8616;
  wire [0:0] act_8617;
  wire [0:0] v_8618;
  wire [0:0] v_8619;
  wire [0:0] v_8620;
  wire [0:0] v_8621;
  wire [0:0] v_8622;
  wire [0:0] v_8623;
  function [0:0] mux_8623(input [0:0] sel);
    case (sel) 0: mux_8623 = 1'h0; 1: mux_8623 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8624;
  function [0:0] mux_8624(input [0:0] sel);
    case (sel) 0: mux_8624 = 1'h0; 1: mux_8624 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8625;
  wire [0:0] v_8626;
  wire [0:0] v_8627;
  wire [0:0] v_8628;
  function [0:0] mux_8628(input [0:0] sel);
    case (sel) 0: mux_8628 = 1'h0; 1: mux_8628 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8629;
  function [0:0] mux_8629(input [0:0] sel);
    case (sel) 0: mux_8629 = 1'h0; 1: mux_8629 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8630;
  wire [0:0] v_8631;
  wire [0:0] v_8632;
  wire [0:0] v_8633;
  wire [0:0] v_8634;
  wire [0:0] v_8635;
  function [0:0] mux_8635(input [0:0] sel);
    case (sel) 0: mux_8635 = 1'h0; 1: mux_8635 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8636;
  function [0:0] mux_8636(input [0:0] sel);
    case (sel) 0: mux_8636 = 1'h0; 1: mux_8636 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8637;
  wire [0:0] v_8638;
  wire [0:0] v_8639;
  wire [0:0] v_8640;
  function [0:0] mux_8640(input [0:0] sel);
    case (sel) 0: mux_8640 = 1'h0; 1: mux_8640 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8641;
  function [0:0] mux_8641(input [0:0] sel);
    case (sel) 0: mux_8641 = 1'h0; 1: mux_8641 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8642;
  wire [0:0] v_8643;
  wire [0:0] v_8644;
  wire [0:0] v_8645;
  wire [0:0] v_8646;
  wire [0:0] v_8647;
  function [0:0] mux_8647(input [0:0] sel);
    case (sel) 0: mux_8647 = 1'h0; 1: mux_8647 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8648;
  wire [0:0] v_8649;
  function [0:0] mux_8649(input [0:0] sel);
    case (sel) 0: mux_8649 = 1'h0; 1: mux_8649 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8650;
  wire [0:0] v_8651;
  wire [0:0] v_8652;
  wire [0:0] v_8653;
  function [0:0] mux_8653(input [0:0] sel);
    case (sel) 0: mux_8653 = 1'h0; 1: mux_8653 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8654;
  function [0:0] mux_8654(input [0:0] sel);
    case (sel) 0: mux_8654 = 1'h0; 1: mux_8654 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8655 = 1'h0;
  wire [0:0] v_8656;
  wire [0:0] v_8657;
  wire [0:0] act_8658;
  wire [0:0] v_8659;
  wire [0:0] v_8660;
  wire [0:0] v_8661;
  reg [0:0] v_8662 = 1'h0;
  wire [0:0] v_8663;
  wire [0:0] v_8664;
  wire [0:0] act_8665;
  wire [0:0] v_8666;
  wire [0:0] v_8667;
  wire [0:0] v_8668;
  reg [0:0] v_8669 = 1'h0;
  wire [0:0] v_8670;
  wire [0:0] v_8671;
  wire [0:0] act_8672;
  wire [0:0] v_8673;
  wire [0:0] v_8674;
  wire [0:0] v_8675;
  wire [0:0] v_8676;
  wire [0:0] v_8677;
  wire [0:0] v_8678;
  function [0:0] mux_8678(input [0:0] sel);
    case (sel) 0: mux_8678 = 1'h0; 1: mux_8678 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8679;
  wire [0:0] v_8680;
  function [0:0] mux_8680(input [0:0] sel);
    case (sel) 0: mux_8680 = 1'h0; 1: mux_8680 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8681;
  wire [0:0] v_8682;
  wire [0:0] v_8683;
  wire [0:0] v_8684;
  function [0:0] mux_8684(input [0:0] sel);
    case (sel) 0: mux_8684 = 1'h0; 1: mux_8684 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8685;
  function [0:0] mux_8685(input [0:0] sel);
    case (sel) 0: mux_8685 = 1'h0; 1: mux_8685 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8686 = 1'h0;
  wire [0:0] v_8687;
  wire [0:0] v_8688;
  wire [0:0] act_8689;
  wire [0:0] v_8690;
  wire [0:0] v_8691;
  wire [0:0] v_8692;
  wire [0:0] v_8693;
  wire [0:0] v_8694;
  wire [0:0] v_8695;
  function [0:0] mux_8695(input [0:0] sel);
    case (sel) 0: mux_8695 = 1'h0; 1: mux_8695 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8696;
  function [0:0] mux_8696(input [0:0] sel);
    case (sel) 0: mux_8696 = 1'h0; 1: mux_8696 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8697;
  wire [0:0] v_8698;
  wire [0:0] v_8699;
  wire [0:0] v_8700;
  function [0:0] mux_8700(input [0:0] sel);
    case (sel) 0: mux_8700 = 1'h0; 1: mux_8700 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8701;
  function [0:0] mux_8701(input [0:0] sel);
    case (sel) 0: mux_8701 = 1'h0; 1: mux_8701 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8702;
  wire [0:0] v_8703;
  wire [0:0] v_8704;
  wire [0:0] v_8705;
  wire [0:0] v_8706;
  wire [0:0] v_8707;
  function [0:0] mux_8707(input [0:0] sel);
    case (sel) 0: mux_8707 = 1'h0; 1: mux_8707 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8708;
  wire [0:0] v_8709;
  function [0:0] mux_8709(input [0:0] sel);
    case (sel) 0: mux_8709 = 1'h0; 1: mux_8709 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8710;
  wire [0:0] v_8711;
  wire [0:0] v_8712;
  wire [0:0] v_8713;
  function [0:0] mux_8713(input [0:0] sel);
    case (sel) 0: mux_8713 = 1'h0; 1: mux_8713 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8714;
  function [0:0] mux_8714(input [0:0] sel);
    case (sel) 0: mux_8714 = 1'h0; 1: mux_8714 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8715 = 1'h0;
  wire [0:0] v_8716;
  wire [0:0] v_8717;
  wire [0:0] act_8718;
  wire [0:0] v_8719;
  wire [0:0] v_8720;
  wire [0:0] v_8721;
  reg [0:0] v_8722 = 1'h0;
  wire [0:0] v_8723;
  wire [0:0] v_8724;
  wire [0:0] act_8725;
  wire [0:0] v_8726;
  wire [0:0] v_8727;
  wire [0:0] v_8728;
  wire [0:0] v_8729;
  wire [0:0] v_8730;
  wire [0:0] v_8731;
  function [0:0] mux_8731(input [0:0] sel);
    case (sel) 0: mux_8731 = 1'h0; 1: mux_8731 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8732;
  wire [0:0] v_8733;
  function [0:0] mux_8733(input [0:0] sel);
    case (sel) 0: mux_8733 = 1'h0; 1: mux_8733 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8734;
  wire [0:0] v_8735;
  wire [0:0] v_8736;
  wire [0:0] v_8737;
  function [0:0] mux_8737(input [0:0] sel);
    case (sel) 0: mux_8737 = 1'h0; 1: mux_8737 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8738;
  function [0:0] mux_8738(input [0:0] sel);
    case (sel) 0: mux_8738 = 1'h0; 1: mux_8738 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8739 = 1'h0;
  wire [0:0] v_8740;
  wire [0:0] v_8741;
  wire [0:0] act_8742;
  wire [0:0] v_8743;
  wire [0:0] v_8744;
  wire [0:0] v_8745;
  wire [0:0] v_8746;
  wire [0:0] v_8747;
  wire [0:0] v_8748;
  function [0:0] mux_8748(input [0:0] sel);
    case (sel) 0: mux_8748 = 1'h0; 1: mux_8748 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8749;
  function [0:0] mux_8749(input [0:0] sel);
    case (sel) 0: mux_8749 = 1'h0; 1: mux_8749 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8750;
  wire [0:0] v_8751;
  wire [0:0] v_8752;
  wire [0:0] v_8753;
  function [0:0] mux_8753(input [0:0] sel);
    case (sel) 0: mux_8753 = 1'h0; 1: mux_8753 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8754;
  function [0:0] mux_8754(input [0:0] sel);
    case (sel) 0: mux_8754 = 1'h0; 1: mux_8754 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8755;
  wire [0:0] v_8756;
  wire [0:0] v_8757;
  wire [0:0] v_8758;
  wire [0:0] v_8759;
  wire [0:0] v_8760;
  function [0:0] mux_8760(input [0:0] sel);
    case (sel) 0: mux_8760 = 1'h0; 1: mux_8760 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8761;
  function [0:0] mux_8761(input [0:0] sel);
    case (sel) 0: mux_8761 = 1'h0; 1: mux_8761 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8762;
  wire [0:0] v_8763;
  wire [0:0] v_8764;
  wire [0:0] v_8765;
  function [0:0] mux_8765(input [0:0] sel);
    case (sel) 0: mux_8765 = 1'h0; 1: mux_8765 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8766;
  function [0:0] mux_8766(input [0:0] sel);
    case (sel) 0: mux_8766 = 1'h0; 1: mux_8766 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8767;
  wire [0:0] v_8768;
  wire [0:0] v_8769;
  wire [0:0] v_8770;
  wire [0:0] v_8771;
  wire [0:0] v_8772;
  function [0:0] mux_8772(input [0:0] sel);
    case (sel) 0: mux_8772 = 1'h0; 1: mux_8772 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8773;
  function [0:0] mux_8773(input [0:0] sel);
    case (sel) 0: mux_8773 = 1'h0; 1: mux_8773 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8774;
  wire [0:0] v_8775;
  wire [0:0] v_8776;
  wire [0:0] v_8777;
  function [0:0] mux_8777(input [0:0] sel);
    case (sel) 0: mux_8777 = 1'h0; 1: mux_8777 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8778;
  function [0:0] mux_8778(input [0:0] sel);
    case (sel) 0: mux_8778 = 1'h0; 1: mux_8778 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8779;
  wire [0:0] v_8780;
  wire [0:0] v_8781;
  wire [0:0] v_8782;
  wire [0:0] v_8783;
  wire [0:0] v_8784;
  function [0:0] mux_8784(input [0:0] sel);
    case (sel) 0: mux_8784 = 1'h0; 1: mux_8784 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8785;
  function [0:0] mux_8785(input [0:0] sel);
    case (sel) 0: mux_8785 = 1'h0; 1: mux_8785 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8786;
  wire [0:0] v_8787;
  wire [0:0] v_8788;
  wire [0:0] v_8789;
  function [0:0] mux_8789(input [0:0] sel);
    case (sel) 0: mux_8789 = 1'h0; 1: mux_8789 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8790;
  function [0:0] mux_8790(input [0:0] sel);
    case (sel) 0: mux_8790 = 1'h0; 1: mux_8790 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8791;
  wire [0:0] v_8792;
  wire [0:0] v_8793;
  wire [0:0] v_8794;
  wire [0:0] v_8795;
  wire [0:0] v_8796;
  function [0:0] mux_8796(input [0:0] sel);
    case (sel) 0: mux_8796 = 1'h0; 1: mux_8796 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8797;
  function [0:0] mux_8797(input [0:0] sel);
    case (sel) 0: mux_8797 = 1'h0; 1: mux_8797 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8798;
  wire [0:0] v_8799;
  wire [0:0] v_8800;
  wire [0:0] v_8801;
  function [0:0] mux_8801(input [0:0] sel);
    case (sel) 0: mux_8801 = 1'h0; 1: mux_8801 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8802;
  function [0:0] mux_8802(input [0:0] sel);
    case (sel) 0: mux_8802 = 1'h0; 1: mux_8802 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8803;
  wire [0:0] v_8804;
  wire [0:0] v_8805;
  wire [0:0] v_8806;
  wire [0:0] v_8807;
  wire [0:0] v_8808;
  function [0:0] mux_8808(input [0:0] sel);
    case (sel) 0: mux_8808 = 1'h0; 1: mux_8808 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8809;
  wire [0:0] v_8810;
  function [0:0] mux_8810(input [0:0] sel);
    case (sel) 0: mux_8810 = 1'h0; 1: mux_8810 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8811;
  wire [0:0] v_8812;
  wire [0:0] v_8813;
  wire [0:0] v_8814;
  function [0:0] mux_8814(input [0:0] sel);
    case (sel) 0: mux_8814 = 1'h0; 1: mux_8814 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8815;
  function [0:0] mux_8815(input [0:0] sel);
    case (sel) 0: mux_8815 = 1'h0; 1: mux_8815 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8816 = 1'h0;
  wire [0:0] v_8817;
  wire [0:0] v_8818;
  wire [0:0] act_8819;
  wire [0:0] v_8820;
  wire [0:0] v_8821;
  wire [0:0] v_8822;
  reg [0:0] v_8823 = 1'h0;
  wire [0:0] v_8824;
  wire [0:0] v_8825;
  wire [0:0] act_8826;
  wire [0:0] v_8827;
  wire [0:0] v_8828;
  wire [0:0] v_8829;
  reg [0:0] v_8830 = 1'h0;
  wire [0:0] v_8831;
  wire [0:0] v_8832;
  wire [0:0] act_8833;
  wire [0:0] v_8834;
  wire [0:0] v_8835;
  wire [0:0] v_8836;
  reg [0:0] v_8837 = 1'h0;
  wire [0:0] v_8838;
  wire [0:0] v_8839;
  wire [0:0] act_8840;
  wire [0:0] v_8841;
  wire [0:0] v_8842;
  wire [0:0] v_8843;
  reg [0:0] v_8844 = 1'h0;
  wire [0:0] v_8845;
  wire [0:0] v_8846;
  wire [0:0] act_8847;
  wire [0:0] v_8848;
  wire [0:0] v_8849;
  wire [0:0] v_8850;
  reg [0:0] v_8851 = 1'h0;
  wire [0:0] v_8852;
  wire [0:0] v_8853;
  wire [0:0] act_8854;
  wire [0:0] v_8855;
  wire [0:0] v_8856;
  wire [0:0] v_8857;
  wire [0:0] v_8858;
  wire [0:0] v_8859;
  wire [0:0] v_8860;
  function [0:0] mux_8860(input [0:0] sel);
    case (sel) 0: mux_8860 = 1'h0; 1: mux_8860 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8861;
  wire [0:0] v_8862;
  function [0:0] mux_8862(input [0:0] sel);
    case (sel) 0: mux_8862 = 1'h0; 1: mux_8862 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8863;
  wire [0:0] v_8864;
  wire [0:0] v_8865;
  wire [0:0] v_8866;
  function [0:0] mux_8866(input [0:0] sel);
    case (sel) 0: mux_8866 = 1'h0; 1: mux_8866 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8867;
  function [0:0] mux_8867(input [0:0] sel);
    case (sel) 0: mux_8867 = 1'h0; 1: mux_8867 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8868 = 1'h0;
  wire [0:0] v_8869;
  wire [0:0] v_8870;
  wire [0:0] act_8871;
  wire [0:0] v_8872;
  wire [0:0] v_8873;
  wire [0:0] v_8874;
  wire [0:0] v_8875;
  wire [0:0] v_8876;
  wire [0:0] v_8877;
  function [0:0] mux_8877(input [0:0] sel);
    case (sel) 0: mux_8877 = 1'h0; 1: mux_8877 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8878;
  function [0:0] mux_8878(input [0:0] sel);
    case (sel) 0: mux_8878 = 1'h0; 1: mux_8878 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8879;
  wire [0:0] v_8880;
  wire [0:0] v_8881;
  wire [0:0] v_8882;
  function [0:0] mux_8882(input [0:0] sel);
    case (sel) 0: mux_8882 = 1'h0; 1: mux_8882 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8883;
  function [0:0] mux_8883(input [0:0] sel);
    case (sel) 0: mux_8883 = 1'h0; 1: mux_8883 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8884;
  wire [0:0] v_8885;
  wire [0:0] v_8886;
  wire [0:0] v_8887;
  wire [0:0] v_8888;
  wire [0:0] v_8889;
  function [0:0] mux_8889(input [0:0] sel);
    case (sel) 0: mux_8889 = 1'h0; 1: mux_8889 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8890;
  wire [0:0] v_8891;
  function [0:0] mux_8891(input [0:0] sel);
    case (sel) 0: mux_8891 = 1'h0; 1: mux_8891 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8892;
  wire [0:0] v_8893;
  wire [0:0] v_8894;
  wire [0:0] v_8895;
  function [0:0] mux_8895(input [0:0] sel);
    case (sel) 0: mux_8895 = 1'h0; 1: mux_8895 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8896;
  function [0:0] mux_8896(input [0:0] sel);
    case (sel) 0: mux_8896 = 1'h0; 1: mux_8896 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8897 = 1'h0;
  wire [0:0] v_8898;
  wire [0:0] v_8899;
  wire [0:0] act_8900;
  wire [0:0] v_8901;
  wire [0:0] v_8902;
  wire [0:0] v_8903;
  reg [0:0] v_8904 = 1'h0;
  wire [0:0] v_8905;
  wire [0:0] v_8906;
  wire [0:0] act_8907;
  wire [0:0] v_8908;
  wire [0:0] v_8909;
  wire [0:0] v_8910;
  wire [0:0] v_8911;
  wire [0:0] v_8912;
  wire [0:0] v_8913;
  function [0:0] mux_8913(input [0:0] sel);
    case (sel) 0: mux_8913 = 1'h0; 1: mux_8913 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8914;
  wire [0:0] v_8915;
  function [0:0] mux_8915(input [0:0] sel);
    case (sel) 0: mux_8915 = 1'h0; 1: mux_8915 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8916;
  wire [0:0] v_8917;
  wire [0:0] v_8918;
  wire [0:0] v_8919;
  function [0:0] mux_8919(input [0:0] sel);
    case (sel) 0: mux_8919 = 1'h0; 1: mux_8919 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8920;
  function [0:0] mux_8920(input [0:0] sel);
    case (sel) 0: mux_8920 = 1'h0; 1: mux_8920 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8921 = 1'h0;
  wire [0:0] v_8922;
  wire [0:0] v_8923;
  wire [0:0] act_8924;
  wire [0:0] v_8925;
  wire [0:0] v_8926;
  wire [0:0] v_8927;
  wire [0:0] v_8928;
  wire [0:0] v_8929;
  wire [0:0] v_8930;
  function [0:0] mux_8930(input [0:0] sel);
    case (sel) 0: mux_8930 = 1'h0; 1: mux_8930 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8931;
  function [0:0] mux_8931(input [0:0] sel);
    case (sel) 0: mux_8931 = 1'h0; 1: mux_8931 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8932;
  wire [0:0] v_8933;
  wire [0:0] v_8934;
  wire [0:0] v_8935;
  function [0:0] mux_8935(input [0:0] sel);
    case (sel) 0: mux_8935 = 1'h0; 1: mux_8935 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8936;
  function [0:0] mux_8936(input [0:0] sel);
    case (sel) 0: mux_8936 = 1'h0; 1: mux_8936 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8937;
  wire [0:0] v_8938;
  wire [0:0] v_8939;
  wire [0:0] v_8940;
  wire [0:0] v_8941;
  wire [0:0] v_8942;
  function [0:0] mux_8942(input [0:0] sel);
    case (sel) 0: mux_8942 = 1'h0; 1: mux_8942 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8943;
  function [0:0] mux_8943(input [0:0] sel);
    case (sel) 0: mux_8943 = 1'h0; 1: mux_8943 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8944;
  wire [0:0] v_8945;
  wire [0:0] v_8946;
  wire [0:0] v_8947;
  function [0:0] mux_8947(input [0:0] sel);
    case (sel) 0: mux_8947 = 1'h0; 1: mux_8947 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8948;
  function [0:0] mux_8948(input [0:0] sel);
    case (sel) 0: mux_8948 = 1'h0; 1: mux_8948 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8949;
  wire [0:0] v_8950;
  wire [0:0] v_8951;
  wire [0:0] v_8952;
  wire [0:0] v_8953;
  wire [0:0] v_8954;
  function [0:0] mux_8954(input [0:0] sel);
    case (sel) 0: mux_8954 = 1'h0; 1: mux_8954 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8955;
  wire [0:0] v_8956;
  function [0:0] mux_8956(input [0:0] sel);
    case (sel) 0: mux_8956 = 1'h0; 1: mux_8956 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8957;
  wire [0:0] v_8958;
  wire [0:0] v_8959;
  wire [0:0] v_8960;
  function [0:0] mux_8960(input [0:0] sel);
    case (sel) 0: mux_8960 = 1'h0; 1: mux_8960 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8961;
  function [0:0] mux_8961(input [0:0] sel);
    case (sel) 0: mux_8961 = 1'h0; 1: mux_8961 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8962 = 1'h0;
  wire [0:0] v_8963;
  wire [0:0] v_8964;
  wire [0:0] act_8965;
  wire [0:0] v_8966;
  wire [0:0] v_8967;
  wire [0:0] v_8968;
  reg [0:0] v_8969 = 1'h0;
  wire [0:0] v_8970;
  wire [0:0] v_8971;
  wire [0:0] act_8972;
  wire [0:0] v_8973;
  wire [0:0] v_8974;
  wire [0:0] v_8975;
  reg [0:0] v_8976 = 1'h0;
  wire [0:0] v_8977;
  wire [0:0] v_8978;
  wire [0:0] act_8979;
  wire [0:0] v_8980;
  wire [0:0] v_8981;
  wire [0:0] v_8982;
  wire [0:0] v_8983;
  wire [0:0] v_8984;
  wire [0:0] v_8985;
  function [0:0] mux_8985(input [0:0] sel);
    case (sel) 0: mux_8985 = 1'h0; 1: mux_8985 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8986;
  wire [0:0] v_8987;
  function [0:0] mux_8987(input [0:0] sel);
    case (sel) 0: mux_8987 = 1'h0; 1: mux_8987 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_8988;
  wire [0:0] v_8989;
  wire [0:0] v_8990;
  wire [0:0] v_8991;
  function [0:0] mux_8991(input [0:0] sel);
    case (sel) 0: mux_8991 = 1'h0; 1: mux_8991 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_8992;
  function [0:0] mux_8992(input [0:0] sel);
    case (sel) 0: mux_8992 = 1'h0; 1: mux_8992 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_8993 = 1'h0;
  wire [0:0] v_8994;
  wire [0:0] v_8995;
  wire [0:0] act_8996;
  wire [0:0] v_8997;
  wire [0:0] v_8998;
  wire [0:0] v_8999;
  wire [0:0] v_9000;
  wire [0:0] v_9001;
  wire [0:0] v_9002;
  function [0:0] mux_9002(input [0:0] sel);
    case (sel) 0: mux_9002 = 1'h0; 1: mux_9002 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9003;
  function [0:0] mux_9003(input [0:0] sel);
    case (sel) 0: mux_9003 = 1'h0; 1: mux_9003 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9004;
  wire [0:0] v_9005;
  wire [0:0] v_9006;
  wire [0:0] v_9007;
  function [0:0] mux_9007(input [0:0] sel);
    case (sel) 0: mux_9007 = 1'h0; 1: mux_9007 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9008;
  function [0:0] mux_9008(input [0:0] sel);
    case (sel) 0: mux_9008 = 1'h0; 1: mux_9008 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9009;
  wire [0:0] v_9010;
  wire [0:0] v_9011;
  wire [0:0] v_9012;
  wire [0:0] v_9013;
  wire [0:0] v_9014;
  function [0:0] mux_9014(input [0:0] sel);
    case (sel) 0: mux_9014 = 1'h0; 1: mux_9014 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9015;
  wire [0:0] v_9016;
  function [0:0] mux_9016(input [0:0] sel);
    case (sel) 0: mux_9016 = 1'h0; 1: mux_9016 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9017;
  wire [0:0] v_9018;
  wire [0:0] v_9019;
  wire [0:0] v_9020;
  function [0:0] mux_9020(input [0:0] sel);
    case (sel) 0: mux_9020 = 1'h0; 1: mux_9020 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9021;
  function [0:0] mux_9021(input [0:0] sel);
    case (sel) 0: mux_9021 = 1'h0; 1: mux_9021 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9022 = 1'h0;
  wire [0:0] v_9023;
  wire [0:0] v_9024;
  wire [0:0] act_9025;
  wire [0:0] v_9026;
  wire [0:0] v_9027;
  wire [0:0] v_9028;
  reg [0:0] v_9029 = 1'h0;
  wire [0:0] v_9030;
  wire [0:0] v_9031;
  wire [0:0] act_9032;
  wire [0:0] v_9033;
  wire [0:0] v_9034;
  wire [0:0] v_9035;
  wire [0:0] v_9036;
  wire [0:0] v_9037;
  wire [0:0] v_9038;
  function [0:0] mux_9038(input [0:0] sel);
    case (sel) 0: mux_9038 = 1'h0; 1: mux_9038 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9039;
  wire [0:0] v_9040;
  function [0:0] mux_9040(input [0:0] sel);
    case (sel) 0: mux_9040 = 1'h0; 1: mux_9040 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9041;
  wire [0:0] v_9042;
  wire [0:0] v_9043;
  wire [0:0] v_9044;
  function [0:0] mux_9044(input [0:0] sel);
    case (sel) 0: mux_9044 = 1'h0; 1: mux_9044 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9045;
  function [0:0] mux_9045(input [0:0] sel);
    case (sel) 0: mux_9045 = 1'h0; 1: mux_9045 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9046 = 1'h0;
  wire [0:0] v_9047;
  wire [0:0] v_9048;
  wire [0:0] act_9049;
  wire [0:0] v_9050;
  wire [0:0] v_9051;
  wire [0:0] v_9052;
  wire [0:0] v_9053;
  wire [0:0] v_9054;
  wire [0:0] v_9055;
  function [0:0] mux_9055(input [0:0] sel);
    case (sel) 0: mux_9055 = 1'h0; 1: mux_9055 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9056;
  function [0:0] mux_9056(input [0:0] sel);
    case (sel) 0: mux_9056 = 1'h0; 1: mux_9056 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9057;
  wire [0:0] v_9058;
  wire [0:0] v_9059;
  wire [0:0] v_9060;
  function [0:0] mux_9060(input [0:0] sel);
    case (sel) 0: mux_9060 = 1'h0; 1: mux_9060 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9061;
  function [0:0] mux_9061(input [0:0] sel);
    case (sel) 0: mux_9061 = 1'h0; 1: mux_9061 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9062;
  wire [0:0] v_9063;
  wire [0:0] v_9064;
  wire [0:0] v_9065;
  wire [0:0] v_9066;
  wire [0:0] v_9067;
  function [0:0] mux_9067(input [0:0] sel);
    case (sel) 0: mux_9067 = 1'h0; 1: mux_9067 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9068;
  function [0:0] mux_9068(input [0:0] sel);
    case (sel) 0: mux_9068 = 1'h0; 1: mux_9068 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9069;
  wire [0:0] v_9070;
  wire [0:0] v_9071;
  wire [0:0] v_9072;
  function [0:0] mux_9072(input [0:0] sel);
    case (sel) 0: mux_9072 = 1'h0; 1: mux_9072 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9073;
  function [0:0] mux_9073(input [0:0] sel);
    case (sel) 0: mux_9073 = 1'h0; 1: mux_9073 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9074;
  wire [0:0] v_9075;
  wire [0:0] v_9076;
  wire [0:0] v_9077;
  wire [0:0] v_9078;
  wire [0:0] v_9079;
  function [0:0] mux_9079(input [0:0] sel);
    case (sel) 0: mux_9079 = 1'h0; 1: mux_9079 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9080;
  function [0:0] mux_9080(input [0:0] sel);
    case (sel) 0: mux_9080 = 1'h0; 1: mux_9080 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9081;
  wire [0:0] v_9082;
  wire [0:0] v_9083;
  wire [0:0] v_9084;
  function [0:0] mux_9084(input [0:0] sel);
    case (sel) 0: mux_9084 = 1'h0; 1: mux_9084 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9085;
  function [0:0] mux_9085(input [0:0] sel);
    case (sel) 0: mux_9085 = 1'h0; 1: mux_9085 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9086;
  wire [0:0] v_9087;
  wire [0:0] v_9088;
  wire [0:0] v_9089;
  wire [0:0] v_9090;
  wire [0:0] v_9091;
  function [0:0] mux_9091(input [0:0] sel);
    case (sel) 0: mux_9091 = 1'h0; 1: mux_9091 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9092;
  wire [0:0] v_9093;
  function [0:0] mux_9093(input [0:0] sel);
    case (sel) 0: mux_9093 = 1'h0; 1: mux_9093 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9094;
  wire [0:0] v_9095;
  wire [0:0] v_9096;
  wire [0:0] v_9097;
  function [0:0] mux_9097(input [0:0] sel);
    case (sel) 0: mux_9097 = 1'h0; 1: mux_9097 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9098;
  function [0:0] mux_9098(input [0:0] sel);
    case (sel) 0: mux_9098 = 1'h0; 1: mux_9098 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9099 = 1'h0;
  wire [0:0] v_9100;
  wire [0:0] v_9101;
  wire [0:0] act_9102;
  wire [0:0] v_9103;
  wire [0:0] v_9104;
  wire [0:0] v_9105;
  reg [0:0] v_9106 = 1'h0;
  wire [0:0] v_9107;
  wire [0:0] v_9108;
  wire [0:0] act_9109;
  wire [0:0] v_9110;
  wire [0:0] v_9111;
  wire [0:0] v_9112;
  reg [0:0] v_9113 = 1'h0;
  wire [0:0] v_9114;
  wire [0:0] v_9115;
  wire [0:0] act_9116;
  wire [0:0] v_9117;
  wire [0:0] v_9118;
  wire [0:0] v_9119;
  reg [0:0] v_9120 = 1'h0;
  wire [0:0] v_9121;
  wire [0:0] v_9122;
  wire [0:0] act_9123;
  wire [0:0] v_9124;
  wire [0:0] v_9125;
  wire [0:0] v_9126;
  wire [0:0] v_9127;
  wire [0:0] v_9128;
  wire [0:0] v_9129;
  function [0:0] mux_9129(input [0:0] sel);
    case (sel) 0: mux_9129 = 1'h0; 1: mux_9129 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9130;
  wire [0:0] v_9131;
  function [0:0] mux_9131(input [0:0] sel);
    case (sel) 0: mux_9131 = 1'h0; 1: mux_9131 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9132;
  wire [0:0] v_9133;
  wire [0:0] v_9134;
  wire [0:0] v_9135;
  function [0:0] mux_9135(input [0:0] sel);
    case (sel) 0: mux_9135 = 1'h0; 1: mux_9135 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9136;
  function [0:0] mux_9136(input [0:0] sel);
    case (sel) 0: mux_9136 = 1'h0; 1: mux_9136 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9137 = 1'h0;
  wire [0:0] v_9138;
  wire [0:0] v_9139;
  wire [0:0] act_9140;
  wire [0:0] v_9141;
  wire [0:0] v_9142;
  wire [0:0] v_9143;
  wire [0:0] v_9144;
  wire [0:0] v_9145;
  wire [0:0] v_9146;
  function [0:0] mux_9146(input [0:0] sel);
    case (sel) 0: mux_9146 = 1'h0; 1: mux_9146 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9147;
  function [0:0] mux_9147(input [0:0] sel);
    case (sel) 0: mux_9147 = 1'h0; 1: mux_9147 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9148;
  wire [0:0] v_9149;
  wire [0:0] v_9150;
  wire [0:0] v_9151;
  function [0:0] mux_9151(input [0:0] sel);
    case (sel) 0: mux_9151 = 1'h0; 1: mux_9151 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9152;
  function [0:0] mux_9152(input [0:0] sel);
    case (sel) 0: mux_9152 = 1'h0; 1: mux_9152 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9153;
  wire [0:0] v_9154;
  wire [0:0] v_9155;
  wire [0:0] v_9156;
  wire [0:0] v_9157;
  wire [0:0] v_9158;
  function [0:0] mux_9158(input [0:0] sel);
    case (sel) 0: mux_9158 = 1'h0; 1: mux_9158 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9159;
  wire [0:0] v_9160;
  function [0:0] mux_9160(input [0:0] sel);
    case (sel) 0: mux_9160 = 1'h0; 1: mux_9160 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9161;
  wire [0:0] v_9162;
  wire [0:0] v_9163;
  wire [0:0] v_9164;
  function [0:0] mux_9164(input [0:0] sel);
    case (sel) 0: mux_9164 = 1'h0; 1: mux_9164 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9165;
  function [0:0] mux_9165(input [0:0] sel);
    case (sel) 0: mux_9165 = 1'h0; 1: mux_9165 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9166 = 1'h0;
  wire [0:0] v_9167;
  wire [0:0] v_9168;
  wire [0:0] act_9169;
  wire [0:0] v_9170;
  wire [0:0] v_9171;
  wire [0:0] v_9172;
  reg [0:0] v_9173 = 1'h0;
  wire [0:0] v_9174;
  wire [0:0] v_9175;
  wire [0:0] act_9176;
  wire [0:0] v_9177;
  wire [0:0] v_9178;
  wire [0:0] v_9179;
  wire [0:0] v_9180;
  wire [0:0] v_9181;
  wire [0:0] v_9182;
  function [0:0] mux_9182(input [0:0] sel);
    case (sel) 0: mux_9182 = 1'h0; 1: mux_9182 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9183;
  wire [0:0] v_9184;
  function [0:0] mux_9184(input [0:0] sel);
    case (sel) 0: mux_9184 = 1'h0; 1: mux_9184 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9185;
  wire [0:0] v_9186;
  wire [0:0] v_9187;
  wire [0:0] v_9188;
  function [0:0] mux_9188(input [0:0] sel);
    case (sel) 0: mux_9188 = 1'h0; 1: mux_9188 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9189;
  function [0:0] mux_9189(input [0:0] sel);
    case (sel) 0: mux_9189 = 1'h0; 1: mux_9189 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9190 = 1'h0;
  wire [0:0] v_9191;
  wire [0:0] v_9192;
  wire [0:0] act_9193;
  wire [0:0] v_9194;
  wire [0:0] v_9195;
  wire [0:0] v_9196;
  wire [0:0] v_9197;
  wire [0:0] v_9198;
  wire [0:0] v_9199;
  function [0:0] mux_9199(input [0:0] sel);
    case (sel) 0: mux_9199 = 1'h0; 1: mux_9199 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9200;
  function [0:0] mux_9200(input [0:0] sel);
    case (sel) 0: mux_9200 = 1'h0; 1: mux_9200 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9201;
  wire [0:0] v_9202;
  wire [0:0] v_9203;
  wire [0:0] v_9204;
  function [0:0] mux_9204(input [0:0] sel);
    case (sel) 0: mux_9204 = 1'h0; 1: mux_9204 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9205;
  function [0:0] mux_9205(input [0:0] sel);
    case (sel) 0: mux_9205 = 1'h0; 1: mux_9205 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9206;
  wire [0:0] v_9207;
  wire [0:0] v_9208;
  wire [0:0] v_9209;
  wire [0:0] v_9210;
  wire [0:0] v_9211;
  function [0:0] mux_9211(input [0:0] sel);
    case (sel) 0: mux_9211 = 1'h0; 1: mux_9211 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9212;
  function [0:0] mux_9212(input [0:0] sel);
    case (sel) 0: mux_9212 = 1'h0; 1: mux_9212 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9213;
  wire [0:0] v_9214;
  wire [0:0] v_9215;
  wire [0:0] v_9216;
  function [0:0] mux_9216(input [0:0] sel);
    case (sel) 0: mux_9216 = 1'h0; 1: mux_9216 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9217;
  function [0:0] mux_9217(input [0:0] sel);
    case (sel) 0: mux_9217 = 1'h0; 1: mux_9217 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9218;
  wire [0:0] v_9219;
  wire [0:0] v_9220;
  wire [0:0] v_9221;
  wire [0:0] v_9222;
  wire [0:0] v_9223;
  function [0:0] mux_9223(input [0:0] sel);
    case (sel) 0: mux_9223 = 1'h0; 1: mux_9223 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9224;
  wire [0:0] v_9225;
  function [0:0] mux_9225(input [0:0] sel);
    case (sel) 0: mux_9225 = 1'h0; 1: mux_9225 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9226;
  wire [0:0] v_9227;
  wire [0:0] v_9228;
  wire [0:0] v_9229;
  function [0:0] mux_9229(input [0:0] sel);
    case (sel) 0: mux_9229 = 1'h0; 1: mux_9229 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9230;
  function [0:0] mux_9230(input [0:0] sel);
    case (sel) 0: mux_9230 = 1'h0; 1: mux_9230 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9231 = 1'h0;
  wire [0:0] v_9232;
  wire [0:0] v_9233;
  wire [0:0] act_9234;
  wire [0:0] v_9235;
  wire [0:0] v_9236;
  wire [0:0] v_9237;
  reg [0:0] v_9238 = 1'h0;
  wire [0:0] v_9239;
  wire [0:0] v_9240;
  wire [0:0] act_9241;
  wire [0:0] v_9242;
  wire [0:0] v_9243;
  wire [0:0] v_9244;
  reg [0:0] v_9245 = 1'h0;
  wire [0:0] v_9246;
  wire [0:0] v_9247;
  wire [0:0] act_9248;
  wire [0:0] v_9249;
  wire [0:0] v_9250;
  wire [0:0] v_9251;
  wire [0:0] v_9252;
  wire [0:0] v_9253;
  wire [0:0] v_9254;
  function [0:0] mux_9254(input [0:0] sel);
    case (sel) 0: mux_9254 = 1'h0; 1: mux_9254 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9255;
  wire [0:0] v_9256;
  function [0:0] mux_9256(input [0:0] sel);
    case (sel) 0: mux_9256 = 1'h0; 1: mux_9256 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9257;
  wire [0:0] v_9258;
  wire [0:0] v_9259;
  wire [0:0] v_9260;
  function [0:0] mux_9260(input [0:0] sel);
    case (sel) 0: mux_9260 = 1'h0; 1: mux_9260 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9261;
  function [0:0] mux_9261(input [0:0] sel);
    case (sel) 0: mux_9261 = 1'h0; 1: mux_9261 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9262 = 1'h0;
  wire [0:0] v_9263;
  wire [0:0] v_9264;
  wire [0:0] act_9265;
  wire [0:0] v_9266;
  wire [0:0] v_9267;
  wire [0:0] v_9268;
  wire [0:0] v_9269;
  wire [0:0] v_9270;
  wire [0:0] v_9271;
  function [0:0] mux_9271(input [0:0] sel);
    case (sel) 0: mux_9271 = 1'h0; 1: mux_9271 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9272;
  function [0:0] mux_9272(input [0:0] sel);
    case (sel) 0: mux_9272 = 1'h0; 1: mux_9272 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9273;
  wire [0:0] v_9274;
  wire [0:0] v_9275;
  wire [0:0] v_9276;
  function [0:0] mux_9276(input [0:0] sel);
    case (sel) 0: mux_9276 = 1'h0; 1: mux_9276 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9277;
  function [0:0] mux_9277(input [0:0] sel);
    case (sel) 0: mux_9277 = 1'h0; 1: mux_9277 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9278;
  wire [0:0] v_9279;
  wire [0:0] v_9280;
  wire [0:0] v_9281;
  wire [0:0] v_9282;
  wire [0:0] v_9283;
  function [0:0] mux_9283(input [0:0] sel);
    case (sel) 0: mux_9283 = 1'h0; 1: mux_9283 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9284;
  wire [0:0] v_9285;
  function [0:0] mux_9285(input [0:0] sel);
    case (sel) 0: mux_9285 = 1'h0; 1: mux_9285 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9286;
  wire [0:0] v_9287;
  wire [0:0] v_9288;
  wire [0:0] v_9289;
  function [0:0] mux_9289(input [0:0] sel);
    case (sel) 0: mux_9289 = 1'h0; 1: mux_9289 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9290;
  function [0:0] mux_9290(input [0:0] sel);
    case (sel) 0: mux_9290 = 1'h0; 1: mux_9290 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9291 = 1'h0;
  wire [0:0] v_9292;
  wire [0:0] v_9293;
  wire [0:0] act_9294;
  wire [0:0] v_9295;
  wire [0:0] v_9296;
  wire [0:0] v_9297;
  reg [0:0] v_9298 = 1'h0;
  wire [0:0] v_9299;
  wire [0:0] v_9300;
  wire [0:0] act_9301;
  wire [0:0] v_9302;
  wire [0:0] v_9303;
  wire [0:0] v_9304;
  wire [0:0] v_9305;
  wire [0:0] v_9306;
  wire [0:0] v_9307;
  function [0:0] mux_9307(input [0:0] sel);
    case (sel) 0: mux_9307 = 1'h0; 1: mux_9307 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9308;
  wire [0:0] v_9309;
  function [0:0] mux_9309(input [0:0] sel);
    case (sel) 0: mux_9309 = 1'h0; 1: mux_9309 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9310;
  wire [0:0] v_9311;
  wire [0:0] v_9312;
  wire [0:0] v_9313;
  function [0:0] mux_9313(input [0:0] sel);
    case (sel) 0: mux_9313 = 1'h0; 1: mux_9313 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9314;
  function [0:0] mux_9314(input [0:0] sel);
    case (sel) 0: mux_9314 = 1'h0; 1: mux_9314 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9315 = 1'h0;
  wire [0:0] v_9316;
  wire [0:0] v_9317;
  wire [0:0] act_9318;
  wire [0:0] v_9319;
  wire [0:0] v_9320;
  wire [0:0] v_9321;
  wire [0:0] v_9322;
  wire [0:0] v_9323;
  wire [0:0] v_9324;
  function [0:0] mux_9324(input [0:0] sel);
    case (sel) 0: mux_9324 = 1'h0; 1: mux_9324 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9325;
  function [0:0] mux_9325(input [0:0] sel);
    case (sel) 0: mux_9325 = 1'h0; 1: mux_9325 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9326;
  wire [0:0] v_9327;
  wire [0:0] v_9328;
  wire [0:0] v_9329;
  function [0:0] mux_9329(input [0:0] sel);
    case (sel) 0: mux_9329 = 1'h0; 1: mux_9329 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9330;
  function [0:0] mux_9330(input [0:0] sel);
    case (sel) 0: mux_9330 = 1'h0; 1: mux_9330 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9331;
  wire [0:0] v_9332;
  wire [0:0] v_9333;
  wire [0:0] v_9334;
  wire [0:0] v_9335;
  wire [0:0] v_9336;
  function [0:0] mux_9336(input [0:0] sel);
    case (sel) 0: mux_9336 = 1'h0; 1: mux_9336 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9337;
  function [0:0] mux_9337(input [0:0] sel);
    case (sel) 0: mux_9337 = 1'h0; 1: mux_9337 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9338;
  wire [0:0] v_9339;
  wire [0:0] v_9340;
  wire [0:0] v_9341;
  function [0:0] mux_9341(input [0:0] sel);
    case (sel) 0: mux_9341 = 1'h0; 1: mux_9341 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9342;
  function [0:0] mux_9342(input [0:0] sel);
    case (sel) 0: mux_9342 = 1'h0; 1: mux_9342 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9343;
  wire [0:0] v_9344;
  wire [0:0] v_9345;
  wire [0:0] v_9346;
  wire [0:0] v_9347;
  wire [0:0] v_9348;
  function [0:0] mux_9348(input [0:0] sel);
    case (sel) 0: mux_9348 = 1'h0; 1: mux_9348 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9349;
  function [0:0] mux_9349(input [0:0] sel);
    case (sel) 0: mux_9349 = 1'h0; 1: mux_9349 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9350;
  wire [0:0] v_9351;
  wire [0:0] v_9352;
  wire [0:0] v_9353;
  function [0:0] mux_9353(input [0:0] sel);
    case (sel) 0: mux_9353 = 1'h0; 1: mux_9353 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9354;
  function [0:0] mux_9354(input [0:0] sel);
    case (sel) 0: mux_9354 = 1'h0; 1: mux_9354 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9355;
  wire [0:0] v_9356;
  wire [0:0] v_9357;
  wire [0:0] v_9358;
  wire [0:0] v_9359;
  wire [0:0] v_9360;
  function [0:0] mux_9360(input [0:0] sel);
    case (sel) 0: mux_9360 = 1'h0; 1: mux_9360 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9361;
  function [0:0] mux_9361(input [0:0] sel);
    case (sel) 0: mux_9361 = 1'h0; 1: mux_9361 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9362;
  wire [0:0] v_9363;
  wire [0:0] v_9364;
  wire [0:0] v_9365;
  function [0:0] mux_9365(input [0:0] sel);
    case (sel) 0: mux_9365 = 1'h0; 1: mux_9365 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9366;
  function [0:0] mux_9366(input [0:0] sel);
    case (sel) 0: mux_9366 = 1'h0; 1: mux_9366 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9367;
  wire [0:0] v_9368;
  wire [0:0] v_9369;
  wire [0:0] v_9370;
  wire [0:0] v_9371;
  wire [0:0] v_9372;
  function [0:0] mux_9372(input [0:0] sel);
    case (sel) 0: mux_9372 = 1'h0; 1: mux_9372 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9373;
  wire [0:0] v_9374;
  function [0:0] mux_9374(input [0:0] sel);
    case (sel) 0: mux_9374 = 1'h0; 1: mux_9374 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9375;
  wire [0:0] v_9376;
  wire [0:0] v_9377;
  wire [0:0] v_9378;
  function [0:0] mux_9378(input [0:0] sel);
    case (sel) 0: mux_9378 = 1'h0; 1: mux_9378 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9379;
  function [0:0] mux_9379(input [0:0] sel);
    case (sel) 0: mux_9379 = 1'h0; 1: mux_9379 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9380 = 1'h0;
  wire [0:0] v_9381;
  wire [0:0] v_9382;
  wire [0:0] act_9383;
  wire [0:0] v_9384;
  wire [0:0] v_9385;
  wire [0:0] v_9386;
  reg [0:0] v_9387 = 1'h0;
  wire [0:0] v_9388;
  wire [0:0] v_9389;
  wire [0:0] act_9390;
  wire [0:0] v_9391;
  wire [0:0] v_9392;
  wire [0:0] v_9393;
  reg [0:0] v_9394 = 1'h0;
  wire [0:0] v_9395;
  wire [0:0] v_9396;
  wire [0:0] act_9397;
  wire [0:0] v_9398;
  wire [0:0] v_9399;
  wire [0:0] v_9400;
  reg [0:0] v_9401 = 1'h0;
  wire [0:0] v_9402;
  wire [0:0] v_9403;
  wire [0:0] act_9404;
  wire [0:0] v_9405;
  wire [0:0] v_9406;
  wire [0:0] v_9407;
  reg [0:0] v_9408 = 1'h0;
  wire [0:0] v_9409;
  wire [0:0] v_9410;
  wire [0:0] act_9411;
  wire [0:0] v_9412;
  wire [0:0] v_9413;
  wire [0:0] v_9414;
  wire [0:0] v_9415;
  wire [0:0] v_9416;
  wire [0:0] v_9417;
  function [0:0] mux_9417(input [0:0] sel);
    case (sel) 0: mux_9417 = 1'h0; 1: mux_9417 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9418;
  wire [0:0] v_9419;
  function [0:0] mux_9419(input [0:0] sel);
    case (sel) 0: mux_9419 = 1'h0; 1: mux_9419 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9420;
  wire [0:0] v_9421;
  wire [0:0] v_9422;
  wire [0:0] v_9423;
  function [0:0] mux_9423(input [0:0] sel);
    case (sel) 0: mux_9423 = 1'h0; 1: mux_9423 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9424;
  function [0:0] mux_9424(input [0:0] sel);
    case (sel) 0: mux_9424 = 1'h0; 1: mux_9424 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9425 = 1'h0;
  wire [0:0] v_9426;
  wire [0:0] v_9427;
  wire [0:0] act_9428;
  wire [0:0] v_9429;
  wire [0:0] v_9430;
  wire [0:0] v_9431;
  wire [0:0] v_9432;
  wire [0:0] v_9433;
  wire [0:0] v_9434;
  function [0:0] mux_9434(input [0:0] sel);
    case (sel) 0: mux_9434 = 1'h0; 1: mux_9434 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9435;
  function [0:0] mux_9435(input [0:0] sel);
    case (sel) 0: mux_9435 = 1'h0; 1: mux_9435 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9436;
  wire [0:0] v_9437;
  wire [0:0] v_9438;
  wire [0:0] v_9439;
  function [0:0] mux_9439(input [0:0] sel);
    case (sel) 0: mux_9439 = 1'h0; 1: mux_9439 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9440;
  function [0:0] mux_9440(input [0:0] sel);
    case (sel) 0: mux_9440 = 1'h0; 1: mux_9440 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9441;
  wire [0:0] v_9442;
  wire [0:0] v_9443;
  wire [0:0] v_9444;
  wire [0:0] v_9445;
  wire [0:0] v_9446;
  function [0:0] mux_9446(input [0:0] sel);
    case (sel) 0: mux_9446 = 1'h0; 1: mux_9446 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9447;
  wire [0:0] v_9448;
  function [0:0] mux_9448(input [0:0] sel);
    case (sel) 0: mux_9448 = 1'h0; 1: mux_9448 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9449;
  wire [0:0] v_9450;
  wire [0:0] v_9451;
  wire [0:0] v_9452;
  function [0:0] mux_9452(input [0:0] sel);
    case (sel) 0: mux_9452 = 1'h0; 1: mux_9452 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9453;
  function [0:0] mux_9453(input [0:0] sel);
    case (sel) 0: mux_9453 = 1'h0; 1: mux_9453 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9454 = 1'h0;
  wire [0:0] v_9455;
  wire [0:0] v_9456;
  wire [0:0] act_9457;
  wire [0:0] v_9458;
  wire [0:0] v_9459;
  wire [0:0] v_9460;
  reg [0:0] v_9461 = 1'h0;
  wire [0:0] v_9462;
  wire [0:0] v_9463;
  wire [0:0] act_9464;
  wire [0:0] v_9465;
  wire [0:0] v_9466;
  wire [0:0] v_9467;
  wire [0:0] v_9468;
  wire [0:0] v_9469;
  wire [0:0] v_9470;
  function [0:0] mux_9470(input [0:0] sel);
    case (sel) 0: mux_9470 = 1'h0; 1: mux_9470 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9471;
  wire [0:0] v_9472;
  function [0:0] mux_9472(input [0:0] sel);
    case (sel) 0: mux_9472 = 1'h0; 1: mux_9472 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9473;
  wire [0:0] v_9474;
  wire [0:0] v_9475;
  wire [0:0] v_9476;
  function [0:0] mux_9476(input [0:0] sel);
    case (sel) 0: mux_9476 = 1'h0; 1: mux_9476 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9477;
  function [0:0] mux_9477(input [0:0] sel);
    case (sel) 0: mux_9477 = 1'h0; 1: mux_9477 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9478 = 1'h0;
  wire [0:0] v_9479;
  wire [0:0] v_9480;
  wire [0:0] act_9481;
  wire [0:0] v_9482;
  wire [0:0] v_9483;
  wire [0:0] v_9484;
  wire [0:0] v_9485;
  wire [0:0] v_9486;
  wire [0:0] v_9487;
  function [0:0] mux_9487(input [0:0] sel);
    case (sel) 0: mux_9487 = 1'h0; 1: mux_9487 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9488;
  function [0:0] mux_9488(input [0:0] sel);
    case (sel) 0: mux_9488 = 1'h0; 1: mux_9488 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9489;
  wire [0:0] v_9490;
  wire [0:0] v_9491;
  wire [0:0] v_9492;
  function [0:0] mux_9492(input [0:0] sel);
    case (sel) 0: mux_9492 = 1'h0; 1: mux_9492 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9493;
  function [0:0] mux_9493(input [0:0] sel);
    case (sel) 0: mux_9493 = 1'h0; 1: mux_9493 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9494;
  wire [0:0] v_9495;
  wire [0:0] v_9496;
  wire [0:0] v_9497;
  wire [0:0] v_9498;
  wire [0:0] v_9499;
  function [0:0] mux_9499(input [0:0] sel);
    case (sel) 0: mux_9499 = 1'h0; 1: mux_9499 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9500;
  function [0:0] mux_9500(input [0:0] sel);
    case (sel) 0: mux_9500 = 1'h0; 1: mux_9500 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9501;
  wire [0:0] v_9502;
  wire [0:0] v_9503;
  wire [0:0] v_9504;
  function [0:0] mux_9504(input [0:0] sel);
    case (sel) 0: mux_9504 = 1'h0; 1: mux_9504 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9505;
  function [0:0] mux_9505(input [0:0] sel);
    case (sel) 0: mux_9505 = 1'h0; 1: mux_9505 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9506;
  wire [0:0] v_9507;
  wire [0:0] v_9508;
  wire [0:0] v_9509;
  wire [0:0] v_9510;
  wire [0:0] v_9511;
  function [0:0] mux_9511(input [0:0] sel);
    case (sel) 0: mux_9511 = 1'h0; 1: mux_9511 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9512;
  wire [0:0] v_9513;
  function [0:0] mux_9513(input [0:0] sel);
    case (sel) 0: mux_9513 = 1'h0; 1: mux_9513 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9514;
  wire [0:0] v_9515;
  wire [0:0] v_9516;
  wire [0:0] v_9517;
  function [0:0] mux_9517(input [0:0] sel);
    case (sel) 0: mux_9517 = 1'h0; 1: mux_9517 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9518;
  function [0:0] mux_9518(input [0:0] sel);
    case (sel) 0: mux_9518 = 1'h0; 1: mux_9518 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9519 = 1'h0;
  wire [0:0] v_9520;
  wire [0:0] v_9521;
  wire [0:0] act_9522;
  wire [0:0] v_9523;
  wire [0:0] v_9524;
  wire [0:0] v_9525;
  reg [0:0] v_9526 = 1'h0;
  wire [0:0] v_9527;
  wire [0:0] v_9528;
  wire [0:0] act_9529;
  wire [0:0] v_9530;
  wire [0:0] v_9531;
  wire [0:0] v_9532;
  reg [0:0] v_9533 = 1'h0;
  wire [0:0] v_9534;
  wire [0:0] v_9535;
  wire [0:0] act_9536;
  wire [0:0] v_9537;
  wire [0:0] v_9538;
  wire [0:0] v_9539;
  wire [0:0] v_9540;
  wire [0:0] v_9541;
  wire [0:0] v_9542;
  function [0:0] mux_9542(input [0:0] sel);
    case (sel) 0: mux_9542 = 1'h0; 1: mux_9542 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9543;
  wire [0:0] v_9544;
  function [0:0] mux_9544(input [0:0] sel);
    case (sel) 0: mux_9544 = 1'h0; 1: mux_9544 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9545;
  wire [0:0] v_9546;
  wire [0:0] v_9547;
  wire [0:0] v_9548;
  function [0:0] mux_9548(input [0:0] sel);
    case (sel) 0: mux_9548 = 1'h0; 1: mux_9548 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9549;
  function [0:0] mux_9549(input [0:0] sel);
    case (sel) 0: mux_9549 = 1'h0; 1: mux_9549 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9550 = 1'h0;
  wire [0:0] v_9551;
  wire [0:0] v_9552;
  wire [0:0] act_9553;
  wire [0:0] v_9554;
  wire [0:0] v_9555;
  wire [0:0] v_9556;
  wire [0:0] v_9557;
  wire [0:0] v_9558;
  wire [0:0] v_9559;
  function [0:0] mux_9559(input [0:0] sel);
    case (sel) 0: mux_9559 = 1'h0; 1: mux_9559 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9560;
  function [0:0] mux_9560(input [0:0] sel);
    case (sel) 0: mux_9560 = 1'h0; 1: mux_9560 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9561;
  wire [0:0] v_9562;
  wire [0:0] v_9563;
  wire [0:0] v_9564;
  function [0:0] mux_9564(input [0:0] sel);
    case (sel) 0: mux_9564 = 1'h0; 1: mux_9564 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9565;
  function [0:0] mux_9565(input [0:0] sel);
    case (sel) 0: mux_9565 = 1'h0; 1: mux_9565 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9566;
  wire [0:0] v_9567;
  wire [0:0] v_9568;
  wire [0:0] v_9569;
  wire [0:0] v_9570;
  wire [0:0] v_9571;
  function [0:0] mux_9571(input [0:0] sel);
    case (sel) 0: mux_9571 = 1'h0; 1: mux_9571 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9572;
  wire [0:0] v_9573;
  function [0:0] mux_9573(input [0:0] sel);
    case (sel) 0: mux_9573 = 1'h0; 1: mux_9573 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9574;
  wire [0:0] v_9575;
  wire [0:0] v_9576;
  wire [0:0] v_9577;
  function [0:0] mux_9577(input [0:0] sel);
    case (sel) 0: mux_9577 = 1'h0; 1: mux_9577 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9578;
  function [0:0] mux_9578(input [0:0] sel);
    case (sel) 0: mux_9578 = 1'h0; 1: mux_9578 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9579 = 1'h0;
  wire [0:0] v_9580;
  wire [0:0] v_9581;
  wire [0:0] act_9582;
  wire [0:0] v_9583;
  wire [0:0] v_9584;
  wire [0:0] v_9585;
  reg [0:0] v_9586 = 1'h0;
  wire [0:0] v_9587;
  wire [0:0] v_9588;
  wire [0:0] act_9589;
  wire [0:0] v_9590;
  wire [0:0] v_9591;
  wire [0:0] v_9592;
  wire [0:0] v_9593;
  wire [0:0] v_9594;
  wire [0:0] v_9595;
  function [0:0] mux_9595(input [0:0] sel);
    case (sel) 0: mux_9595 = 1'h0; 1: mux_9595 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9596;
  wire [0:0] v_9597;
  function [0:0] mux_9597(input [0:0] sel);
    case (sel) 0: mux_9597 = 1'h0; 1: mux_9597 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9598;
  wire [0:0] v_9599;
  wire [0:0] v_9600;
  wire [0:0] v_9601;
  function [0:0] mux_9601(input [0:0] sel);
    case (sel) 0: mux_9601 = 1'h0; 1: mux_9601 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9602;
  function [0:0] mux_9602(input [0:0] sel);
    case (sel) 0: mux_9602 = 1'h0; 1: mux_9602 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9603 = 1'h0;
  wire [0:0] v_9604;
  wire [0:0] v_9605;
  wire [0:0] act_9606;
  wire [0:0] v_9607;
  wire [0:0] v_9608;
  wire [0:0] v_9609;
  wire [0:0] v_9610;
  wire [0:0] v_9611;
  wire [0:0] v_9612;
  function [0:0] mux_9612(input [0:0] sel);
    case (sel) 0: mux_9612 = 1'h0; 1: mux_9612 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9613;
  function [0:0] mux_9613(input [0:0] sel);
    case (sel) 0: mux_9613 = 1'h0; 1: mux_9613 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9614;
  wire [0:0] v_9615;
  wire [0:0] v_9616;
  wire [0:0] v_9617;
  function [0:0] mux_9617(input [0:0] sel);
    case (sel) 0: mux_9617 = 1'h0; 1: mux_9617 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9618;
  function [0:0] mux_9618(input [0:0] sel);
    case (sel) 0: mux_9618 = 1'h0; 1: mux_9618 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9619;
  wire [0:0] v_9620;
  wire [0:0] v_9621;
  wire [0:0] v_9622;
  wire [0:0] v_9623;
  wire [0:0] v_9624;
  function [0:0] mux_9624(input [0:0] sel);
    case (sel) 0: mux_9624 = 1'h0; 1: mux_9624 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9625;
  function [0:0] mux_9625(input [0:0] sel);
    case (sel) 0: mux_9625 = 1'h0; 1: mux_9625 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9626;
  wire [0:0] v_9627;
  wire [0:0] v_9628;
  wire [0:0] v_9629;
  function [0:0] mux_9629(input [0:0] sel);
    case (sel) 0: mux_9629 = 1'h0; 1: mux_9629 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9630;
  function [0:0] mux_9630(input [0:0] sel);
    case (sel) 0: mux_9630 = 1'h0; 1: mux_9630 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9631;
  wire [0:0] v_9632;
  wire [0:0] v_9633;
  wire [0:0] v_9634;
  wire [0:0] v_9635;
  wire [0:0] v_9636;
  function [0:0] mux_9636(input [0:0] sel);
    case (sel) 0: mux_9636 = 1'h0; 1: mux_9636 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9637;
  function [0:0] mux_9637(input [0:0] sel);
    case (sel) 0: mux_9637 = 1'h0; 1: mux_9637 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9638;
  wire [0:0] v_9639;
  wire [0:0] v_9640;
  wire [0:0] v_9641;
  function [0:0] mux_9641(input [0:0] sel);
    case (sel) 0: mux_9641 = 1'h0; 1: mux_9641 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9642;
  function [0:0] mux_9642(input [0:0] sel);
    case (sel) 0: mux_9642 = 1'h0; 1: mux_9642 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9643;
  wire [0:0] v_9644;
  wire [0:0] v_9645;
  wire [0:0] v_9646;
  wire [0:0] v_9647;
  wire [0:0] v_9648;
  function [0:0] mux_9648(input [0:0] sel);
    case (sel) 0: mux_9648 = 1'h0; 1: mux_9648 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9649;
  wire [0:0] v_9650;
  function [0:0] mux_9650(input [0:0] sel);
    case (sel) 0: mux_9650 = 1'h0; 1: mux_9650 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9651;
  wire [0:0] v_9652;
  wire [0:0] v_9653;
  wire [0:0] v_9654;
  function [0:0] mux_9654(input [0:0] sel);
    case (sel) 0: mux_9654 = 1'h0; 1: mux_9654 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9655;
  function [0:0] mux_9655(input [0:0] sel);
    case (sel) 0: mux_9655 = 1'h0; 1: mux_9655 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9656 = 1'h0;
  wire [0:0] v_9657;
  wire [0:0] v_9658;
  wire [0:0] act_9659;
  wire [0:0] v_9660;
  wire [0:0] v_9661;
  wire [0:0] v_9662;
  reg [0:0] v_9663 = 1'h0;
  wire [0:0] v_9664;
  wire [0:0] v_9665;
  wire [0:0] act_9666;
  wire [0:0] v_9667;
  wire [0:0] v_9668;
  wire [0:0] v_9669;
  reg [0:0] v_9670 = 1'h0;
  wire [0:0] v_9671;
  wire [0:0] v_9672;
  wire [0:0] act_9673;
  wire [0:0] v_9674;
  wire [0:0] v_9675;
  wire [0:0] v_9676;
  reg [0:0] v_9677 = 1'h0;
  wire [0:0] v_9678;
  wire [0:0] v_9679;
  wire [0:0] act_9680;
  wire [0:0] v_9681;
  wire [0:0] v_9682;
  wire [0:0] v_9683;
  wire [0:0] v_9684;
  wire [0:0] v_9685;
  wire [0:0] v_9686;
  function [0:0] mux_9686(input [0:0] sel);
    case (sel) 0: mux_9686 = 1'h0; 1: mux_9686 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9687;
  wire [0:0] v_9688;
  function [0:0] mux_9688(input [0:0] sel);
    case (sel) 0: mux_9688 = 1'h0; 1: mux_9688 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9689;
  wire [0:0] v_9690;
  wire [0:0] v_9691;
  wire [0:0] v_9692;
  function [0:0] mux_9692(input [0:0] sel);
    case (sel) 0: mux_9692 = 1'h0; 1: mux_9692 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9693;
  function [0:0] mux_9693(input [0:0] sel);
    case (sel) 0: mux_9693 = 1'h0; 1: mux_9693 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9694 = 1'h0;
  wire [0:0] v_9695;
  wire [0:0] v_9696;
  wire [0:0] act_9697;
  wire [0:0] v_9698;
  wire [0:0] v_9699;
  wire [0:0] v_9700;
  wire [0:0] v_9701;
  wire [0:0] v_9702;
  wire [0:0] v_9703;
  function [0:0] mux_9703(input [0:0] sel);
    case (sel) 0: mux_9703 = 1'h0; 1: mux_9703 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9704;
  function [0:0] mux_9704(input [0:0] sel);
    case (sel) 0: mux_9704 = 1'h0; 1: mux_9704 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9705;
  wire [0:0] v_9706;
  wire [0:0] v_9707;
  wire [0:0] v_9708;
  function [0:0] mux_9708(input [0:0] sel);
    case (sel) 0: mux_9708 = 1'h0; 1: mux_9708 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9709;
  function [0:0] mux_9709(input [0:0] sel);
    case (sel) 0: mux_9709 = 1'h0; 1: mux_9709 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9710;
  wire [0:0] v_9711;
  wire [0:0] v_9712;
  wire [0:0] v_9713;
  wire [0:0] v_9714;
  wire [0:0] v_9715;
  function [0:0] mux_9715(input [0:0] sel);
    case (sel) 0: mux_9715 = 1'h0; 1: mux_9715 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9716;
  wire [0:0] v_9717;
  function [0:0] mux_9717(input [0:0] sel);
    case (sel) 0: mux_9717 = 1'h0; 1: mux_9717 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9718;
  wire [0:0] v_9719;
  wire [0:0] v_9720;
  wire [0:0] v_9721;
  function [0:0] mux_9721(input [0:0] sel);
    case (sel) 0: mux_9721 = 1'h0; 1: mux_9721 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9722;
  function [0:0] mux_9722(input [0:0] sel);
    case (sel) 0: mux_9722 = 1'h0; 1: mux_9722 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9723 = 1'h0;
  wire [0:0] v_9724;
  wire [0:0] v_9725;
  wire [0:0] act_9726;
  wire [0:0] v_9727;
  wire [0:0] v_9728;
  wire [0:0] v_9729;
  reg [0:0] v_9730 = 1'h0;
  wire [0:0] v_9731;
  wire [0:0] v_9732;
  wire [0:0] act_9733;
  wire [0:0] v_9734;
  wire [0:0] v_9735;
  wire [0:0] v_9736;
  wire [0:0] v_9737;
  wire [0:0] v_9738;
  wire [0:0] v_9739;
  function [0:0] mux_9739(input [0:0] sel);
    case (sel) 0: mux_9739 = 1'h0; 1: mux_9739 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9740;
  wire [0:0] v_9741;
  function [0:0] mux_9741(input [0:0] sel);
    case (sel) 0: mux_9741 = 1'h0; 1: mux_9741 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9742;
  wire [0:0] v_9743;
  wire [0:0] v_9744;
  wire [0:0] v_9745;
  function [0:0] mux_9745(input [0:0] sel);
    case (sel) 0: mux_9745 = 1'h0; 1: mux_9745 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9746;
  function [0:0] mux_9746(input [0:0] sel);
    case (sel) 0: mux_9746 = 1'h0; 1: mux_9746 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9747 = 1'h0;
  wire [0:0] v_9748;
  wire [0:0] v_9749;
  wire [0:0] act_9750;
  wire [0:0] v_9751;
  wire [0:0] v_9752;
  wire [0:0] v_9753;
  wire [0:0] v_9754;
  wire [0:0] v_9755;
  wire [0:0] v_9756;
  function [0:0] mux_9756(input [0:0] sel);
    case (sel) 0: mux_9756 = 1'h0; 1: mux_9756 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9757;
  function [0:0] mux_9757(input [0:0] sel);
    case (sel) 0: mux_9757 = 1'h0; 1: mux_9757 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9758;
  wire [0:0] v_9759;
  wire [0:0] v_9760;
  wire [0:0] v_9761;
  function [0:0] mux_9761(input [0:0] sel);
    case (sel) 0: mux_9761 = 1'h0; 1: mux_9761 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9762;
  function [0:0] mux_9762(input [0:0] sel);
    case (sel) 0: mux_9762 = 1'h0; 1: mux_9762 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9763;
  wire [0:0] v_9764;
  wire [0:0] v_9765;
  wire [0:0] v_9766;
  wire [0:0] v_9767;
  wire [0:0] v_9768;
  function [0:0] mux_9768(input [0:0] sel);
    case (sel) 0: mux_9768 = 1'h0; 1: mux_9768 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9769;
  function [0:0] mux_9769(input [0:0] sel);
    case (sel) 0: mux_9769 = 1'h0; 1: mux_9769 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9770;
  wire [0:0] v_9771;
  wire [0:0] v_9772;
  wire [0:0] v_9773;
  function [0:0] mux_9773(input [0:0] sel);
    case (sel) 0: mux_9773 = 1'h0; 1: mux_9773 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9774;
  function [0:0] mux_9774(input [0:0] sel);
    case (sel) 0: mux_9774 = 1'h0; 1: mux_9774 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9775;
  wire [0:0] v_9776;
  wire [0:0] v_9777;
  wire [0:0] v_9778;
  wire [0:0] v_9779;
  wire [0:0] v_9780;
  function [0:0] mux_9780(input [0:0] sel);
    case (sel) 0: mux_9780 = 1'h0; 1: mux_9780 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9781;
  wire [0:0] v_9782;
  function [0:0] mux_9782(input [0:0] sel);
    case (sel) 0: mux_9782 = 1'h0; 1: mux_9782 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9783;
  wire [0:0] v_9784;
  wire [0:0] v_9785;
  wire [0:0] v_9786;
  function [0:0] mux_9786(input [0:0] sel);
    case (sel) 0: mux_9786 = 1'h0; 1: mux_9786 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9787;
  function [0:0] mux_9787(input [0:0] sel);
    case (sel) 0: mux_9787 = 1'h0; 1: mux_9787 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9788 = 1'h0;
  wire [0:0] v_9789;
  wire [0:0] v_9790;
  wire [0:0] act_9791;
  wire [0:0] v_9792;
  wire [0:0] v_9793;
  wire [0:0] v_9794;
  reg [0:0] v_9795 = 1'h0;
  wire [0:0] v_9796;
  wire [0:0] v_9797;
  wire [0:0] act_9798;
  wire [0:0] v_9799;
  wire [0:0] v_9800;
  wire [0:0] v_9801;
  reg [0:0] v_9802 = 1'h0;
  wire [0:0] v_9803;
  wire [0:0] v_9804;
  wire [0:0] act_9805;
  wire [0:0] v_9806;
  wire [0:0] v_9807;
  wire [0:0] v_9808;
  wire [0:0] v_9809;
  wire [0:0] v_9810;
  wire [0:0] v_9811;
  function [0:0] mux_9811(input [0:0] sel);
    case (sel) 0: mux_9811 = 1'h0; 1: mux_9811 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9812;
  wire [0:0] v_9813;
  function [0:0] mux_9813(input [0:0] sel);
    case (sel) 0: mux_9813 = 1'h0; 1: mux_9813 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9814;
  wire [0:0] v_9815;
  wire [0:0] v_9816;
  wire [0:0] v_9817;
  function [0:0] mux_9817(input [0:0] sel);
    case (sel) 0: mux_9817 = 1'h0; 1: mux_9817 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9818;
  function [0:0] mux_9818(input [0:0] sel);
    case (sel) 0: mux_9818 = 1'h0; 1: mux_9818 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9819 = 1'h0;
  wire [0:0] v_9820;
  wire [0:0] v_9821;
  wire [0:0] act_9822;
  wire [0:0] v_9823;
  wire [0:0] v_9824;
  wire [0:0] v_9825;
  wire [0:0] v_9826;
  wire [0:0] v_9827;
  wire [0:0] v_9828;
  function [0:0] mux_9828(input [0:0] sel);
    case (sel) 0: mux_9828 = 1'h0; 1: mux_9828 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9829;
  function [0:0] mux_9829(input [0:0] sel);
    case (sel) 0: mux_9829 = 1'h0; 1: mux_9829 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9830;
  wire [0:0] v_9831;
  wire [0:0] v_9832;
  wire [0:0] v_9833;
  function [0:0] mux_9833(input [0:0] sel);
    case (sel) 0: mux_9833 = 1'h0; 1: mux_9833 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9834;
  function [0:0] mux_9834(input [0:0] sel);
    case (sel) 0: mux_9834 = 1'h0; 1: mux_9834 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9835;
  wire [0:0] v_9836;
  wire [0:0] v_9837;
  wire [0:0] v_9838;
  wire [0:0] v_9839;
  wire [0:0] v_9840;
  function [0:0] mux_9840(input [0:0] sel);
    case (sel) 0: mux_9840 = 1'h0; 1: mux_9840 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9841;
  wire [0:0] v_9842;
  function [0:0] mux_9842(input [0:0] sel);
    case (sel) 0: mux_9842 = 1'h0; 1: mux_9842 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9843;
  wire [0:0] v_9844;
  wire [0:0] v_9845;
  wire [0:0] v_9846;
  function [0:0] mux_9846(input [0:0] sel);
    case (sel) 0: mux_9846 = 1'h0; 1: mux_9846 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9847;
  function [0:0] mux_9847(input [0:0] sel);
    case (sel) 0: mux_9847 = 1'h0; 1: mux_9847 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9848 = 1'h0;
  wire [0:0] v_9849;
  wire [0:0] v_9850;
  wire [0:0] act_9851;
  wire [0:0] v_9852;
  wire [0:0] v_9853;
  wire [0:0] v_9854;
  reg [0:0] v_9855 = 1'h0;
  wire [0:0] v_9856;
  wire [0:0] v_9857;
  wire [0:0] act_9858;
  wire [0:0] v_9859;
  wire [0:0] v_9860;
  wire [0:0] v_9861;
  wire [0:0] v_9862;
  wire [0:0] v_9863;
  wire [0:0] v_9864;
  function [0:0] mux_9864(input [0:0] sel);
    case (sel) 0: mux_9864 = 1'h0; 1: mux_9864 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9865;
  wire [0:0] v_9866;
  function [0:0] mux_9866(input [0:0] sel);
    case (sel) 0: mux_9866 = 1'h0; 1: mux_9866 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9867;
  wire [0:0] v_9868;
  wire [0:0] v_9869;
  wire [0:0] v_9870;
  function [0:0] mux_9870(input [0:0] sel);
    case (sel) 0: mux_9870 = 1'h0; 1: mux_9870 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9871;
  function [0:0] mux_9871(input [0:0] sel);
    case (sel) 0: mux_9871 = 1'h0; 1: mux_9871 = 1'h0;
    endcase
  endfunction
  reg [0:0] v_9872 = 1'h0;
  wire [0:0] v_9873;
  wire [0:0] v_9874;
  wire [0:0] act_9875;
  wire [0:0] v_9876;
  wire [0:0] v_9877;
  wire [0:0] v_9878;
  wire [0:0] v_9879;
  wire [0:0] v_9880;
  wire [0:0] v_9881;
  function [0:0] mux_9881(input [0:0] sel);
    case (sel) 0: mux_9881 = 1'h0; 1: mux_9881 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9882;
  function [0:0] mux_9882(input [0:0] sel);
    case (sel) 0: mux_9882 = 1'h0; 1: mux_9882 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9883;
  wire [0:0] v_9884;
  wire [0:0] v_9885;
  wire [0:0] v_9886;
  function [0:0] mux_9886(input [0:0] sel);
    case (sel) 0: mux_9886 = 1'h0; 1: mux_9886 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9887;
  function [0:0] mux_9887(input [0:0] sel);
    case (sel) 0: mux_9887 = 1'h0; 1: mux_9887 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9888;
  wire [0:0] v_9889;
  wire [0:0] v_9890;
  wire [0:0] v_9891;
  wire [0:0] v_9892;
  wire [0:0] v_9893;
  function [0:0] mux_9893(input [0:0] sel);
    case (sel) 0: mux_9893 = 1'h0; 1: mux_9893 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9894;
  function [0:0] mux_9894(input [0:0] sel);
    case (sel) 0: mux_9894 = 1'h0; 1: mux_9894 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9895;
  wire [0:0] v_9896;
  wire [0:0] v_9897;
  wire [0:0] v_9898;
  function [0:0] mux_9898(input [0:0] sel);
    case (sel) 0: mux_9898 = 1'h0; 1: mux_9898 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9899;
  function [0:0] mux_9899(input [0:0] sel);
    case (sel) 0: mux_9899 = 1'h0; 1: mux_9899 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9900;
  wire [0:0] v_9901;
  wire [0:0] v_9902;
  wire [0:0] v_9903;
  wire [0:0] v_9904;
  wire [0:0] v_9905;
  function [0:0] mux_9905(input [0:0] sel);
    case (sel) 0: mux_9905 = 1'h0; 1: mux_9905 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9906;
  function [0:0] mux_9906(input [0:0] sel);
    case (sel) 0: mux_9906 = 1'h0; 1: mux_9906 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9907;
  wire [0:0] v_9908;
  wire [0:0] v_9909;
  wire [0:0] v_9910;
  function [0:0] mux_9910(input [0:0] sel);
    case (sel) 0: mux_9910 = 1'h0; 1: mux_9910 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9911;
  function [0:0] mux_9911(input [0:0] sel);
    case (sel) 0: mux_9911 = 1'h0; 1: mux_9911 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9912;
  wire [0:0] v_9913;
  wire [0:0] v_9914;
  wire [0:0] v_9915;
  wire [0:0] v_9916;
  wire [0:0] v_9917;
  function [0:0] mux_9917(input [0:0] sel);
    case (sel) 0: mux_9917 = 1'h0; 1: mux_9917 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9918;
  function [0:0] mux_9918(input [0:0] sel);
    case (sel) 0: mux_9918 = 1'h0; 1: mux_9918 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9919;
  wire [0:0] v_9920;
  wire [0:0] v_9921;
  wire [0:0] v_9922;
  function [0:0] mux_9922(input [0:0] sel);
    case (sel) 0: mux_9922 = 1'h0; 1: mux_9922 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9923;
  function [0:0] mux_9923(input [0:0] sel);
    case (sel) 0: mux_9923 = 1'h0; 1: mux_9923 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9924;
  wire [0:0] v_9925;
  wire [0:0] v_9926;
  wire [0:0] v_9927;
  wire [0:0] v_9928;
  wire [0:0] v_9929;
  function [0:0] mux_9929(input [0:0] sel);
    case (sel) 0: mux_9929 = 1'h0; 1: mux_9929 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9930;
  function [0:0] mux_9930(input [0:0] sel);
    case (sel) 0: mux_9930 = 1'h0; 1: mux_9930 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9931;
  wire [0:0] v_9932;
  wire [0:0] v_9933;
  wire [0:0] v_9934;
  function [0:0] mux_9934(input [0:0] sel);
    case (sel) 0: mux_9934 = 1'h0; 1: mux_9934 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9935;
  function [0:0] mux_9935(input [0:0] sel);
    case (sel) 0: mux_9935 = 1'h0; 1: mux_9935 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9936;
  wire [0:0] v_9937;
  wire [0:0] v_9938;
  wire [0:0] v_9939;
  wire [0:0] v_9940;
  wire [0:0] v_9941;
  function [0:0] mux_9941(input [0:0] sel);
    case (sel) 0: mux_9941 = 1'h0; 1: mux_9941 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9942;
  function [0:0] mux_9942(input [0:0] sel);
    case (sel) 0: mux_9942 = 1'h0; 1: mux_9942 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9943;
  wire [0:0] v_9944;
  wire [0:0] v_9945;
  wire [0:0] v_9946;
  function [0:0] mux_9946(input [0:0] sel);
    case (sel) 0: mux_9946 = 1'h0; 1: mux_9946 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9947;
  function [0:0] mux_9947(input [0:0] sel);
    case (sel) 0: mux_9947 = 1'h0; 1: mux_9947 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9948;
  wire [0:0] v_9949;
  wire [0:0] v_9950;
  wire [0:0] v_9951;
  wire [0:0] v_9952;
  wire [0:0] v_9953;
  function [0:0] mux_9953(input [0:0] sel);
    case (sel) 0: mux_9953 = 1'h0; 1: mux_9953 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9954;
  function [0:0] mux_9954(input [0:0] sel);
    case (sel) 0: mux_9954 = 1'h0; 1: mux_9954 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9955;
  wire [0:0] v_9956;
  wire [0:0] v_9957;
  wire [0:0] v_9958;
  function [0:0] mux_9958(input [0:0] sel);
    case (sel) 0: mux_9958 = 1'h0; 1: mux_9958 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9959;
  function [0:0] mux_9959(input [0:0] sel);
    case (sel) 0: mux_9959 = 1'h0; 1: mux_9959 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9960;
  wire [0:0] v_9961;
  wire [0:0] v_9962;
  wire [0:0] v_9963;
  wire [0:0] v_9964;
  wire [0:0] v_9965;
  function [0:0] mux_9965(input [0:0] sel);
    case (sel) 0: mux_9965 = 1'h0; 1: mux_9965 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9966;
  function [0:0] mux_9966(input [0:0] sel);
    case (sel) 0: mux_9966 = 1'h0; 1: mux_9966 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9967;
  wire [0:0] v_9968;
  wire [0:0] v_9969;
  wire [0:0] v_9970;
  function [0:0] mux_9970(input [0:0] sel);
    case (sel) 0: mux_9970 = 1'h0; 1: mux_9970 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9971;
  function [0:0] mux_9971(input [0:0] sel);
    case (sel) 0: mux_9971 = 1'h0; 1: mux_9971 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9972;
  wire [0:0] v_9973;
  wire [0:0] v_9974;
  wire [0:0] v_9975;
  wire [0:0] v_9976;
  wire [0:0] v_9977;
  function [0:0] mux_9977(input [0:0] sel);
    case (sel) 0: mux_9977 = 1'h0; 1: mux_9977 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9978;
  wire [0:0] v_9979;
  wire [0:0] v_9980;
  function [0:0] mux_9980(input [0:0] sel);
    case (sel) 0: mux_9980 = 1'h0; 1: mux_9980 = 1'h0;
    endcase
  endfunction
  wire [0:0] v_9981;
  wire [0:0] v_9982;
  wire [0:0] v_9983;
  wire [0:0] v_9984;
  function [0:0] mux_9984(input [0:0] sel);
    case (sel) 0: mux_9984 = 1'h0; 1: mux_9984 = 1'h1;
    endcase
  endfunction
  wire [0:0] v_9985;
  function [0:0] mux_9985(input [0:0] sel);
    case (sel) 0: mux_9985 = 1'h0; 1: mux_9985 = 1'h0;
    endcase
  endfunction
  reg [7:0] v_9987 = 8'h0;
  wire [7:0] v_9988;
  wire [7:0] v_9989;
  function [7:0] mux_9989(input [0:0] sel);
    case (sel) 0: mux_9989 = 8'h0; 1: mux_9989 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_9990;
  wire [7:0] v_9991;
  wire [7:0] v_9992;
  function [7:0] mux_9992(input [0:0] sel);
    case (sel) 0: mux_9992 = 8'h0; 1: mux_9992 = v_9993;
    endcase
  endfunction
  reg [7:0] v_9993 = 8'h0;
  wire [7:0] v_9994;
  wire [7:0] v_9995;
  function [7:0] mux_9995(input [0:0] sel);
    case (sel) 0: mux_9995 = 8'h0; 1: mux_9995 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_9996;
  wire [7:0] v_9997;
  wire [7:0] v_9998;
  function [7:0] mux_9998(input [0:0] sel);
    case (sel) 0: mux_9998 = 8'h0; 1: mux_9998 = v_9999;
    endcase
  endfunction
  reg [7:0] v_9999 = 8'h0;
  wire [7:0] v_10000;
  wire [7:0] v_10001;
  function [7:0] mux_10001(input [0:0] sel);
    case (sel) 0: mux_10001 = 8'h0; 1: mux_10001 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10002;
  wire [7:0] v_10003;
  wire [7:0] v_10004;
  function [7:0] mux_10004(input [0:0] sel);
    case (sel) 0: mux_10004 = 8'h0; 1: mux_10004 = v_10005;
    endcase
  endfunction
  reg [7:0] v_10005 = 8'h0;
  wire [7:0] v_10006;
  wire [7:0] v_10007;
  function [7:0] mux_10007(input [0:0] sel);
    case (sel) 0: mux_10007 = 8'h0; 1: mux_10007 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10008;
  wire [7:0] v_10009;
  wire [7:0] v_10010;
  function [7:0] mux_10010(input [0:0] sel);
    case (sel) 0: mux_10010 = 8'h0; 1: mux_10010 = v_10011;
    endcase
  endfunction
  reg [7:0] v_10011 = 8'h0;
  wire [7:0] v_10012;
  wire [7:0] v_10013;
  function [7:0] mux_10013(input [0:0] sel);
    case (sel) 0: mux_10013 = 8'h0; 1: mux_10013 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10014;
  wire [7:0] v_10015;
  wire [7:0] v_10016;
  function [7:0] mux_10016(input [0:0] sel);
    case (sel) 0: mux_10016 = 8'h0; 1: mux_10016 = v_10017;
    endcase
  endfunction
  reg [7:0] v_10017 = 8'h0;
  wire [7:0] v_10018;
  wire [7:0] v_10019;
  function [7:0] mux_10019(input [0:0] sel);
    case (sel) 0: mux_10019 = 8'h0; 1: mux_10019 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10020;
  wire [7:0] v_10021;
  wire [7:0] v_10022;
  function [7:0] mux_10022(input [0:0] sel);
    case (sel) 0: mux_10022 = 8'h0; 1: mux_10022 = v_10023;
    endcase
  endfunction
  reg [7:0] v_10023 = 8'h0;
  wire [7:0] v_10024;
  wire [7:0] v_10025;
  function [7:0] mux_10025(input [0:0] sel);
    case (sel) 0: mux_10025 = 8'h0; 1: mux_10025 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10026;
  wire [7:0] v_10027;
  wire [7:0] v_10028;
  function [7:0] mux_10028(input [0:0] sel);
    case (sel) 0: mux_10028 = 8'h0; 1: mux_10028 = v_10029;
    endcase
  endfunction
  reg [7:0] v_10029 = 8'h0;
  wire [7:0] v_10030;
  wire [7:0] v_10031;
  function [7:0] mux_10031(input [0:0] sel);
    case (sel) 0: mux_10031 = 8'h0; 1: mux_10031 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10032;
  wire [7:0] v_10033;
  wire [7:0] v_10034;
  function [7:0] mux_10034(input [0:0] sel);
    case (sel) 0: mux_10034 = 8'h0; 1: mux_10034 = v_10035;
    endcase
  endfunction
  reg [7:0] v_10035 = 8'h0;
  wire [7:0] v_10036;
  wire [7:0] v_10037;
  function [7:0] mux_10037(input [0:0] sel);
    case (sel) 0: mux_10037 = 8'h0; 1: mux_10037 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10038;
  wire [7:0] v_10039;
  wire [7:0] v_10040;
  function [7:0] mux_10040(input [0:0] sel);
    case (sel) 0: mux_10040 = 8'h0; 1: mux_10040 = vout_peek_2013;
    endcase
  endfunction
  wire [7:0] v_10041;
  function [7:0] mux_10041(input [0:0] sel);
    case (sel) 0: mux_10041 = 8'h0; 1: mux_10041 = vout_peek_2005;
    endcase
  endfunction
  wire [7:0] v_10042;
  function [7:0] mux_10042(input [0:0] sel);
    case (sel) 0: mux_10042 = 8'h0; 1: mux_10042 = v_10043;
    endcase
  endfunction
  reg [7:0] v_10043 = 8'h0;
  wire [7:0] v_10044;
  wire [7:0] v_10045;
  function [7:0] mux_10045(input [0:0] sel);
    case (sel) 0: mux_10045 = 8'h0; 1: mux_10045 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10046;
  wire [7:0] v_10047;
  wire [7:0] v_10048;
  function [7:0] mux_10048(input [0:0] sel);
    case (sel) 0: mux_10048 = 8'h0; 1: mux_10048 = vout_peek_1999;
    endcase
  endfunction
  wire [7:0] v_10049;
  function [7:0] mux_10049(input [0:0] sel);
    case (sel) 0: mux_10049 = 8'h0; 1: mux_10049 = vout_peek_1991;
    endcase
  endfunction
  wire [7:0] v_10050;
  function [7:0] mux_10050(input [0:0] sel);
    case (sel) 0: mux_10050 = 8'h0; 1: mux_10050 = v_10051;
    endcase
  endfunction
  reg [7:0] v_10051 = 8'h0;
  wire [7:0] v_10052;
  wire [7:0] v_10053;
  function [7:0] mux_10053(input [0:0] sel);
    case (sel) 0: mux_10053 = 8'h0; 1: mux_10053 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10054;
  wire [7:0] v_10055;
  wire [7:0] v_10056;
  function [7:0] mux_10056(input [0:0] sel);
    case (sel) 0: mux_10056 = 8'h0; 1: mux_10056 = v_10057;
    endcase
  endfunction
  reg [7:0] v_10057 = 8'h0;
  wire [7:0] v_10058;
  wire [7:0] v_10059;
  function [7:0] mux_10059(input [0:0] sel);
    case (sel) 0: mux_10059 = 8'h0; 1: mux_10059 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10060;
  wire [7:0] v_10061;
  wire [7:0] v_10062;
  function [7:0] mux_10062(input [0:0] sel);
    case (sel) 0: mux_10062 = 8'h0; 1: mux_10062 = vout_peek_1985;
    endcase
  endfunction
  wire [7:0] v_10063;
  function [7:0] mux_10063(input [0:0] sel);
    case (sel) 0: mux_10063 = 8'h0; 1: mux_10063 = vout_peek_1977;
    endcase
  endfunction
  wire [7:0] v_10064;
  function [7:0] mux_10064(input [0:0] sel);
    case (sel) 0: mux_10064 = 8'h0; 1: mux_10064 = v_10065;
    endcase
  endfunction
  reg [7:0] v_10065 = 8'h0;
  wire [7:0] v_10066;
  wire [7:0] v_10067;
  function [7:0] mux_10067(input [0:0] sel);
    case (sel) 0: mux_10067 = 8'h0; 1: mux_10067 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10068;
  wire [7:0] v_10069;
  wire [7:0] v_10070;
  function [7:0] mux_10070(input [0:0] sel);
    case (sel) 0: mux_10070 = 8'h0; 1: mux_10070 = vout_peek_1971;
    endcase
  endfunction
  wire [7:0] v_10071;
  function [7:0] mux_10071(input [0:0] sel);
    case (sel) 0: mux_10071 = 8'h0; 1: mux_10071 = vout_peek_1963;
    endcase
  endfunction
  wire [7:0] v_10072;
  function [7:0] mux_10072(input [0:0] sel);
    case (sel) 0: mux_10072 = 8'h0; 1: mux_10072 = v_10073;
    endcase
  endfunction
  reg [7:0] v_10073 = 8'h0;
  wire [7:0] v_10074;
  wire [7:0] v_10075;
  function [7:0] mux_10075(input [0:0] sel);
    case (sel) 0: mux_10075 = 8'h0; 1: mux_10075 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10076;
  wire [7:0] v_10077;
  wire [7:0] v_10078;
  function [7:0] mux_10078(input [0:0] sel);
    case (sel) 0: mux_10078 = 8'h0; 1: mux_10078 = v_10079;
    endcase
  endfunction
  reg [7:0] v_10079 = 8'h0;
  wire [7:0] v_10080;
  wire [7:0] v_10081;
  function [7:0] mux_10081(input [0:0] sel);
    case (sel) 0: mux_10081 = 8'h0; 1: mux_10081 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10082;
  wire [7:0] v_10083;
  wire [7:0] v_10084;
  function [7:0] mux_10084(input [0:0] sel);
    case (sel) 0: mux_10084 = 8'h0; 1: mux_10084 = v_10085;
    endcase
  endfunction
  reg [7:0] v_10085 = 8'h0;
  wire [7:0] v_10086;
  wire [7:0] v_10087;
  function [7:0] mux_10087(input [0:0] sel);
    case (sel) 0: mux_10087 = 8'h0; 1: mux_10087 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10088;
  wire [7:0] v_10089;
  wire [7:0] v_10090;
  function [7:0] mux_10090(input [0:0] sel);
    case (sel) 0: mux_10090 = 8'h0; 1: mux_10090 = vout_peek_1957;
    endcase
  endfunction
  wire [7:0] v_10091;
  function [7:0] mux_10091(input [0:0] sel);
    case (sel) 0: mux_10091 = 8'h0; 1: mux_10091 = vout_peek_1949;
    endcase
  endfunction
  wire [7:0] v_10092;
  function [7:0] mux_10092(input [0:0] sel);
    case (sel) 0: mux_10092 = 8'h0; 1: mux_10092 = v_10093;
    endcase
  endfunction
  reg [7:0] v_10093 = 8'h0;
  wire [7:0] v_10094;
  wire [7:0] v_10095;
  function [7:0] mux_10095(input [0:0] sel);
    case (sel) 0: mux_10095 = 8'h0; 1: mux_10095 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10096;
  wire [7:0] v_10097;
  wire [7:0] v_10098;
  function [7:0] mux_10098(input [0:0] sel);
    case (sel) 0: mux_10098 = 8'h0; 1: mux_10098 = vout_peek_1943;
    endcase
  endfunction
  wire [7:0] v_10099;
  function [7:0] mux_10099(input [0:0] sel);
    case (sel) 0: mux_10099 = 8'h0; 1: mux_10099 = vout_peek_1935;
    endcase
  endfunction
  wire [7:0] v_10100;
  function [7:0] mux_10100(input [0:0] sel);
    case (sel) 0: mux_10100 = 8'h0; 1: mux_10100 = v_10101;
    endcase
  endfunction
  reg [7:0] v_10101 = 8'h0;
  wire [7:0] v_10102;
  wire [7:0] v_10103;
  function [7:0] mux_10103(input [0:0] sel);
    case (sel) 0: mux_10103 = 8'h0; 1: mux_10103 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10104;
  wire [7:0] v_10105;
  wire [7:0] v_10106;
  function [7:0] mux_10106(input [0:0] sel);
    case (sel) 0: mux_10106 = 8'h0; 1: mux_10106 = v_10107;
    endcase
  endfunction
  reg [7:0] v_10107 = 8'h0;
  wire [7:0] v_10108;
  wire [7:0] v_10109;
  function [7:0] mux_10109(input [0:0] sel);
    case (sel) 0: mux_10109 = 8'h0; 1: mux_10109 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10110;
  wire [7:0] v_10111;
  wire [7:0] v_10112;
  function [7:0] mux_10112(input [0:0] sel);
    case (sel) 0: mux_10112 = 8'h0; 1: mux_10112 = vout_peek_1929;
    endcase
  endfunction
  wire [7:0] v_10113;
  function [7:0] mux_10113(input [0:0] sel);
    case (sel) 0: mux_10113 = 8'h0; 1: mux_10113 = vout_peek_1921;
    endcase
  endfunction
  wire [7:0] v_10114;
  function [7:0] mux_10114(input [0:0] sel);
    case (sel) 0: mux_10114 = 8'h0; 1: mux_10114 = v_10115;
    endcase
  endfunction
  reg [7:0] v_10115 = 8'h0;
  wire [7:0] v_10116;
  wire [7:0] v_10117;
  function [7:0] mux_10117(input [0:0] sel);
    case (sel) 0: mux_10117 = 8'h0; 1: mux_10117 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10118;
  wire [7:0] v_10119;
  wire [7:0] v_10120;
  function [7:0] mux_10120(input [0:0] sel);
    case (sel) 0: mux_10120 = 8'h0; 1: mux_10120 = vout_peek_1915;
    endcase
  endfunction
  wire [7:0] v_10121;
  function [7:0] mux_10121(input [0:0] sel);
    case (sel) 0: mux_10121 = 8'h0; 1: mux_10121 = vout_peek_1907;
    endcase
  endfunction
  wire [7:0] v_10122;
  function [7:0] mux_10122(input [0:0] sel);
    case (sel) 0: mux_10122 = 8'h0; 1: mux_10122 = v_10123;
    endcase
  endfunction
  reg [7:0] v_10123 = 8'h0;
  wire [7:0] v_10124;
  wire [7:0] v_10125;
  function [7:0] mux_10125(input [0:0] sel);
    case (sel) 0: mux_10125 = 8'h0; 1: mux_10125 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10126;
  wire [7:0] v_10127;
  wire [7:0] v_10128;
  function [7:0] mux_10128(input [0:0] sel);
    case (sel) 0: mux_10128 = 8'h0; 1: mux_10128 = v_10129;
    endcase
  endfunction
  reg [7:0] v_10129 = 8'h0;
  wire [7:0] v_10130;
  wire [7:0] v_10131;
  function [7:0] mux_10131(input [0:0] sel);
    case (sel) 0: mux_10131 = 8'h0; 1: mux_10131 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10132;
  wire [7:0] v_10133;
  wire [7:0] v_10134;
  function [7:0] mux_10134(input [0:0] sel);
    case (sel) 0: mux_10134 = 8'h0; 1: mux_10134 = v_10135;
    endcase
  endfunction
  reg [7:0] v_10135 = 8'h0;
  wire [7:0] v_10136;
  wire [7:0] v_10137;
  function [7:0] mux_10137(input [0:0] sel);
    case (sel) 0: mux_10137 = 8'h0; 1: mux_10137 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10138;
  wire [7:0] v_10139;
  wire [7:0] v_10140;
  function [7:0] mux_10140(input [0:0] sel);
    case (sel) 0: mux_10140 = 8'h0; 1: mux_10140 = v_10141;
    endcase
  endfunction
  reg [7:0] v_10141 = 8'h0;
  wire [7:0] v_10142;
  wire [7:0] v_10143;
  function [7:0] mux_10143(input [0:0] sel);
    case (sel) 0: mux_10143 = 8'h0; 1: mux_10143 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10144;
  wire [7:0] v_10145;
  wire [7:0] v_10146;
  function [7:0] mux_10146(input [0:0] sel);
    case (sel) 0: mux_10146 = 8'h0; 1: mux_10146 = vout_peek_1901;
    endcase
  endfunction
  wire [7:0] v_10147;
  function [7:0] mux_10147(input [0:0] sel);
    case (sel) 0: mux_10147 = 8'h0; 1: mux_10147 = vout_peek_1893;
    endcase
  endfunction
  wire [7:0] v_10148;
  function [7:0] mux_10148(input [0:0] sel);
    case (sel) 0: mux_10148 = 8'h0; 1: mux_10148 = v_10149;
    endcase
  endfunction
  reg [7:0] v_10149 = 8'h0;
  wire [7:0] v_10150;
  wire [7:0] v_10151;
  function [7:0] mux_10151(input [0:0] sel);
    case (sel) 0: mux_10151 = 8'h0; 1: mux_10151 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10152;
  wire [7:0] v_10153;
  wire [7:0] v_10154;
  function [7:0] mux_10154(input [0:0] sel);
    case (sel) 0: mux_10154 = 8'h0; 1: mux_10154 = vout_peek_1887;
    endcase
  endfunction
  wire [7:0] v_10155;
  function [7:0] mux_10155(input [0:0] sel);
    case (sel) 0: mux_10155 = 8'h0; 1: mux_10155 = vout_peek_1879;
    endcase
  endfunction
  wire [7:0] v_10156;
  function [7:0] mux_10156(input [0:0] sel);
    case (sel) 0: mux_10156 = 8'h0; 1: mux_10156 = v_10157;
    endcase
  endfunction
  reg [7:0] v_10157 = 8'h0;
  wire [7:0] v_10158;
  wire [7:0] v_10159;
  function [7:0] mux_10159(input [0:0] sel);
    case (sel) 0: mux_10159 = 8'h0; 1: mux_10159 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10160;
  wire [7:0] v_10161;
  wire [7:0] v_10162;
  function [7:0] mux_10162(input [0:0] sel);
    case (sel) 0: mux_10162 = 8'h0; 1: mux_10162 = v_10163;
    endcase
  endfunction
  reg [7:0] v_10163 = 8'h0;
  wire [7:0] v_10164;
  wire [7:0] v_10165;
  function [7:0] mux_10165(input [0:0] sel);
    case (sel) 0: mux_10165 = 8'h0; 1: mux_10165 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10166;
  wire [7:0] v_10167;
  wire [7:0] v_10168;
  function [7:0] mux_10168(input [0:0] sel);
    case (sel) 0: mux_10168 = 8'h0; 1: mux_10168 = vout_peek_1873;
    endcase
  endfunction
  wire [7:0] v_10169;
  function [7:0] mux_10169(input [0:0] sel);
    case (sel) 0: mux_10169 = 8'h0; 1: mux_10169 = vout_peek_1865;
    endcase
  endfunction
  wire [7:0] v_10170;
  function [7:0] mux_10170(input [0:0] sel);
    case (sel) 0: mux_10170 = 8'h0; 1: mux_10170 = v_10171;
    endcase
  endfunction
  reg [7:0] v_10171 = 8'h0;
  wire [7:0] v_10172;
  wire [7:0] v_10173;
  function [7:0] mux_10173(input [0:0] sel);
    case (sel) 0: mux_10173 = 8'h0; 1: mux_10173 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10174;
  wire [7:0] v_10175;
  wire [7:0] v_10176;
  function [7:0] mux_10176(input [0:0] sel);
    case (sel) 0: mux_10176 = 8'h0; 1: mux_10176 = vout_peek_1859;
    endcase
  endfunction
  wire [7:0] v_10177;
  function [7:0] mux_10177(input [0:0] sel);
    case (sel) 0: mux_10177 = 8'h0; 1: mux_10177 = vout_peek_1851;
    endcase
  endfunction
  wire [7:0] v_10178;
  function [7:0] mux_10178(input [0:0] sel);
    case (sel) 0: mux_10178 = 8'h0; 1: mux_10178 = v_10179;
    endcase
  endfunction
  reg [7:0] v_10179 = 8'h0;
  wire [7:0] v_10180;
  wire [7:0] v_10181;
  function [7:0] mux_10181(input [0:0] sel);
    case (sel) 0: mux_10181 = 8'h0; 1: mux_10181 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10182;
  wire [7:0] v_10183;
  wire [7:0] v_10184;
  function [7:0] mux_10184(input [0:0] sel);
    case (sel) 0: mux_10184 = 8'h0; 1: mux_10184 = v_10185;
    endcase
  endfunction
  reg [7:0] v_10185 = 8'h0;
  wire [7:0] v_10186;
  wire [7:0] v_10187;
  function [7:0] mux_10187(input [0:0] sel);
    case (sel) 0: mux_10187 = 8'h0; 1: mux_10187 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10188;
  wire [7:0] v_10189;
  wire [7:0] v_10190;
  function [7:0] mux_10190(input [0:0] sel);
    case (sel) 0: mux_10190 = 8'h0; 1: mux_10190 = v_10191;
    endcase
  endfunction
  reg [7:0] v_10191 = 8'h0;
  wire [7:0] v_10192;
  wire [7:0] v_10193;
  function [7:0] mux_10193(input [0:0] sel);
    case (sel) 0: mux_10193 = 8'h0; 1: mux_10193 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10194;
  wire [7:0] v_10195;
  wire [7:0] v_10196;
  function [7:0] mux_10196(input [0:0] sel);
    case (sel) 0: mux_10196 = 8'h0; 1: mux_10196 = vout_peek_1845;
    endcase
  endfunction
  wire [7:0] v_10197;
  function [7:0] mux_10197(input [0:0] sel);
    case (sel) 0: mux_10197 = 8'h0; 1: mux_10197 = vout_peek_1837;
    endcase
  endfunction
  wire [7:0] v_10198;
  function [7:0] mux_10198(input [0:0] sel);
    case (sel) 0: mux_10198 = 8'h0; 1: mux_10198 = v_10199;
    endcase
  endfunction
  reg [7:0] v_10199 = 8'h0;
  wire [7:0] v_10200;
  wire [7:0] v_10201;
  function [7:0] mux_10201(input [0:0] sel);
    case (sel) 0: mux_10201 = 8'h0; 1: mux_10201 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10202;
  wire [7:0] v_10203;
  wire [7:0] v_10204;
  function [7:0] mux_10204(input [0:0] sel);
    case (sel) 0: mux_10204 = 8'h0; 1: mux_10204 = vout_peek_1831;
    endcase
  endfunction
  wire [7:0] v_10205;
  function [7:0] mux_10205(input [0:0] sel);
    case (sel) 0: mux_10205 = 8'h0; 1: mux_10205 = vout_peek_1823;
    endcase
  endfunction
  wire [7:0] v_10206;
  function [7:0] mux_10206(input [0:0] sel);
    case (sel) 0: mux_10206 = 8'h0; 1: mux_10206 = v_10207;
    endcase
  endfunction
  reg [7:0] v_10207 = 8'h0;
  wire [7:0] v_10208;
  wire [7:0] v_10209;
  function [7:0] mux_10209(input [0:0] sel);
    case (sel) 0: mux_10209 = 8'h0; 1: mux_10209 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10210;
  wire [7:0] v_10211;
  wire [7:0] v_10212;
  function [7:0] mux_10212(input [0:0] sel);
    case (sel) 0: mux_10212 = 8'h0; 1: mux_10212 = v_10213;
    endcase
  endfunction
  reg [7:0] v_10213 = 8'h0;
  wire [7:0] v_10214;
  wire [7:0] v_10215;
  function [7:0] mux_10215(input [0:0] sel);
    case (sel) 0: mux_10215 = 8'h0; 1: mux_10215 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10216;
  wire [7:0] v_10217;
  wire [7:0] v_10218;
  function [7:0] mux_10218(input [0:0] sel);
    case (sel) 0: mux_10218 = 8'h0; 1: mux_10218 = vout_peek_1817;
    endcase
  endfunction
  wire [7:0] v_10219;
  function [7:0] mux_10219(input [0:0] sel);
    case (sel) 0: mux_10219 = 8'h0; 1: mux_10219 = vout_peek_1809;
    endcase
  endfunction
  wire [7:0] v_10220;
  function [7:0] mux_10220(input [0:0] sel);
    case (sel) 0: mux_10220 = 8'h0; 1: mux_10220 = v_10221;
    endcase
  endfunction
  reg [7:0] v_10221 = 8'h0;
  wire [7:0] v_10222;
  wire [7:0] v_10223;
  function [7:0] mux_10223(input [0:0] sel);
    case (sel) 0: mux_10223 = 8'h0; 1: mux_10223 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10224;
  wire [7:0] v_10225;
  wire [7:0] v_10226;
  function [7:0] mux_10226(input [0:0] sel);
    case (sel) 0: mux_10226 = 8'h0; 1: mux_10226 = vout_peek_1803;
    endcase
  endfunction
  wire [7:0] v_10227;
  function [7:0] mux_10227(input [0:0] sel);
    case (sel) 0: mux_10227 = 8'h0; 1: mux_10227 = vout_peek_1795;
    endcase
  endfunction
  wire [7:0] v_10228;
  function [7:0] mux_10228(input [0:0] sel);
    case (sel) 0: mux_10228 = 8'h0; 1: mux_10228 = v_10229;
    endcase
  endfunction
  reg [7:0] v_10229 = 8'h0;
  wire [7:0] v_10230;
  wire [7:0] v_10231;
  function [7:0] mux_10231(input [0:0] sel);
    case (sel) 0: mux_10231 = 8'h0; 1: mux_10231 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10232;
  wire [7:0] v_10233;
  wire [7:0] v_10234;
  function [7:0] mux_10234(input [0:0] sel);
    case (sel) 0: mux_10234 = 8'h0; 1: mux_10234 = v_10235;
    endcase
  endfunction
  reg [7:0] v_10235 = 8'h0;
  wire [7:0] v_10236;
  wire [7:0] v_10237;
  function [7:0] mux_10237(input [0:0] sel);
    case (sel) 0: mux_10237 = 8'h0; 1: mux_10237 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10238;
  wire [7:0] v_10239;
  wire [7:0] v_10240;
  function [7:0] mux_10240(input [0:0] sel);
    case (sel) 0: mux_10240 = 8'h0; 1: mux_10240 = v_10241;
    endcase
  endfunction
  reg [7:0] v_10241 = 8'h0;
  wire [7:0] v_10242;
  wire [7:0] v_10243;
  function [7:0] mux_10243(input [0:0] sel);
    case (sel) 0: mux_10243 = 8'h0; 1: mux_10243 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10244;
  wire [7:0] v_10245;
  wire [7:0] v_10246;
  function [7:0] mux_10246(input [0:0] sel);
    case (sel) 0: mux_10246 = 8'h0; 1: mux_10246 = v_10247;
    endcase
  endfunction
  reg [7:0] v_10247 = 8'h0;
  wire [7:0] v_10248;
  wire [7:0] v_10249;
  function [7:0] mux_10249(input [0:0] sel);
    case (sel) 0: mux_10249 = 8'h0; 1: mux_10249 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10250;
  wire [7:0] v_10251;
  wire [7:0] v_10252;
  function [7:0] mux_10252(input [0:0] sel);
    case (sel) 0: mux_10252 = 8'h0; 1: mux_10252 = v_10253;
    endcase
  endfunction
  reg [7:0] v_10253 = 8'h0;
  wire [7:0] v_10254;
  wire [7:0] v_10255;
  function [7:0] mux_10255(input [0:0] sel);
    case (sel) 0: mux_10255 = 8'h0; 1: mux_10255 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10256;
  wire [7:0] v_10257;
  wire [7:0] v_10258;
  function [7:0] mux_10258(input [0:0] sel);
    case (sel) 0: mux_10258 = 8'h0; 1: mux_10258 = vout_peek_1789;
    endcase
  endfunction
  wire [7:0] v_10259;
  function [7:0] mux_10259(input [0:0] sel);
    case (sel) 0: mux_10259 = 8'h0; 1: mux_10259 = vout_peek_1781;
    endcase
  endfunction
  wire [7:0] v_10260;
  function [7:0] mux_10260(input [0:0] sel);
    case (sel) 0: mux_10260 = 8'h0; 1: mux_10260 = v_10261;
    endcase
  endfunction
  reg [7:0] v_10261 = 8'h0;
  wire [7:0] v_10262;
  wire [7:0] v_10263;
  function [7:0] mux_10263(input [0:0] sel);
    case (sel) 0: mux_10263 = 8'h0; 1: mux_10263 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10264;
  wire [7:0] v_10265;
  wire [7:0] v_10266;
  function [7:0] mux_10266(input [0:0] sel);
    case (sel) 0: mux_10266 = 8'h0; 1: mux_10266 = vout_peek_1775;
    endcase
  endfunction
  wire [7:0] v_10267;
  function [7:0] mux_10267(input [0:0] sel);
    case (sel) 0: mux_10267 = 8'h0; 1: mux_10267 = vout_peek_1767;
    endcase
  endfunction
  wire [7:0] v_10268;
  function [7:0] mux_10268(input [0:0] sel);
    case (sel) 0: mux_10268 = 8'h0; 1: mux_10268 = v_10269;
    endcase
  endfunction
  reg [7:0] v_10269 = 8'h0;
  wire [7:0] v_10270;
  wire [7:0] v_10271;
  function [7:0] mux_10271(input [0:0] sel);
    case (sel) 0: mux_10271 = 8'h0; 1: mux_10271 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10272;
  wire [7:0] v_10273;
  wire [7:0] v_10274;
  function [7:0] mux_10274(input [0:0] sel);
    case (sel) 0: mux_10274 = 8'h0; 1: mux_10274 = v_10275;
    endcase
  endfunction
  reg [7:0] v_10275 = 8'h0;
  wire [7:0] v_10276;
  wire [7:0] v_10277;
  function [7:0] mux_10277(input [0:0] sel);
    case (sel) 0: mux_10277 = 8'h0; 1: mux_10277 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10278;
  wire [7:0] v_10279;
  wire [7:0] v_10280;
  function [7:0] mux_10280(input [0:0] sel);
    case (sel) 0: mux_10280 = 8'h0; 1: mux_10280 = vout_peek_1761;
    endcase
  endfunction
  wire [7:0] v_10281;
  function [7:0] mux_10281(input [0:0] sel);
    case (sel) 0: mux_10281 = 8'h0; 1: mux_10281 = vout_peek_1753;
    endcase
  endfunction
  wire [7:0] v_10282;
  function [7:0] mux_10282(input [0:0] sel);
    case (sel) 0: mux_10282 = 8'h0; 1: mux_10282 = v_10283;
    endcase
  endfunction
  reg [7:0] v_10283 = 8'h0;
  wire [7:0] v_10284;
  wire [7:0] v_10285;
  function [7:0] mux_10285(input [0:0] sel);
    case (sel) 0: mux_10285 = 8'h0; 1: mux_10285 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10286;
  wire [7:0] v_10287;
  wire [7:0] v_10288;
  function [7:0] mux_10288(input [0:0] sel);
    case (sel) 0: mux_10288 = 8'h0; 1: mux_10288 = vout_peek_1747;
    endcase
  endfunction
  wire [7:0] v_10289;
  function [7:0] mux_10289(input [0:0] sel);
    case (sel) 0: mux_10289 = 8'h0; 1: mux_10289 = vout_peek_1739;
    endcase
  endfunction
  wire [7:0] v_10290;
  function [7:0] mux_10290(input [0:0] sel);
    case (sel) 0: mux_10290 = 8'h0; 1: mux_10290 = v_10291;
    endcase
  endfunction
  reg [7:0] v_10291 = 8'h0;
  wire [7:0] v_10292;
  wire [7:0] v_10293;
  function [7:0] mux_10293(input [0:0] sel);
    case (sel) 0: mux_10293 = 8'h0; 1: mux_10293 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10294;
  wire [7:0] v_10295;
  wire [7:0] v_10296;
  function [7:0] mux_10296(input [0:0] sel);
    case (sel) 0: mux_10296 = 8'h0; 1: mux_10296 = v_10297;
    endcase
  endfunction
  reg [7:0] v_10297 = 8'h0;
  wire [7:0] v_10298;
  wire [7:0] v_10299;
  function [7:0] mux_10299(input [0:0] sel);
    case (sel) 0: mux_10299 = 8'h0; 1: mux_10299 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10300;
  wire [7:0] v_10301;
  wire [7:0] v_10302;
  function [7:0] mux_10302(input [0:0] sel);
    case (sel) 0: mux_10302 = 8'h0; 1: mux_10302 = v_10303;
    endcase
  endfunction
  reg [7:0] v_10303 = 8'h0;
  wire [7:0] v_10304;
  wire [7:0] v_10305;
  function [7:0] mux_10305(input [0:0] sel);
    case (sel) 0: mux_10305 = 8'h0; 1: mux_10305 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10306;
  wire [7:0] v_10307;
  wire [7:0] v_10308;
  function [7:0] mux_10308(input [0:0] sel);
    case (sel) 0: mux_10308 = 8'h0; 1: mux_10308 = vout_peek_1733;
    endcase
  endfunction
  wire [7:0] v_10309;
  function [7:0] mux_10309(input [0:0] sel);
    case (sel) 0: mux_10309 = 8'h0; 1: mux_10309 = vout_peek_1725;
    endcase
  endfunction
  wire [7:0] v_10310;
  function [7:0] mux_10310(input [0:0] sel);
    case (sel) 0: mux_10310 = 8'h0; 1: mux_10310 = v_10311;
    endcase
  endfunction
  reg [7:0] v_10311 = 8'h0;
  wire [7:0] v_10312;
  wire [7:0] v_10313;
  function [7:0] mux_10313(input [0:0] sel);
    case (sel) 0: mux_10313 = 8'h0; 1: mux_10313 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10314;
  wire [7:0] v_10315;
  wire [7:0] v_10316;
  function [7:0] mux_10316(input [0:0] sel);
    case (sel) 0: mux_10316 = 8'h0; 1: mux_10316 = vout_peek_1719;
    endcase
  endfunction
  wire [7:0] v_10317;
  function [7:0] mux_10317(input [0:0] sel);
    case (sel) 0: mux_10317 = 8'h0; 1: mux_10317 = vout_peek_1711;
    endcase
  endfunction
  wire [7:0] v_10318;
  function [7:0] mux_10318(input [0:0] sel);
    case (sel) 0: mux_10318 = 8'h0; 1: mux_10318 = v_10319;
    endcase
  endfunction
  reg [7:0] v_10319 = 8'h0;
  wire [7:0] v_10320;
  wire [7:0] v_10321;
  function [7:0] mux_10321(input [0:0] sel);
    case (sel) 0: mux_10321 = 8'h0; 1: mux_10321 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10322;
  wire [7:0] v_10323;
  wire [7:0] v_10324;
  function [7:0] mux_10324(input [0:0] sel);
    case (sel) 0: mux_10324 = 8'h0; 1: mux_10324 = v_10325;
    endcase
  endfunction
  reg [7:0] v_10325 = 8'h0;
  wire [7:0] v_10326;
  wire [7:0] v_10327;
  function [7:0] mux_10327(input [0:0] sel);
    case (sel) 0: mux_10327 = 8'h0; 1: mux_10327 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10328;
  wire [7:0] v_10329;
  wire [7:0] v_10330;
  function [7:0] mux_10330(input [0:0] sel);
    case (sel) 0: mux_10330 = 8'h0; 1: mux_10330 = vout_peek_1705;
    endcase
  endfunction
  wire [7:0] v_10331;
  function [7:0] mux_10331(input [0:0] sel);
    case (sel) 0: mux_10331 = 8'h0; 1: mux_10331 = vout_peek_1697;
    endcase
  endfunction
  wire [7:0] v_10332;
  function [7:0] mux_10332(input [0:0] sel);
    case (sel) 0: mux_10332 = 8'h0; 1: mux_10332 = v_10333;
    endcase
  endfunction
  reg [7:0] v_10333 = 8'h0;
  wire [7:0] v_10334;
  wire [7:0] v_10335;
  function [7:0] mux_10335(input [0:0] sel);
    case (sel) 0: mux_10335 = 8'h0; 1: mux_10335 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10336;
  wire [7:0] v_10337;
  wire [7:0] v_10338;
  function [7:0] mux_10338(input [0:0] sel);
    case (sel) 0: mux_10338 = 8'h0; 1: mux_10338 = vout_peek_1691;
    endcase
  endfunction
  wire [7:0] v_10339;
  function [7:0] mux_10339(input [0:0] sel);
    case (sel) 0: mux_10339 = 8'h0; 1: mux_10339 = vout_peek_1683;
    endcase
  endfunction
  wire [7:0] v_10340;
  function [7:0] mux_10340(input [0:0] sel);
    case (sel) 0: mux_10340 = 8'h0; 1: mux_10340 = v_10341;
    endcase
  endfunction
  reg [7:0] v_10341 = 8'h0;
  wire [7:0] v_10342;
  wire [7:0] v_10343;
  function [7:0] mux_10343(input [0:0] sel);
    case (sel) 0: mux_10343 = 8'h0; 1: mux_10343 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10344;
  wire [7:0] v_10345;
  wire [7:0] v_10346;
  function [7:0] mux_10346(input [0:0] sel);
    case (sel) 0: mux_10346 = 8'h0; 1: mux_10346 = v_10347;
    endcase
  endfunction
  reg [7:0] v_10347 = 8'h0;
  wire [7:0] v_10348;
  wire [7:0] v_10349;
  function [7:0] mux_10349(input [0:0] sel);
    case (sel) 0: mux_10349 = 8'h0; 1: mux_10349 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10350;
  wire [7:0] v_10351;
  wire [7:0] v_10352;
  function [7:0] mux_10352(input [0:0] sel);
    case (sel) 0: mux_10352 = 8'h0; 1: mux_10352 = v_10353;
    endcase
  endfunction
  reg [7:0] v_10353 = 8'h0;
  wire [7:0] v_10354;
  wire [7:0] v_10355;
  function [7:0] mux_10355(input [0:0] sel);
    case (sel) 0: mux_10355 = 8'h0; 1: mux_10355 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10356;
  wire [7:0] v_10357;
  wire [7:0] v_10358;
  function [7:0] mux_10358(input [0:0] sel);
    case (sel) 0: mux_10358 = 8'h0; 1: mux_10358 = v_10359;
    endcase
  endfunction
  reg [7:0] v_10359 = 8'h0;
  wire [7:0] v_10360;
  wire [7:0] v_10361;
  function [7:0] mux_10361(input [0:0] sel);
    case (sel) 0: mux_10361 = 8'h0; 1: mux_10361 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10362;
  wire [7:0] v_10363;
  wire [7:0] v_10364;
  function [7:0] mux_10364(input [0:0] sel);
    case (sel) 0: mux_10364 = 8'h0; 1: mux_10364 = vout_peek_1677;
    endcase
  endfunction
  wire [7:0] v_10365;
  function [7:0] mux_10365(input [0:0] sel);
    case (sel) 0: mux_10365 = 8'h0; 1: mux_10365 = vout_peek_1669;
    endcase
  endfunction
  wire [7:0] v_10366;
  function [7:0] mux_10366(input [0:0] sel);
    case (sel) 0: mux_10366 = 8'h0; 1: mux_10366 = v_10367;
    endcase
  endfunction
  reg [7:0] v_10367 = 8'h0;
  wire [7:0] v_10368;
  wire [7:0] v_10369;
  function [7:0] mux_10369(input [0:0] sel);
    case (sel) 0: mux_10369 = 8'h0; 1: mux_10369 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10370;
  wire [7:0] v_10371;
  wire [7:0] v_10372;
  function [7:0] mux_10372(input [0:0] sel);
    case (sel) 0: mux_10372 = 8'h0; 1: mux_10372 = vout_peek_1663;
    endcase
  endfunction
  wire [7:0] v_10373;
  function [7:0] mux_10373(input [0:0] sel);
    case (sel) 0: mux_10373 = 8'h0; 1: mux_10373 = vout_peek_1655;
    endcase
  endfunction
  wire [7:0] v_10374;
  function [7:0] mux_10374(input [0:0] sel);
    case (sel) 0: mux_10374 = 8'h0; 1: mux_10374 = v_10375;
    endcase
  endfunction
  reg [7:0] v_10375 = 8'h0;
  wire [7:0] v_10376;
  wire [7:0] v_10377;
  function [7:0] mux_10377(input [0:0] sel);
    case (sel) 0: mux_10377 = 8'h0; 1: mux_10377 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10378;
  wire [7:0] v_10379;
  wire [7:0] v_10380;
  function [7:0] mux_10380(input [0:0] sel);
    case (sel) 0: mux_10380 = 8'h0; 1: mux_10380 = v_10381;
    endcase
  endfunction
  reg [7:0] v_10381 = 8'h0;
  wire [7:0] v_10382;
  wire [7:0] v_10383;
  function [7:0] mux_10383(input [0:0] sel);
    case (sel) 0: mux_10383 = 8'h0; 1: mux_10383 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10384;
  wire [7:0] v_10385;
  wire [7:0] v_10386;
  function [7:0] mux_10386(input [0:0] sel);
    case (sel) 0: mux_10386 = 8'h0; 1: mux_10386 = vout_peek_1649;
    endcase
  endfunction
  wire [7:0] v_10387;
  function [7:0] mux_10387(input [0:0] sel);
    case (sel) 0: mux_10387 = 8'h0; 1: mux_10387 = vout_peek_1641;
    endcase
  endfunction
  wire [7:0] v_10388;
  function [7:0] mux_10388(input [0:0] sel);
    case (sel) 0: mux_10388 = 8'h0; 1: mux_10388 = v_10389;
    endcase
  endfunction
  reg [7:0] v_10389 = 8'h0;
  wire [7:0] v_10390;
  wire [7:0] v_10391;
  function [7:0] mux_10391(input [0:0] sel);
    case (sel) 0: mux_10391 = 8'h0; 1: mux_10391 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10392;
  wire [7:0] v_10393;
  wire [7:0] v_10394;
  function [7:0] mux_10394(input [0:0] sel);
    case (sel) 0: mux_10394 = 8'h0; 1: mux_10394 = vout_peek_1635;
    endcase
  endfunction
  wire [7:0] v_10395;
  function [7:0] mux_10395(input [0:0] sel);
    case (sel) 0: mux_10395 = 8'h0; 1: mux_10395 = vout_peek_1627;
    endcase
  endfunction
  wire [7:0] v_10396;
  function [7:0] mux_10396(input [0:0] sel);
    case (sel) 0: mux_10396 = 8'h0; 1: mux_10396 = v_10397;
    endcase
  endfunction
  reg [7:0] v_10397 = 8'h0;
  wire [7:0] v_10398;
  wire [7:0] v_10399;
  function [7:0] mux_10399(input [0:0] sel);
    case (sel) 0: mux_10399 = 8'h0; 1: mux_10399 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10400;
  wire [7:0] v_10401;
  wire [7:0] v_10402;
  function [7:0] mux_10402(input [0:0] sel);
    case (sel) 0: mux_10402 = 8'h0; 1: mux_10402 = v_10403;
    endcase
  endfunction
  reg [7:0] v_10403 = 8'h0;
  wire [7:0] v_10404;
  wire [7:0] v_10405;
  function [7:0] mux_10405(input [0:0] sel);
    case (sel) 0: mux_10405 = 8'h0; 1: mux_10405 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10406;
  wire [7:0] v_10407;
  wire [7:0] v_10408;
  function [7:0] mux_10408(input [0:0] sel);
    case (sel) 0: mux_10408 = 8'h0; 1: mux_10408 = v_10409;
    endcase
  endfunction
  reg [7:0] v_10409 = 8'h0;
  wire [7:0] v_10410;
  wire [7:0] v_10411;
  function [7:0] mux_10411(input [0:0] sel);
    case (sel) 0: mux_10411 = 8'h0; 1: mux_10411 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10412;
  wire [7:0] v_10413;
  wire [7:0] v_10414;
  function [7:0] mux_10414(input [0:0] sel);
    case (sel) 0: mux_10414 = 8'h0; 1: mux_10414 = vout_peek_1621;
    endcase
  endfunction
  wire [7:0] v_10415;
  function [7:0] mux_10415(input [0:0] sel);
    case (sel) 0: mux_10415 = 8'h0; 1: mux_10415 = vout_peek_1613;
    endcase
  endfunction
  wire [7:0] v_10416;
  function [7:0] mux_10416(input [0:0] sel);
    case (sel) 0: mux_10416 = 8'h0; 1: mux_10416 = v_10417;
    endcase
  endfunction
  reg [7:0] v_10417 = 8'h0;
  wire [7:0] v_10418;
  wire [7:0] v_10419;
  function [7:0] mux_10419(input [0:0] sel);
    case (sel) 0: mux_10419 = 8'h0; 1: mux_10419 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10420;
  wire [7:0] v_10421;
  wire [7:0] v_10422;
  function [7:0] mux_10422(input [0:0] sel);
    case (sel) 0: mux_10422 = 8'h0; 1: mux_10422 = vout_peek_1607;
    endcase
  endfunction
  wire [7:0] v_10423;
  function [7:0] mux_10423(input [0:0] sel);
    case (sel) 0: mux_10423 = 8'h0; 1: mux_10423 = vout_peek_1599;
    endcase
  endfunction
  wire [7:0] v_10424;
  function [7:0] mux_10424(input [0:0] sel);
    case (sel) 0: mux_10424 = 8'h0; 1: mux_10424 = v_10425;
    endcase
  endfunction
  reg [7:0] v_10425 = 8'h0;
  wire [7:0] v_10426;
  wire [7:0] v_10427;
  function [7:0] mux_10427(input [0:0] sel);
    case (sel) 0: mux_10427 = 8'h0; 1: mux_10427 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10428;
  wire [7:0] v_10429;
  wire [7:0] v_10430;
  function [7:0] mux_10430(input [0:0] sel);
    case (sel) 0: mux_10430 = 8'h0; 1: mux_10430 = v_10431;
    endcase
  endfunction
  reg [7:0] v_10431 = 8'h0;
  wire [7:0] v_10432;
  wire [7:0] v_10433;
  function [7:0] mux_10433(input [0:0] sel);
    case (sel) 0: mux_10433 = 8'h0; 1: mux_10433 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10434;
  wire [7:0] v_10435;
  wire [7:0] v_10436;
  function [7:0] mux_10436(input [0:0] sel);
    case (sel) 0: mux_10436 = 8'h0; 1: mux_10436 = vout_peek_1593;
    endcase
  endfunction
  wire [7:0] v_10437;
  function [7:0] mux_10437(input [0:0] sel);
    case (sel) 0: mux_10437 = 8'h0; 1: mux_10437 = vout_peek_1585;
    endcase
  endfunction
  wire [7:0] v_10438;
  function [7:0] mux_10438(input [0:0] sel);
    case (sel) 0: mux_10438 = 8'h0; 1: mux_10438 = v_10439;
    endcase
  endfunction
  reg [7:0] v_10439 = 8'h0;
  wire [7:0] v_10440;
  wire [7:0] v_10441;
  function [7:0] mux_10441(input [0:0] sel);
    case (sel) 0: mux_10441 = 8'h0; 1: mux_10441 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10442;
  wire [7:0] v_10443;
  wire [7:0] v_10444;
  function [7:0] mux_10444(input [0:0] sel);
    case (sel) 0: mux_10444 = 8'h0; 1: mux_10444 = vout_peek_1579;
    endcase
  endfunction
  wire [7:0] v_10445;
  function [7:0] mux_10445(input [0:0] sel);
    case (sel) 0: mux_10445 = 8'h0; 1: mux_10445 = vout_peek_1571;
    endcase
  endfunction
  wire [7:0] v_10446;
  function [7:0] mux_10446(input [0:0] sel);
    case (sel) 0: mux_10446 = 8'h0; 1: mux_10446 = v_10447;
    endcase
  endfunction
  reg [7:0] v_10447 = 8'h0;
  wire [7:0] v_10448;
  wire [7:0] v_10449;
  function [7:0] mux_10449(input [0:0] sel);
    case (sel) 0: mux_10449 = 8'h0; 1: mux_10449 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10450;
  wire [7:0] v_10451;
  wire [7:0] v_10452;
  function [7:0] mux_10452(input [0:0] sel);
    case (sel) 0: mux_10452 = 8'h0; 1: mux_10452 = v_10453;
    endcase
  endfunction
  reg [7:0] v_10453 = 8'h0;
  wire [7:0] v_10454;
  wire [7:0] v_10455;
  function [7:0] mux_10455(input [0:0] sel);
    case (sel) 0: mux_10455 = 8'h0; 1: mux_10455 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10456;
  wire [7:0] v_10457;
  wire [7:0] v_10458;
  function [7:0] mux_10458(input [0:0] sel);
    case (sel) 0: mux_10458 = 8'h0; 1: mux_10458 = v_10459;
    endcase
  endfunction
  reg [7:0] v_10459 = 8'h0;
  wire [7:0] v_10460;
  wire [7:0] v_10461;
  function [7:0] mux_10461(input [0:0] sel);
    case (sel) 0: mux_10461 = 8'h0; 1: mux_10461 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10462;
  wire [7:0] v_10463;
  wire [7:0] v_10464;
  function [7:0] mux_10464(input [0:0] sel);
    case (sel) 0: mux_10464 = 8'h0; 1: mux_10464 = v_10465;
    endcase
  endfunction
  reg [7:0] v_10465 = 8'h0;
  wire [7:0] v_10466;
  wire [7:0] v_10467;
  function [7:0] mux_10467(input [0:0] sel);
    case (sel) 0: mux_10467 = 8'h0; 1: mux_10467 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10468;
  wire [7:0] v_10469;
  wire [7:0] v_10470;
  function [7:0] mux_10470(input [0:0] sel);
    case (sel) 0: mux_10470 = 8'h0; 1: mux_10470 = v_10471;
    endcase
  endfunction
  reg [7:0] v_10471 = 8'h0;
  wire [7:0] v_10472;
  wire [7:0] v_10473;
  function [7:0] mux_10473(input [0:0] sel);
    case (sel) 0: mux_10473 = 8'h0; 1: mux_10473 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10474;
  wire [7:0] v_10475;
  wire [7:0] v_10476;
  function [7:0] mux_10476(input [0:0] sel);
    case (sel) 0: mux_10476 = 8'h0; 1: mux_10476 = v_10477;
    endcase
  endfunction
  reg [7:0] v_10477 = 8'h0;
  wire [7:0] v_10478;
  wire [7:0] v_10479;
  function [7:0] mux_10479(input [0:0] sel);
    case (sel) 0: mux_10479 = 8'h0; 1: mux_10479 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10480;
  wire [7:0] v_10481;
  wire [7:0] v_10482;
  function [7:0] mux_10482(input [0:0] sel);
    case (sel) 0: mux_10482 = 8'h0; 1: mux_10482 = vout_peek_1565;
    endcase
  endfunction
  wire [7:0] v_10483;
  function [7:0] mux_10483(input [0:0] sel);
    case (sel) 0: mux_10483 = 8'h0; 1: mux_10483 = vout_peek_1557;
    endcase
  endfunction
  wire [7:0] v_10484;
  function [7:0] mux_10484(input [0:0] sel);
    case (sel) 0: mux_10484 = 8'h0; 1: mux_10484 = v_10485;
    endcase
  endfunction
  reg [7:0] v_10485 = 8'h0;
  wire [7:0] v_10486;
  wire [7:0] v_10487;
  function [7:0] mux_10487(input [0:0] sel);
    case (sel) 0: mux_10487 = 8'h0; 1: mux_10487 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10488;
  wire [7:0] v_10489;
  wire [7:0] v_10490;
  function [7:0] mux_10490(input [0:0] sel);
    case (sel) 0: mux_10490 = 8'h0; 1: mux_10490 = vout_peek_1551;
    endcase
  endfunction
  wire [7:0] v_10491;
  function [7:0] mux_10491(input [0:0] sel);
    case (sel) 0: mux_10491 = 8'h0; 1: mux_10491 = vout_peek_1543;
    endcase
  endfunction
  wire [7:0] v_10492;
  function [7:0] mux_10492(input [0:0] sel);
    case (sel) 0: mux_10492 = 8'h0; 1: mux_10492 = v_10493;
    endcase
  endfunction
  reg [7:0] v_10493 = 8'h0;
  wire [7:0] v_10494;
  wire [7:0] v_10495;
  function [7:0] mux_10495(input [0:0] sel);
    case (sel) 0: mux_10495 = 8'h0; 1: mux_10495 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10496;
  wire [7:0] v_10497;
  wire [7:0] v_10498;
  function [7:0] mux_10498(input [0:0] sel);
    case (sel) 0: mux_10498 = 8'h0; 1: mux_10498 = v_10499;
    endcase
  endfunction
  reg [7:0] v_10499 = 8'h0;
  wire [7:0] v_10500;
  wire [7:0] v_10501;
  function [7:0] mux_10501(input [0:0] sel);
    case (sel) 0: mux_10501 = 8'h0; 1: mux_10501 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10502;
  wire [7:0] v_10503;
  wire [7:0] v_10504;
  function [7:0] mux_10504(input [0:0] sel);
    case (sel) 0: mux_10504 = 8'h0; 1: mux_10504 = vout_peek_1537;
    endcase
  endfunction
  wire [7:0] v_10505;
  function [7:0] mux_10505(input [0:0] sel);
    case (sel) 0: mux_10505 = 8'h0; 1: mux_10505 = vout_peek_1529;
    endcase
  endfunction
  wire [7:0] v_10506;
  function [7:0] mux_10506(input [0:0] sel);
    case (sel) 0: mux_10506 = 8'h0; 1: mux_10506 = v_10507;
    endcase
  endfunction
  reg [7:0] v_10507 = 8'h0;
  wire [7:0] v_10508;
  wire [7:0] v_10509;
  function [7:0] mux_10509(input [0:0] sel);
    case (sel) 0: mux_10509 = 8'h0; 1: mux_10509 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10510;
  wire [7:0] v_10511;
  wire [7:0] v_10512;
  function [7:0] mux_10512(input [0:0] sel);
    case (sel) 0: mux_10512 = 8'h0; 1: mux_10512 = vout_peek_1523;
    endcase
  endfunction
  wire [7:0] v_10513;
  function [7:0] mux_10513(input [0:0] sel);
    case (sel) 0: mux_10513 = 8'h0; 1: mux_10513 = vout_peek_1515;
    endcase
  endfunction
  wire [7:0] v_10514;
  function [7:0] mux_10514(input [0:0] sel);
    case (sel) 0: mux_10514 = 8'h0; 1: mux_10514 = v_10515;
    endcase
  endfunction
  reg [7:0] v_10515 = 8'h0;
  wire [7:0] v_10516;
  wire [7:0] v_10517;
  function [7:0] mux_10517(input [0:0] sel);
    case (sel) 0: mux_10517 = 8'h0; 1: mux_10517 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10518;
  wire [7:0] v_10519;
  wire [7:0] v_10520;
  function [7:0] mux_10520(input [0:0] sel);
    case (sel) 0: mux_10520 = 8'h0; 1: mux_10520 = v_10521;
    endcase
  endfunction
  reg [7:0] v_10521 = 8'h0;
  wire [7:0] v_10522;
  wire [7:0] v_10523;
  function [7:0] mux_10523(input [0:0] sel);
    case (sel) 0: mux_10523 = 8'h0; 1: mux_10523 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10524;
  wire [7:0] v_10525;
  wire [7:0] v_10526;
  function [7:0] mux_10526(input [0:0] sel);
    case (sel) 0: mux_10526 = 8'h0; 1: mux_10526 = v_10527;
    endcase
  endfunction
  reg [7:0] v_10527 = 8'h0;
  wire [7:0] v_10528;
  wire [7:0] v_10529;
  function [7:0] mux_10529(input [0:0] sel);
    case (sel) 0: mux_10529 = 8'h0; 1: mux_10529 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10530;
  wire [7:0] v_10531;
  wire [7:0] v_10532;
  function [7:0] mux_10532(input [0:0] sel);
    case (sel) 0: mux_10532 = 8'h0; 1: mux_10532 = vout_peek_1509;
    endcase
  endfunction
  wire [7:0] v_10533;
  function [7:0] mux_10533(input [0:0] sel);
    case (sel) 0: mux_10533 = 8'h0; 1: mux_10533 = vout_peek_1501;
    endcase
  endfunction
  wire [7:0] v_10534;
  function [7:0] mux_10534(input [0:0] sel);
    case (sel) 0: mux_10534 = 8'h0; 1: mux_10534 = v_10535;
    endcase
  endfunction
  reg [7:0] v_10535 = 8'h0;
  wire [7:0] v_10536;
  wire [7:0] v_10537;
  function [7:0] mux_10537(input [0:0] sel);
    case (sel) 0: mux_10537 = 8'h0; 1: mux_10537 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10538;
  wire [7:0] v_10539;
  wire [7:0] v_10540;
  function [7:0] mux_10540(input [0:0] sel);
    case (sel) 0: mux_10540 = 8'h0; 1: mux_10540 = vout_peek_1495;
    endcase
  endfunction
  wire [7:0] v_10541;
  function [7:0] mux_10541(input [0:0] sel);
    case (sel) 0: mux_10541 = 8'h0; 1: mux_10541 = vout_peek_1487;
    endcase
  endfunction
  wire [7:0] v_10542;
  function [7:0] mux_10542(input [0:0] sel);
    case (sel) 0: mux_10542 = 8'h0; 1: mux_10542 = v_10543;
    endcase
  endfunction
  reg [7:0] v_10543 = 8'h0;
  wire [7:0] v_10544;
  wire [7:0] v_10545;
  function [7:0] mux_10545(input [0:0] sel);
    case (sel) 0: mux_10545 = 8'h0; 1: mux_10545 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10546;
  wire [7:0] v_10547;
  wire [7:0] v_10548;
  function [7:0] mux_10548(input [0:0] sel);
    case (sel) 0: mux_10548 = 8'h0; 1: mux_10548 = v_10549;
    endcase
  endfunction
  reg [7:0] v_10549 = 8'h0;
  wire [7:0] v_10550;
  wire [7:0] v_10551;
  function [7:0] mux_10551(input [0:0] sel);
    case (sel) 0: mux_10551 = 8'h0; 1: mux_10551 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10552;
  wire [7:0] v_10553;
  wire [7:0] v_10554;
  function [7:0] mux_10554(input [0:0] sel);
    case (sel) 0: mux_10554 = 8'h0; 1: mux_10554 = vout_peek_1481;
    endcase
  endfunction
  wire [7:0] v_10555;
  function [7:0] mux_10555(input [0:0] sel);
    case (sel) 0: mux_10555 = 8'h0; 1: mux_10555 = vout_peek_1473;
    endcase
  endfunction
  wire [7:0] v_10556;
  function [7:0] mux_10556(input [0:0] sel);
    case (sel) 0: mux_10556 = 8'h0; 1: mux_10556 = v_10557;
    endcase
  endfunction
  reg [7:0] v_10557 = 8'h0;
  wire [7:0] v_10558;
  wire [7:0] v_10559;
  function [7:0] mux_10559(input [0:0] sel);
    case (sel) 0: mux_10559 = 8'h0; 1: mux_10559 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10560;
  wire [7:0] v_10561;
  wire [7:0] v_10562;
  function [7:0] mux_10562(input [0:0] sel);
    case (sel) 0: mux_10562 = 8'h0; 1: mux_10562 = vout_peek_1467;
    endcase
  endfunction
  wire [7:0] v_10563;
  function [7:0] mux_10563(input [0:0] sel);
    case (sel) 0: mux_10563 = 8'h0; 1: mux_10563 = vout_peek_1459;
    endcase
  endfunction
  wire [7:0] v_10564;
  function [7:0] mux_10564(input [0:0] sel);
    case (sel) 0: mux_10564 = 8'h0; 1: mux_10564 = v_10565;
    endcase
  endfunction
  reg [7:0] v_10565 = 8'h0;
  wire [7:0] v_10566;
  wire [7:0] v_10567;
  function [7:0] mux_10567(input [0:0] sel);
    case (sel) 0: mux_10567 = 8'h0; 1: mux_10567 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10568;
  wire [7:0] v_10569;
  wire [7:0] v_10570;
  function [7:0] mux_10570(input [0:0] sel);
    case (sel) 0: mux_10570 = 8'h0; 1: mux_10570 = v_10571;
    endcase
  endfunction
  reg [7:0] v_10571 = 8'h0;
  wire [7:0] v_10572;
  wire [7:0] v_10573;
  function [7:0] mux_10573(input [0:0] sel);
    case (sel) 0: mux_10573 = 8'h0; 1: mux_10573 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10574;
  wire [7:0] v_10575;
  wire [7:0] v_10576;
  function [7:0] mux_10576(input [0:0] sel);
    case (sel) 0: mux_10576 = 8'h0; 1: mux_10576 = v_10577;
    endcase
  endfunction
  reg [7:0] v_10577 = 8'h0;
  wire [7:0] v_10578;
  wire [7:0] v_10579;
  function [7:0] mux_10579(input [0:0] sel);
    case (sel) 0: mux_10579 = 8'h0; 1: mux_10579 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10580;
  wire [7:0] v_10581;
  wire [7:0] v_10582;
  function [7:0] mux_10582(input [0:0] sel);
    case (sel) 0: mux_10582 = 8'h0; 1: mux_10582 = v_10583;
    endcase
  endfunction
  reg [7:0] v_10583 = 8'h0;
  wire [7:0] v_10584;
  wire [7:0] v_10585;
  function [7:0] mux_10585(input [0:0] sel);
    case (sel) 0: mux_10585 = 8'h0; 1: mux_10585 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10586;
  wire [7:0] v_10587;
  wire [7:0] v_10588;
  function [7:0] mux_10588(input [0:0] sel);
    case (sel) 0: mux_10588 = 8'h0; 1: mux_10588 = vout_peek_1453;
    endcase
  endfunction
  wire [7:0] v_10589;
  function [7:0] mux_10589(input [0:0] sel);
    case (sel) 0: mux_10589 = 8'h0; 1: mux_10589 = vout_peek_1445;
    endcase
  endfunction
  wire [7:0] v_10590;
  function [7:0] mux_10590(input [0:0] sel);
    case (sel) 0: mux_10590 = 8'h0; 1: mux_10590 = v_10591;
    endcase
  endfunction
  reg [7:0] v_10591 = 8'h0;
  wire [7:0] v_10592;
  wire [7:0] v_10593;
  function [7:0] mux_10593(input [0:0] sel);
    case (sel) 0: mux_10593 = 8'h0; 1: mux_10593 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10594;
  wire [7:0] v_10595;
  wire [7:0] v_10596;
  function [7:0] mux_10596(input [0:0] sel);
    case (sel) 0: mux_10596 = 8'h0; 1: mux_10596 = vout_peek_1439;
    endcase
  endfunction
  wire [7:0] v_10597;
  function [7:0] mux_10597(input [0:0] sel);
    case (sel) 0: mux_10597 = 8'h0; 1: mux_10597 = vout_peek_1431;
    endcase
  endfunction
  wire [7:0] v_10598;
  function [7:0] mux_10598(input [0:0] sel);
    case (sel) 0: mux_10598 = 8'h0; 1: mux_10598 = v_10599;
    endcase
  endfunction
  reg [7:0] v_10599 = 8'h0;
  wire [7:0] v_10600;
  wire [7:0] v_10601;
  function [7:0] mux_10601(input [0:0] sel);
    case (sel) 0: mux_10601 = 8'h0; 1: mux_10601 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10602;
  wire [7:0] v_10603;
  wire [7:0] v_10604;
  function [7:0] mux_10604(input [0:0] sel);
    case (sel) 0: mux_10604 = 8'h0; 1: mux_10604 = v_10605;
    endcase
  endfunction
  reg [7:0] v_10605 = 8'h0;
  wire [7:0] v_10606;
  wire [7:0] v_10607;
  function [7:0] mux_10607(input [0:0] sel);
    case (sel) 0: mux_10607 = 8'h0; 1: mux_10607 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10608;
  wire [7:0] v_10609;
  wire [7:0] v_10610;
  function [7:0] mux_10610(input [0:0] sel);
    case (sel) 0: mux_10610 = 8'h0; 1: mux_10610 = vout_peek_1425;
    endcase
  endfunction
  wire [7:0] v_10611;
  function [7:0] mux_10611(input [0:0] sel);
    case (sel) 0: mux_10611 = 8'h0; 1: mux_10611 = vout_peek_1417;
    endcase
  endfunction
  wire [7:0] v_10612;
  function [7:0] mux_10612(input [0:0] sel);
    case (sel) 0: mux_10612 = 8'h0; 1: mux_10612 = v_10613;
    endcase
  endfunction
  reg [7:0] v_10613 = 8'h0;
  wire [7:0] v_10614;
  wire [7:0] v_10615;
  function [7:0] mux_10615(input [0:0] sel);
    case (sel) 0: mux_10615 = 8'h0; 1: mux_10615 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10616;
  wire [7:0] v_10617;
  wire [7:0] v_10618;
  function [7:0] mux_10618(input [0:0] sel);
    case (sel) 0: mux_10618 = 8'h0; 1: mux_10618 = vout_peek_1411;
    endcase
  endfunction
  wire [7:0] v_10619;
  function [7:0] mux_10619(input [0:0] sel);
    case (sel) 0: mux_10619 = 8'h0; 1: mux_10619 = vout_peek_1403;
    endcase
  endfunction
  wire [7:0] v_10620;
  function [7:0] mux_10620(input [0:0] sel);
    case (sel) 0: mux_10620 = 8'h0; 1: mux_10620 = v_10621;
    endcase
  endfunction
  reg [7:0] v_10621 = 8'h0;
  wire [7:0] v_10622;
  wire [7:0] v_10623;
  function [7:0] mux_10623(input [0:0] sel);
    case (sel) 0: mux_10623 = 8'h0; 1: mux_10623 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10624;
  wire [7:0] v_10625;
  wire [7:0] v_10626;
  function [7:0] mux_10626(input [0:0] sel);
    case (sel) 0: mux_10626 = 8'h0; 1: mux_10626 = v_10627;
    endcase
  endfunction
  reg [7:0] v_10627 = 8'h0;
  wire [7:0] v_10628;
  wire [7:0] v_10629;
  function [7:0] mux_10629(input [0:0] sel);
    case (sel) 0: mux_10629 = 8'h0; 1: mux_10629 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10630;
  wire [7:0] v_10631;
  wire [7:0] v_10632;
  function [7:0] mux_10632(input [0:0] sel);
    case (sel) 0: mux_10632 = 8'h0; 1: mux_10632 = v_10633;
    endcase
  endfunction
  reg [7:0] v_10633 = 8'h0;
  wire [7:0] v_10634;
  wire [7:0] v_10635;
  function [7:0] mux_10635(input [0:0] sel);
    case (sel) 0: mux_10635 = 8'h0; 1: mux_10635 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10636;
  wire [7:0] v_10637;
  wire [7:0] v_10638;
  function [7:0] mux_10638(input [0:0] sel);
    case (sel) 0: mux_10638 = 8'h0; 1: mux_10638 = vout_peek_1397;
    endcase
  endfunction
  wire [7:0] v_10639;
  function [7:0] mux_10639(input [0:0] sel);
    case (sel) 0: mux_10639 = 8'h0; 1: mux_10639 = vout_peek_1389;
    endcase
  endfunction
  wire [7:0] v_10640;
  function [7:0] mux_10640(input [0:0] sel);
    case (sel) 0: mux_10640 = 8'h0; 1: mux_10640 = v_10641;
    endcase
  endfunction
  reg [7:0] v_10641 = 8'h0;
  wire [7:0] v_10642;
  wire [7:0] v_10643;
  function [7:0] mux_10643(input [0:0] sel);
    case (sel) 0: mux_10643 = 8'h0; 1: mux_10643 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10644;
  wire [7:0] v_10645;
  wire [7:0] v_10646;
  function [7:0] mux_10646(input [0:0] sel);
    case (sel) 0: mux_10646 = 8'h0; 1: mux_10646 = vout_peek_1383;
    endcase
  endfunction
  wire [7:0] v_10647;
  function [7:0] mux_10647(input [0:0] sel);
    case (sel) 0: mux_10647 = 8'h0; 1: mux_10647 = vout_peek_1375;
    endcase
  endfunction
  wire [7:0] v_10648;
  function [7:0] mux_10648(input [0:0] sel);
    case (sel) 0: mux_10648 = 8'h0; 1: mux_10648 = v_10649;
    endcase
  endfunction
  reg [7:0] v_10649 = 8'h0;
  wire [7:0] v_10650;
  wire [7:0] v_10651;
  function [7:0] mux_10651(input [0:0] sel);
    case (sel) 0: mux_10651 = 8'h0; 1: mux_10651 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10652;
  wire [7:0] v_10653;
  wire [7:0] v_10654;
  function [7:0] mux_10654(input [0:0] sel);
    case (sel) 0: mux_10654 = 8'h0; 1: mux_10654 = v_10655;
    endcase
  endfunction
  reg [7:0] v_10655 = 8'h0;
  wire [7:0] v_10656;
  wire [7:0] v_10657;
  function [7:0] mux_10657(input [0:0] sel);
    case (sel) 0: mux_10657 = 8'h0; 1: mux_10657 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10658;
  wire [7:0] v_10659;
  wire [7:0] v_10660;
  function [7:0] mux_10660(input [0:0] sel);
    case (sel) 0: mux_10660 = 8'h0; 1: mux_10660 = vout_peek_1369;
    endcase
  endfunction
  wire [7:0] v_10661;
  function [7:0] mux_10661(input [0:0] sel);
    case (sel) 0: mux_10661 = 8'h0; 1: mux_10661 = vout_peek_1361;
    endcase
  endfunction
  wire [7:0] v_10662;
  function [7:0] mux_10662(input [0:0] sel);
    case (sel) 0: mux_10662 = 8'h0; 1: mux_10662 = v_10663;
    endcase
  endfunction
  reg [7:0] v_10663 = 8'h0;
  wire [7:0] v_10664;
  wire [7:0] v_10665;
  function [7:0] mux_10665(input [0:0] sel);
    case (sel) 0: mux_10665 = 8'h0; 1: mux_10665 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10666;
  wire [7:0] v_10667;
  wire [7:0] v_10668;
  function [7:0] mux_10668(input [0:0] sel);
    case (sel) 0: mux_10668 = 8'h0; 1: mux_10668 = vout_peek_1355;
    endcase
  endfunction
  wire [7:0] v_10669;
  function [7:0] mux_10669(input [0:0] sel);
    case (sel) 0: mux_10669 = 8'h0; 1: mux_10669 = vout_peek_1347;
    endcase
  endfunction
  wire [7:0] v_10670;
  function [7:0] mux_10670(input [0:0] sel);
    case (sel) 0: mux_10670 = 8'h0; 1: mux_10670 = v_10671;
    endcase
  endfunction
  reg [7:0] v_10671 = 8'h0;
  wire [7:0] v_10672;
  wire [7:0] v_10673;
  function [7:0] mux_10673(input [0:0] sel);
    case (sel) 0: mux_10673 = 8'h0; 1: mux_10673 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10674;
  wire [7:0] v_10675;
  wire [7:0] v_10676;
  function [7:0] mux_10676(input [0:0] sel);
    case (sel) 0: mux_10676 = 8'h0; 1: mux_10676 = v_10677;
    endcase
  endfunction
  reg [7:0] v_10677 = 8'h0;
  wire [7:0] v_10678;
  wire [7:0] v_10679;
  function [7:0] mux_10679(input [0:0] sel);
    case (sel) 0: mux_10679 = 8'h0; 1: mux_10679 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10680;
  wire [7:0] v_10681;
  wire [7:0] v_10682;
  function [7:0] mux_10682(input [0:0] sel);
    case (sel) 0: mux_10682 = 8'h0; 1: mux_10682 = v_10683;
    endcase
  endfunction
  reg [7:0] v_10683 = 8'h0;
  wire [7:0] v_10684;
  wire [7:0] v_10685;
  function [7:0] mux_10685(input [0:0] sel);
    case (sel) 0: mux_10685 = 8'h0; 1: mux_10685 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10686;
  wire [7:0] v_10687;
  wire [7:0] v_10688;
  function [7:0] mux_10688(input [0:0] sel);
    case (sel) 0: mux_10688 = 8'h0; 1: mux_10688 = v_10689;
    endcase
  endfunction
  reg [7:0] v_10689 = 8'h0;
  wire [7:0] v_10690;
  wire [7:0] v_10691;
  function [7:0] mux_10691(input [0:0] sel);
    case (sel) 0: mux_10691 = 8'h0; 1: mux_10691 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10692;
  wire [7:0] v_10693;
  wire [7:0] v_10694;
  function [7:0] mux_10694(input [0:0] sel);
    case (sel) 0: mux_10694 = 8'h0; 1: mux_10694 = v_10695;
    endcase
  endfunction
  reg [7:0] v_10695 = 8'h0;
  wire [7:0] v_10696;
  wire [7:0] v_10697;
  function [7:0] mux_10697(input [0:0] sel);
    case (sel) 0: mux_10697 = 8'h0; 1: mux_10697 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10698;
  wire [7:0] v_10699;
  wire [7:0] v_10700;
  function [7:0] mux_10700(input [0:0] sel);
    case (sel) 0: mux_10700 = 8'h0; 1: mux_10700 = vout_peek_1341;
    endcase
  endfunction
  wire [7:0] v_10701;
  function [7:0] mux_10701(input [0:0] sel);
    case (sel) 0: mux_10701 = 8'h0; 1: mux_10701 = vout_peek_1333;
    endcase
  endfunction
  wire [7:0] v_10702;
  function [7:0] mux_10702(input [0:0] sel);
    case (sel) 0: mux_10702 = 8'h0; 1: mux_10702 = v_10703;
    endcase
  endfunction
  reg [7:0] v_10703 = 8'h0;
  wire [7:0] v_10704;
  wire [7:0] v_10705;
  function [7:0] mux_10705(input [0:0] sel);
    case (sel) 0: mux_10705 = 8'h0; 1: mux_10705 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10706;
  wire [7:0] v_10707;
  wire [7:0] v_10708;
  function [7:0] mux_10708(input [0:0] sel);
    case (sel) 0: mux_10708 = 8'h0; 1: mux_10708 = vout_peek_1327;
    endcase
  endfunction
  wire [7:0] v_10709;
  function [7:0] mux_10709(input [0:0] sel);
    case (sel) 0: mux_10709 = 8'h0; 1: mux_10709 = vout_peek_1319;
    endcase
  endfunction
  wire [7:0] v_10710;
  function [7:0] mux_10710(input [0:0] sel);
    case (sel) 0: mux_10710 = 8'h0; 1: mux_10710 = v_10711;
    endcase
  endfunction
  reg [7:0] v_10711 = 8'h0;
  wire [7:0] v_10712;
  wire [7:0] v_10713;
  function [7:0] mux_10713(input [0:0] sel);
    case (sel) 0: mux_10713 = 8'h0; 1: mux_10713 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10714;
  wire [7:0] v_10715;
  wire [7:0] v_10716;
  function [7:0] mux_10716(input [0:0] sel);
    case (sel) 0: mux_10716 = 8'h0; 1: mux_10716 = v_10717;
    endcase
  endfunction
  reg [7:0] v_10717 = 8'h0;
  wire [7:0] v_10718;
  wire [7:0] v_10719;
  function [7:0] mux_10719(input [0:0] sel);
    case (sel) 0: mux_10719 = 8'h0; 1: mux_10719 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10720;
  wire [7:0] v_10721;
  wire [7:0] v_10722;
  function [7:0] mux_10722(input [0:0] sel);
    case (sel) 0: mux_10722 = 8'h0; 1: mux_10722 = vout_peek_1313;
    endcase
  endfunction
  wire [7:0] v_10723;
  function [7:0] mux_10723(input [0:0] sel);
    case (sel) 0: mux_10723 = 8'h0; 1: mux_10723 = vout_peek_1305;
    endcase
  endfunction
  wire [7:0] v_10724;
  function [7:0] mux_10724(input [0:0] sel);
    case (sel) 0: mux_10724 = 8'h0; 1: mux_10724 = v_10725;
    endcase
  endfunction
  reg [7:0] v_10725 = 8'h0;
  wire [7:0] v_10726;
  wire [7:0] v_10727;
  function [7:0] mux_10727(input [0:0] sel);
    case (sel) 0: mux_10727 = 8'h0; 1: mux_10727 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10728;
  wire [7:0] v_10729;
  wire [7:0] v_10730;
  function [7:0] mux_10730(input [0:0] sel);
    case (sel) 0: mux_10730 = 8'h0; 1: mux_10730 = vout_peek_1299;
    endcase
  endfunction
  wire [7:0] v_10731;
  function [7:0] mux_10731(input [0:0] sel);
    case (sel) 0: mux_10731 = 8'h0; 1: mux_10731 = vout_peek_1291;
    endcase
  endfunction
  wire [7:0] v_10732;
  function [7:0] mux_10732(input [0:0] sel);
    case (sel) 0: mux_10732 = 8'h0; 1: mux_10732 = v_10733;
    endcase
  endfunction
  reg [7:0] v_10733 = 8'h0;
  wire [7:0] v_10734;
  wire [7:0] v_10735;
  function [7:0] mux_10735(input [0:0] sel);
    case (sel) 0: mux_10735 = 8'h0; 1: mux_10735 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10736;
  wire [7:0] v_10737;
  wire [7:0] v_10738;
  function [7:0] mux_10738(input [0:0] sel);
    case (sel) 0: mux_10738 = 8'h0; 1: mux_10738 = v_10739;
    endcase
  endfunction
  reg [7:0] v_10739 = 8'h0;
  wire [7:0] v_10740;
  wire [7:0] v_10741;
  function [7:0] mux_10741(input [0:0] sel);
    case (sel) 0: mux_10741 = 8'h0; 1: mux_10741 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10742;
  wire [7:0] v_10743;
  wire [7:0] v_10744;
  function [7:0] mux_10744(input [0:0] sel);
    case (sel) 0: mux_10744 = 8'h0; 1: mux_10744 = v_10745;
    endcase
  endfunction
  reg [7:0] v_10745 = 8'h0;
  wire [7:0] v_10746;
  wire [7:0] v_10747;
  function [7:0] mux_10747(input [0:0] sel);
    case (sel) 0: mux_10747 = 8'h0; 1: mux_10747 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10748;
  wire [7:0] v_10749;
  wire [7:0] v_10750;
  function [7:0] mux_10750(input [0:0] sel);
    case (sel) 0: mux_10750 = 8'h0; 1: mux_10750 = vout_peek_1285;
    endcase
  endfunction
  wire [7:0] v_10751;
  function [7:0] mux_10751(input [0:0] sel);
    case (sel) 0: mux_10751 = 8'h0; 1: mux_10751 = vout_peek_1277;
    endcase
  endfunction
  wire [7:0] v_10752;
  function [7:0] mux_10752(input [0:0] sel);
    case (sel) 0: mux_10752 = 8'h0; 1: mux_10752 = v_10753;
    endcase
  endfunction
  reg [7:0] v_10753 = 8'h0;
  wire [7:0] v_10754;
  wire [7:0] v_10755;
  function [7:0] mux_10755(input [0:0] sel);
    case (sel) 0: mux_10755 = 8'h0; 1: mux_10755 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10756;
  wire [7:0] v_10757;
  wire [7:0] v_10758;
  function [7:0] mux_10758(input [0:0] sel);
    case (sel) 0: mux_10758 = 8'h0; 1: mux_10758 = vout_peek_1271;
    endcase
  endfunction
  wire [7:0] v_10759;
  function [7:0] mux_10759(input [0:0] sel);
    case (sel) 0: mux_10759 = 8'h0; 1: mux_10759 = vout_peek_1263;
    endcase
  endfunction
  wire [7:0] v_10760;
  function [7:0] mux_10760(input [0:0] sel);
    case (sel) 0: mux_10760 = 8'h0; 1: mux_10760 = v_10761;
    endcase
  endfunction
  reg [7:0] v_10761 = 8'h0;
  wire [7:0] v_10762;
  wire [7:0] v_10763;
  function [7:0] mux_10763(input [0:0] sel);
    case (sel) 0: mux_10763 = 8'h0; 1: mux_10763 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10764;
  wire [7:0] v_10765;
  wire [7:0] v_10766;
  function [7:0] mux_10766(input [0:0] sel);
    case (sel) 0: mux_10766 = 8'h0; 1: mux_10766 = v_10767;
    endcase
  endfunction
  reg [7:0] v_10767 = 8'h0;
  wire [7:0] v_10768;
  wire [7:0] v_10769;
  function [7:0] mux_10769(input [0:0] sel);
    case (sel) 0: mux_10769 = 8'h0; 1: mux_10769 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10770;
  wire [7:0] v_10771;
  wire [7:0] v_10772;
  function [7:0] mux_10772(input [0:0] sel);
    case (sel) 0: mux_10772 = 8'h0; 1: mux_10772 = vout_peek_1257;
    endcase
  endfunction
  wire [7:0] v_10773;
  function [7:0] mux_10773(input [0:0] sel);
    case (sel) 0: mux_10773 = 8'h0; 1: mux_10773 = vout_peek_1249;
    endcase
  endfunction
  wire [7:0] v_10774;
  function [7:0] mux_10774(input [0:0] sel);
    case (sel) 0: mux_10774 = 8'h0; 1: mux_10774 = v_10775;
    endcase
  endfunction
  reg [7:0] v_10775 = 8'h0;
  wire [7:0] v_10776;
  wire [7:0] v_10777;
  function [7:0] mux_10777(input [0:0] sel);
    case (sel) 0: mux_10777 = 8'h0; 1: mux_10777 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10778;
  wire [7:0] v_10779;
  wire [7:0] v_10780;
  function [7:0] mux_10780(input [0:0] sel);
    case (sel) 0: mux_10780 = 8'h0; 1: mux_10780 = vout_peek_1243;
    endcase
  endfunction
  wire [7:0] v_10781;
  function [7:0] mux_10781(input [0:0] sel);
    case (sel) 0: mux_10781 = 8'h0; 1: mux_10781 = vout_peek_1235;
    endcase
  endfunction
  wire [7:0] v_10782;
  function [7:0] mux_10782(input [0:0] sel);
    case (sel) 0: mux_10782 = 8'h0; 1: mux_10782 = v_10783;
    endcase
  endfunction
  reg [7:0] v_10783 = 8'h0;
  wire [7:0] v_10784;
  wire [7:0] v_10785;
  function [7:0] mux_10785(input [0:0] sel);
    case (sel) 0: mux_10785 = 8'h0; 1: mux_10785 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10786;
  wire [7:0] v_10787;
  wire [7:0] v_10788;
  function [7:0] mux_10788(input [0:0] sel);
    case (sel) 0: mux_10788 = 8'h0; 1: mux_10788 = v_10789;
    endcase
  endfunction
  reg [7:0] v_10789 = 8'h0;
  wire [7:0] v_10790;
  wire [7:0] v_10791;
  function [7:0] mux_10791(input [0:0] sel);
    case (sel) 0: mux_10791 = 8'h0; 1: mux_10791 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10792;
  wire [7:0] v_10793;
  wire [7:0] v_10794;
  function [7:0] mux_10794(input [0:0] sel);
    case (sel) 0: mux_10794 = 8'h0; 1: mux_10794 = v_10795;
    endcase
  endfunction
  reg [7:0] v_10795 = 8'h0;
  wire [7:0] v_10796;
  wire [7:0] v_10797;
  function [7:0] mux_10797(input [0:0] sel);
    case (sel) 0: mux_10797 = 8'h0; 1: mux_10797 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10798;
  wire [7:0] v_10799;
  wire [7:0] v_10800;
  function [7:0] mux_10800(input [0:0] sel);
    case (sel) 0: mux_10800 = 8'h0; 1: mux_10800 = v_10801;
    endcase
  endfunction
  reg [7:0] v_10801 = 8'h0;
  wire [7:0] v_10802;
  wire [7:0] v_10803;
  function [7:0] mux_10803(input [0:0] sel);
    case (sel) 0: mux_10803 = 8'h0; 1: mux_10803 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10804;
  wire [7:0] v_10805;
  wire [7:0] v_10806;
  function [7:0] mux_10806(input [0:0] sel);
    case (sel) 0: mux_10806 = 8'h0; 1: mux_10806 = vout_peek_1229;
    endcase
  endfunction
  wire [7:0] v_10807;
  function [7:0] mux_10807(input [0:0] sel);
    case (sel) 0: mux_10807 = 8'h0; 1: mux_10807 = vout_peek_1221;
    endcase
  endfunction
  wire [7:0] v_10808;
  function [7:0] mux_10808(input [0:0] sel);
    case (sel) 0: mux_10808 = 8'h0; 1: mux_10808 = v_10809;
    endcase
  endfunction
  reg [7:0] v_10809 = 8'h0;
  wire [7:0] v_10810;
  wire [7:0] v_10811;
  function [7:0] mux_10811(input [0:0] sel);
    case (sel) 0: mux_10811 = 8'h0; 1: mux_10811 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10812;
  wire [7:0] v_10813;
  wire [7:0] v_10814;
  function [7:0] mux_10814(input [0:0] sel);
    case (sel) 0: mux_10814 = 8'h0; 1: mux_10814 = vout_peek_1215;
    endcase
  endfunction
  wire [7:0] v_10815;
  function [7:0] mux_10815(input [0:0] sel);
    case (sel) 0: mux_10815 = 8'h0; 1: mux_10815 = vout_peek_1207;
    endcase
  endfunction
  wire [7:0] v_10816;
  function [7:0] mux_10816(input [0:0] sel);
    case (sel) 0: mux_10816 = 8'h0; 1: mux_10816 = v_10817;
    endcase
  endfunction
  reg [7:0] v_10817 = 8'h0;
  wire [7:0] v_10818;
  wire [7:0] v_10819;
  function [7:0] mux_10819(input [0:0] sel);
    case (sel) 0: mux_10819 = 8'h0; 1: mux_10819 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10820;
  wire [7:0] v_10821;
  wire [7:0] v_10822;
  function [7:0] mux_10822(input [0:0] sel);
    case (sel) 0: mux_10822 = 8'h0; 1: mux_10822 = v_10823;
    endcase
  endfunction
  reg [7:0] v_10823 = 8'h0;
  wire [7:0] v_10824;
  wire [7:0] v_10825;
  function [7:0] mux_10825(input [0:0] sel);
    case (sel) 0: mux_10825 = 8'h0; 1: mux_10825 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10826;
  wire [7:0] v_10827;
  wire [7:0] v_10828;
  function [7:0] mux_10828(input [0:0] sel);
    case (sel) 0: mux_10828 = 8'h0; 1: mux_10828 = vout_peek_1201;
    endcase
  endfunction
  wire [7:0] v_10829;
  function [7:0] mux_10829(input [0:0] sel);
    case (sel) 0: mux_10829 = 8'h0; 1: mux_10829 = vout_peek_1193;
    endcase
  endfunction
  wire [7:0] v_10830;
  function [7:0] mux_10830(input [0:0] sel);
    case (sel) 0: mux_10830 = 8'h0; 1: mux_10830 = v_10831;
    endcase
  endfunction
  reg [7:0] v_10831 = 8'h0;
  wire [7:0] v_10832;
  wire [7:0] v_10833;
  function [7:0] mux_10833(input [0:0] sel);
    case (sel) 0: mux_10833 = 8'h0; 1: mux_10833 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10834;
  wire [7:0] v_10835;
  wire [7:0] v_10836;
  function [7:0] mux_10836(input [0:0] sel);
    case (sel) 0: mux_10836 = 8'h0; 1: mux_10836 = vout_peek_1187;
    endcase
  endfunction
  wire [7:0] v_10837;
  function [7:0] mux_10837(input [0:0] sel);
    case (sel) 0: mux_10837 = 8'h0; 1: mux_10837 = vout_peek_1179;
    endcase
  endfunction
  wire [7:0] v_10838;
  function [7:0] mux_10838(input [0:0] sel);
    case (sel) 0: mux_10838 = 8'h0; 1: mux_10838 = v_10839;
    endcase
  endfunction
  reg [7:0] v_10839 = 8'h0;
  wire [7:0] v_10840;
  wire [7:0] v_10841;
  function [7:0] mux_10841(input [0:0] sel);
    case (sel) 0: mux_10841 = 8'h0; 1: mux_10841 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10842;
  wire [7:0] v_10843;
  wire [7:0] v_10844;
  function [7:0] mux_10844(input [0:0] sel);
    case (sel) 0: mux_10844 = 8'h0; 1: mux_10844 = v_10845;
    endcase
  endfunction
  reg [7:0] v_10845 = 8'h0;
  wire [7:0] v_10846;
  wire [7:0] v_10847;
  function [7:0] mux_10847(input [0:0] sel);
    case (sel) 0: mux_10847 = 8'h0; 1: mux_10847 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10848;
  wire [7:0] v_10849;
  wire [7:0] v_10850;
  function [7:0] mux_10850(input [0:0] sel);
    case (sel) 0: mux_10850 = 8'h0; 1: mux_10850 = v_10851;
    endcase
  endfunction
  reg [7:0] v_10851 = 8'h0;
  wire [7:0] v_10852;
  wire [7:0] v_10853;
  function [7:0] mux_10853(input [0:0] sel);
    case (sel) 0: mux_10853 = 8'h0; 1: mux_10853 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10854;
  wire [7:0] v_10855;
  wire [7:0] v_10856;
  function [7:0] mux_10856(input [0:0] sel);
    case (sel) 0: mux_10856 = 8'h0; 1: mux_10856 = vout_peek_1173;
    endcase
  endfunction
  wire [7:0] v_10857;
  function [7:0] mux_10857(input [0:0] sel);
    case (sel) 0: mux_10857 = 8'h0; 1: mux_10857 = vout_peek_1165;
    endcase
  endfunction
  wire [7:0] v_10858;
  function [7:0] mux_10858(input [0:0] sel);
    case (sel) 0: mux_10858 = 8'h0; 1: mux_10858 = v_10859;
    endcase
  endfunction
  reg [7:0] v_10859 = 8'h0;
  wire [7:0] v_10860;
  wire [7:0] v_10861;
  function [7:0] mux_10861(input [0:0] sel);
    case (sel) 0: mux_10861 = 8'h0; 1: mux_10861 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10862;
  wire [7:0] v_10863;
  wire [7:0] v_10864;
  function [7:0] mux_10864(input [0:0] sel);
    case (sel) 0: mux_10864 = 8'h0; 1: mux_10864 = vout_peek_1159;
    endcase
  endfunction
  wire [7:0] v_10865;
  function [7:0] mux_10865(input [0:0] sel);
    case (sel) 0: mux_10865 = 8'h0; 1: mux_10865 = vout_peek_1151;
    endcase
  endfunction
  wire [7:0] v_10866;
  function [7:0] mux_10866(input [0:0] sel);
    case (sel) 0: mux_10866 = 8'h0; 1: mux_10866 = v_10867;
    endcase
  endfunction
  reg [7:0] v_10867 = 8'h0;
  wire [7:0] v_10868;
  wire [7:0] v_10869;
  function [7:0] mux_10869(input [0:0] sel);
    case (sel) 0: mux_10869 = 8'h0; 1: mux_10869 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10870;
  wire [7:0] v_10871;
  wire [7:0] v_10872;
  function [7:0] mux_10872(input [0:0] sel);
    case (sel) 0: mux_10872 = 8'h0; 1: mux_10872 = v_10873;
    endcase
  endfunction
  reg [7:0] v_10873 = 8'h0;
  wire [7:0] v_10874;
  wire [7:0] v_10875;
  function [7:0] mux_10875(input [0:0] sel);
    case (sel) 0: mux_10875 = 8'h0; 1: mux_10875 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10876;
  wire [7:0] v_10877;
  wire [7:0] v_10878;
  function [7:0] mux_10878(input [0:0] sel);
    case (sel) 0: mux_10878 = 8'h0; 1: mux_10878 = vout_peek_1145;
    endcase
  endfunction
  wire [7:0] v_10879;
  function [7:0] mux_10879(input [0:0] sel);
    case (sel) 0: mux_10879 = 8'h0; 1: mux_10879 = vout_peek_1137;
    endcase
  endfunction
  wire [7:0] v_10880;
  function [7:0] mux_10880(input [0:0] sel);
    case (sel) 0: mux_10880 = 8'h0; 1: mux_10880 = v_10881;
    endcase
  endfunction
  reg [7:0] v_10881 = 8'h0;
  wire [7:0] v_10882;
  wire [7:0] v_10883;
  function [7:0] mux_10883(input [0:0] sel);
    case (sel) 0: mux_10883 = 8'h0; 1: mux_10883 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10884;
  wire [7:0] v_10885;
  wire [7:0] v_10886;
  function [7:0] mux_10886(input [0:0] sel);
    case (sel) 0: mux_10886 = 8'h0; 1: mux_10886 = vout_peek_1131;
    endcase
  endfunction
  wire [7:0] v_10887;
  function [7:0] mux_10887(input [0:0] sel);
    case (sel) 0: mux_10887 = 8'h0; 1: mux_10887 = vout_peek_1123;
    endcase
  endfunction
  wire [7:0] v_10888;
  function [7:0] mux_10888(input [0:0] sel);
    case (sel) 0: mux_10888 = 8'h0; 1: mux_10888 = v_10889;
    endcase
  endfunction
  reg [7:0] v_10889 = 8'h0;
  wire [7:0] v_10890;
  wire [7:0] v_10891;
  function [7:0] mux_10891(input [0:0] sel);
    case (sel) 0: mux_10891 = 8'h0; 1: mux_10891 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10892;
  wire [7:0] v_10893;
  wire [7:0] v_10894;
  function [7:0] mux_10894(input [0:0] sel);
    case (sel) 0: mux_10894 = 8'h0; 1: mux_10894 = v_10895;
    endcase
  endfunction
  reg [7:0] v_10895 = 8'h0;
  wire [7:0] v_10896;
  wire [7:0] v_10897;
  function [7:0] mux_10897(input [0:0] sel);
    case (sel) 0: mux_10897 = 8'h0; 1: mux_10897 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10898;
  wire [7:0] v_10899;
  wire [7:0] v_10900;
  function [7:0] mux_10900(input [0:0] sel);
    case (sel) 0: mux_10900 = 8'h0; 1: mux_10900 = v_10901;
    endcase
  endfunction
  reg [7:0] v_10901 = 8'h0;
  wire [7:0] v_10902;
  wire [7:0] v_10903;
  function [7:0] mux_10903(input [0:0] sel);
    case (sel) 0: mux_10903 = 8'h0; 1: mux_10903 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10904;
  wire [7:0] v_10905;
  wire [7:0] v_10906;
  function [7:0] mux_10906(input [0:0] sel);
    case (sel) 0: mux_10906 = 8'h0; 1: mux_10906 = v_10907;
    endcase
  endfunction
  reg [7:0] v_10907 = 8'h0;
  wire [7:0] v_10908;
  wire [7:0] v_10909;
  function [7:0] mux_10909(input [0:0] sel);
    case (sel) 0: mux_10909 = 8'h0; 1: mux_10909 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10910;
  wire [7:0] v_10911;
  wire [7:0] v_10912;
  function [7:0] mux_10912(input [0:0] sel);
    case (sel) 0: mux_10912 = 8'h0; 1: mux_10912 = v_10913;
    endcase
  endfunction
  reg [7:0] v_10913 = 8'h0;
  wire [7:0] v_10914;
  wire [7:0] v_10915;
  function [7:0] mux_10915(input [0:0] sel);
    case (sel) 0: mux_10915 = 8'h0; 1: mux_10915 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10916;
  wire [7:0] v_10917;
  wire [7:0] v_10918;
  function [7:0] mux_10918(input [0:0] sel);
    case (sel) 0: mux_10918 = 8'h0; 1: mux_10918 = v_10919;
    endcase
  endfunction
  reg [7:0] v_10919 = 8'h0;
  wire [7:0] v_10920;
  wire [7:0] v_10921;
  function [7:0] mux_10921(input [0:0] sel);
    case (sel) 0: mux_10921 = 8'h0; 1: mux_10921 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10922;
  wire [7:0] v_10923;
  wire [7:0] v_10924;
  function [7:0] mux_10924(input [0:0] sel);
    case (sel) 0: mux_10924 = 8'h0; 1: mux_10924 = v_10925;
    endcase
  endfunction
  reg [7:0] v_10925 = 8'h0;
  wire [7:0] v_10926;
  wire [7:0] v_10927;
  function [7:0] mux_10927(input [0:0] sel);
    case (sel) 0: mux_10927 = 8'h0; 1: mux_10927 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10928;
  wire [7:0] v_10929;
  wire [7:0] v_10930;
  function [7:0] mux_10930(input [0:0] sel);
    case (sel) 0: mux_10930 = 8'h0; 1: mux_10930 = vout_peek_1117;
    endcase
  endfunction
  wire [7:0] v_10931;
  function [7:0] mux_10931(input [0:0] sel);
    case (sel) 0: mux_10931 = 8'h0; 1: mux_10931 = vout_peek_1109;
    endcase
  endfunction
  wire [7:0] v_10932;
  function [7:0] mux_10932(input [0:0] sel);
    case (sel) 0: mux_10932 = 8'h0; 1: mux_10932 = v_10933;
    endcase
  endfunction
  reg [7:0] v_10933 = 8'h0;
  wire [7:0] v_10934;
  wire [7:0] v_10935;
  function [7:0] mux_10935(input [0:0] sel);
    case (sel) 0: mux_10935 = 8'h0; 1: mux_10935 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10936;
  wire [7:0] v_10937;
  wire [7:0] v_10938;
  function [7:0] mux_10938(input [0:0] sel);
    case (sel) 0: mux_10938 = 8'h0; 1: mux_10938 = vout_peek_1103;
    endcase
  endfunction
  wire [7:0] v_10939;
  function [7:0] mux_10939(input [0:0] sel);
    case (sel) 0: mux_10939 = 8'h0; 1: mux_10939 = vout_peek_1095;
    endcase
  endfunction
  wire [7:0] v_10940;
  function [7:0] mux_10940(input [0:0] sel);
    case (sel) 0: mux_10940 = 8'h0; 1: mux_10940 = v_10941;
    endcase
  endfunction
  reg [7:0] v_10941 = 8'h0;
  wire [7:0] v_10942;
  wire [7:0] v_10943;
  function [7:0] mux_10943(input [0:0] sel);
    case (sel) 0: mux_10943 = 8'h0; 1: mux_10943 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10944;
  wire [7:0] v_10945;
  wire [7:0] v_10946;
  function [7:0] mux_10946(input [0:0] sel);
    case (sel) 0: mux_10946 = 8'h0; 1: mux_10946 = v_10947;
    endcase
  endfunction
  reg [7:0] v_10947 = 8'h0;
  wire [7:0] v_10948;
  wire [7:0] v_10949;
  function [7:0] mux_10949(input [0:0] sel);
    case (sel) 0: mux_10949 = 8'h0; 1: mux_10949 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10950;
  wire [7:0] v_10951;
  wire [7:0] v_10952;
  function [7:0] mux_10952(input [0:0] sel);
    case (sel) 0: mux_10952 = 8'h0; 1: mux_10952 = vout_peek_1089;
    endcase
  endfunction
  wire [7:0] v_10953;
  function [7:0] mux_10953(input [0:0] sel);
    case (sel) 0: mux_10953 = 8'h0; 1: mux_10953 = vout_peek_1081;
    endcase
  endfunction
  wire [7:0] v_10954;
  function [7:0] mux_10954(input [0:0] sel);
    case (sel) 0: mux_10954 = 8'h0; 1: mux_10954 = v_10955;
    endcase
  endfunction
  reg [7:0] v_10955 = 8'h0;
  wire [7:0] v_10956;
  wire [7:0] v_10957;
  function [7:0] mux_10957(input [0:0] sel);
    case (sel) 0: mux_10957 = 8'h0; 1: mux_10957 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10958;
  wire [7:0] v_10959;
  wire [7:0] v_10960;
  function [7:0] mux_10960(input [0:0] sel);
    case (sel) 0: mux_10960 = 8'h0; 1: mux_10960 = vout_peek_1075;
    endcase
  endfunction
  wire [7:0] v_10961;
  function [7:0] mux_10961(input [0:0] sel);
    case (sel) 0: mux_10961 = 8'h0; 1: mux_10961 = vout_peek_1067;
    endcase
  endfunction
  wire [7:0] v_10962;
  function [7:0] mux_10962(input [0:0] sel);
    case (sel) 0: mux_10962 = 8'h0; 1: mux_10962 = v_10963;
    endcase
  endfunction
  reg [7:0] v_10963 = 8'h0;
  wire [7:0] v_10964;
  wire [7:0] v_10965;
  function [7:0] mux_10965(input [0:0] sel);
    case (sel) 0: mux_10965 = 8'h0; 1: mux_10965 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10966;
  wire [7:0] v_10967;
  wire [7:0] v_10968;
  function [7:0] mux_10968(input [0:0] sel);
    case (sel) 0: mux_10968 = 8'h0; 1: mux_10968 = v_10969;
    endcase
  endfunction
  reg [7:0] v_10969 = 8'h0;
  wire [7:0] v_10970;
  wire [7:0] v_10971;
  function [7:0] mux_10971(input [0:0] sel);
    case (sel) 0: mux_10971 = 8'h0; 1: mux_10971 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10972;
  wire [7:0] v_10973;
  wire [7:0] v_10974;
  function [7:0] mux_10974(input [0:0] sel);
    case (sel) 0: mux_10974 = 8'h0; 1: mux_10974 = v_10975;
    endcase
  endfunction
  reg [7:0] v_10975 = 8'h0;
  wire [7:0] v_10976;
  wire [7:0] v_10977;
  function [7:0] mux_10977(input [0:0] sel);
    case (sel) 0: mux_10977 = 8'h0; 1: mux_10977 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10978;
  wire [7:0] v_10979;
  wire [7:0] v_10980;
  function [7:0] mux_10980(input [0:0] sel);
    case (sel) 0: mux_10980 = 8'h0; 1: mux_10980 = vout_peek_1061;
    endcase
  endfunction
  wire [7:0] v_10981;
  function [7:0] mux_10981(input [0:0] sel);
    case (sel) 0: mux_10981 = 8'h0; 1: mux_10981 = vout_peek_1053;
    endcase
  endfunction
  wire [7:0] v_10982;
  function [7:0] mux_10982(input [0:0] sel);
    case (sel) 0: mux_10982 = 8'h0; 1: mux_10982 = v_10983;
    endcase
  endfunction
  reg [7:0] v_10983 = 8'h0;
  wire [7:0] v_10984;
  wire [7:0] v_10985;
  function [7:0] mux_10985(input [0:0] sel);
    case (sel) 0: mux_10985 = 8'h0; 1: mux_10985 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10986;
  wire [7:0] v_10987;
  wire [7:0] v_10988;
  function [7:0] mux_10988(input [0:0] sel);
    case (sel) 0: mux_10988 = 8'h0; 1: mux_10988 = vout_peek_1047;
    endcase
  endfunction
  wire [7:0] v_10989;
  function [7:0] mux_10989(input [0:0] sel);
    case (sel) 0: mux_10989 = 8'h0; 1: mux_10989 = vout_peek_1039;
    endcase
  endfunction
  wire [7:0] v_10990;
  function [7:0] mux_10990(input [0:0] sel);
    case (sel) 0: mux_10990 = 8'h0; 1: mux_10990 = v_10991;
    endcase
  endfunction
  reg [7:0] v_10991 = 8'h0;
  wire [7:0] v_10992;
  wire [7:0] v_10993;
  function [7:0] mux_10993(input [0:0] sel);
    case (sel) 0: mux_10993 = 8'h0; 1: mux_10993 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_10994;
  wire [7:0] v_10995;
  wire [7:0] v_10996;
  function [7:0] mux_10996(input [0:0] sel);
    case (sel) 0: mux_10996 = 8'h0; 1: mux_10996 = v_10997;
    endcase
  endfunction
  reg [7:0] v_10997 = 8'h0;
  wire [7:0] v_10998;
  wire [7:0] v_10999;
  function [7:0] mux_10999(input [0:0] sel);
    case (sel) 0: mux_10999 = 8'h0; 1: mux_10999 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11000;
  wire [7:0] v_11001;
  wire [7:0] v_11002;
  function [7:0] mux_11002(input [0:0] sel);
    case (sel) 0: mux_11002 = 8'h0; 1: mux_11002 = vout_peek_1033;
    endcase
  endfunction
  wire [7:0] v_11003;
  function [7:0] mux_11003(input [0:0] sel);
    case (sel) 0: mux_11003 = 8'h0; 1: mux_11003 = vout_peek_1025;
    endcase
  endfunction
  wire [7:0] v_11004;
  function [7:0] mux_11004(input [0:0] sel);
    case (sel) 0: mux_11004 = 8'h0; 1: mux_11004 = v_11005;
    endcase
  endfunction
  reg [7:0] v_11005 = 8'h0;
  wire [7:0] v_11006;
  wire [7:0] v_11007;
  function [7:0] mux_11007(input [0:0] sel);
    case (sel) 0: mux_11007 = 8'h0; 1: mux_11007 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11008;
  wire [7:0] v_11009;
  wire [7:0] v_11010;
  function [7:0] mux_11010(input [0:0] sel);
    case (sel) 0: mux_11010 = 8'h0; 1: mux_11010 = vout_peek_1019;
    endcase
  endfunction
  wire [7:0] v_11011;
  function [7:0] mux_11011(input [0:0] sel);
    case (sel) 0: mux_11011 = 8'h0; 1: mux_11011 = vout_peek_1011;
    endcase
  endfunction
  wire [7:0] v_11012;
  function [7:0] mux_11012(input [0:0] sel);
    case (sel) 0: mux_11012 = 8'h0; 1: mux_11012 = v_11013;
    endcase
  endfunction
  reg [7:0] v_11013 = 8'h0;
  wire [7:0] v_11014;
  wire [7:0] v_11015;
  function [7:0] mux_11015(input [0:0] sel);
    case (sel) 0: mux_11015 = 8'h0; 1: mux_11015 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11016;
  wire [7:0] v_11017;
  wire [7:0] v_11018;
  function [7:0] mux_11018(input [0:0] sel);
    case (sel) 0: mux_11018 = 8'h0; 1: mux_11018 = v_11019;
    endcase
  endfunction
  reg [7:0] v_11019 = 8'h0;
  wire [7:0] v_11020;
  wire [7:0] v_11021;
  function [7:0] mux_11021(input [0:0] sel);
    case (sel) 0: mux_11021 = 8'h0; 1: mux_11021 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11022;
  wire [7:0] v_11023;
  wire [7:0] v_11024;
  function [7:0] mux_11024(input [0:0] sel);
    case (sel) 0: mux_11024 = 8'h0; 1: mux_11024 = v_11025;
    endcase
  endfunction
  reg [7:0] v_11025 = 8'h0;
  wire [7:0] v_11026;
  wire [7:0] v_11027;
  function [7:0] mux_11027(input [0:0] sel);
    case (sel) 0: mux_11027 = 8'h0; 1: mux_11027 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11028;
  wire [7:0] v_11029;
  wire [7:0] v_11030;
  function [7:0] mux_11030(input [0:0] sel);
    case (sel) 0: mux_11030 = 8'h0; 1: mux_11030 = v_11031;
    endcase
  endfunction
  reg [7:0] v_11031 = 8'h0;
  wire [7:0] v_11032;
  wire [7:0] v_11033;
  function [7:0] mux_11033(input [0:0] sel);
    case (sel) 0: mux_11033 = 8'h0; 1: mux_11033 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11034;
  wire [7:0] v_11035;
  wire [7:0] v_11036;
  function [7:0] mux_11036(input [0:0] sel);
    case (sel) 0: mux_11036 = 8'h0; 1: mux_11036 = vout_peek_1005;
    endcase
  endfunction
  wire [7:0] v_11037;
  function [7:0] mux_11037(input [0:0] sel);
    case (sel) 0: mux_11037 = 8'h0; 1: mux_11037 = vout_peek_997;
    endcase
  endfunction
  wire [7:0] v_11038;
  function [7:0] mux_11038(input [0:0] sel);
    case (sel) 0: mux_11038 = 8'h0; 1: mux_11038 = v_11039;
    endcase
  endfunction
  reg [7:0] v_11039 = 8'h0;
  wire [7:0] v_11040;
  wire [7:0] v_11041;
  function [7:0] mux_11041(input [0:0] sel);
    case (sel) 0: mux_11041 = 8'h0; 1: mux_11041 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11042;
  wire [7:0] v_11043;
  wire [7:0] v_11044;
  function [7:0] mux_11044(input [0:0] sel);
    case (sel) 0: mux_11044 = 8'h0; 1: mux_11044 = vout_peek_991;
    endcase
  endfunction
  wire [7:0] v_11045;
  function [7:0] mux_11045(input [0:0] sel);
    case (sel) 0: mux_11045 = 8'h0; 1: mux_11045 = vout_peek_983;
    endcase
  endfunction
  wire [7:0] v_11046;
  function [7:0] mux_11046(input [0:0] sel);
    case (sel) 0: mux_11046 = 8'h0; 1: mux_11046 = v_11047;
    endcase
  endfunction
  reg [7:0] v_11047 = 8'h0;
  wire [7:0] v_11048;
  wire [7:0] v_11049;
  function [7:0] mux_11049(input [0:0] sel);
    case (sel) 0: mux_11049 = 8'h0; 1: mux_11049 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11050;
  wire [7:0] v_11051;
  wire [7:0] v_11052;
  function [7:0] mux_11052(input [0:0] sel);
    case (sel) 0: mux_11052 = 8'h0; 1: mux_11052 = v_11053;
    endcase
  endfunction
  reg [7:0] v_11053 = 8'h0;
  wire [7:0] v_11054;
  wire [7:0] v_11055;
  function [7:0] mux_11055(input [0:0] sel);
    case (sel) 0: mux_11055 = 8'h0; 1: mux_11055 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11056;
  wire [7:0] v_11057;
  wire [7:0] v_11058;
  function [7:0] mux_11058(input [0:0] sel);
    case (sel) 0: mux_11058 = 8'h0; 1: mux_11058 = vout_peek_977;
    endcase
  endfunction
  wire [7:0] v_11059;
  function [7:0] mux_11059(input [0:0] sel);
    case (sel) 0: mux_11059 = 8'h0; 1: mux_11059 = vout_peek_969;
    endcase
  endfunction
  wire [7:0] v_11060;
  function [7:0] mux_11060(input [0:0] sel);
    case (sel) 0: mux_11060 = 8'h0; 1: mux_11060 = v_11061;
    endcase
  endfunction
  reg [7:0] v_11061 = 8'h0;
  wire [7:0] v_11062;
  wire [7:0] v_11063;
  function [7:0] mux_11063(input [0:0] sel);
    case (sel) 0: mux_11063 = 8'h0; 1: mux_11063 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11064;
  wire [7:0] v_11065;
  wire [7:0] v_11066;
  function [7:0] mux_11066(input [0:0] sel);
    case (sel) 0: mux_11066 = 8'h0; 1: mux_11066 = vout_peek_963;
    endcase
  endfunction
  wire [7:0] v_11067;
  function [7:0] mux_11067(input [0:0] sel);
    case (sel) 0: mux_11067 = 8'h0; 1: mux_11067 = vout_peek_955;
    endcase
  endfunction
  wire [7:0] v_11068;
  function [7:0] mux_11068(input [0:0] sel);
    case (sel) 0: mux_11068 = 8'h0; 1: mux_11068 = v_11069;
    endcase
  endfunction
  reg [7:0] v_11069 = 8'h0;
  wire [7:0] v_11070;
  wire [7:0] v_11071;
  function [7:0] mux_11071(input [0:0] sel);
    case (sel) 0: mux_11071 = 8'h0; 1: mux_11071 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11072;
  wire [7:0] v_11073;
  wire [7:0] v_11074;
  function [7:0] mux_11074(input [0:0] sel);
    case (sel) 0: mux_11074 = 8'h0; 1: mux_11074 = v_11075;
    endcase
  endfunction
  reg [7:0] v_11075 = 8'h0;
  wire [7:0] v_11076;
  wire [7:0] v_11077;
  function [7:0] mux_11077(input [0:0] sel);
    case (sel) 0: mux_11077 = 8'h0; 1: mux_11077 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11078;
  wire [7:0] v_11079;
  wire [7:0] v_11080;
  function [7:0] mux_11080(input [0:0] sel);
    case (sel) 0: mux_11080 = 8'h0; 1: mux_11080 = v_11081;
    endcase
  endfunction
  reg [7:0] v_11081 = 8'h0;
  wire [7:0] v_11082;
  wire [7:0] v_11083;
  function [7:0] mux_11083(input [0:0] sel);
    case (sel) 0: mux_11083 = 8'h0; 1: mux_11083 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11084;
  wire [7:0] v_11085;
  wire [7:0] v_11086;
  function [7:0] mux_11086(input [0:0] sel);
    case (sel) 0: mux_11086 = 8'h0; 1: mux_11086 = vout_peek_949;
    endcase
  endfunction
  wire [7:0] v_11087;
  function [7:0] mux_11087(input [0:0] sel);
    case (sel) 0: mux_11087 = 8'h0; 1: mux_11087 = vout_peek_941;
    endcase
  endfunction
  wire [7:0] v_11088;
  function [7:0] mux_11088(input [0:0] sel);
    case (sel) 0: mux_11088 = 8'h0; 1: mux_11088 = v_11089;
    endcase
  endfunction
  reg [7:0] v_11089 = 8'h0;
  wire [7:0] v_11090;
  wire [7:0] v_11091;
  function [7:0] mux_11091(input [0:0] sel);
    case (sel) 0: mux_11091 = 8'h0; 1: mux_11091 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11092;
  wire [7:0] v_11093;
  wire [7:0] v_11094;
  function [7:0] mux_11094(input [0:0] sel);
    case (sel) 0: mux_11094 = 8'h0; 1: mux_11094 = vout_peek_935;
    endcase
  endfunction
  wire [7:0] v_11095;
  function [7:0] mux_11095(input [0:0] sel);
    case (sel) 0: mux_11095 = 8'h0; 1: mux_11095 = vout_peek_927;
    endcase
  endfunction
  wire [7:0] v_11096;
  function [7:0] mux_11096(input [0:0] sel);
    case (sel) 0: mux_11096 = 8'h0; 1: mux_11096 = v_11097;
    endcase
  endfunction
  reg [7:0] v_11097 = 8'h0;
  wire [7:0] v_11098;
  wire [7:0] v_11099;
  function [7:0] mux_11099(input [0:0] sel);
    case (sel) 0: mux_11099 = 8'h0; 1: mux_11099 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11100;
  wire [7:0] v_11101;
  wire [7:0] v_11102;
  function [7:0] mux_11102(input [0:0] sel);
    case (sel) 0: mux_11102 = 8'h0; 1: mux_11102 = v_11103;
    endcase
  endfunction
  reg [7:0] v_11103 = 8'h0;
  wire [7:0] v_11104;
  wire [7:0] v_11105;
  function [7:0] mux_11105(input [0:0] sel);
    case (sel) 0: mux_11105 = 8'h0; 1: mux_11105 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11106;
  wire [7:0] v_11107;
  wire [7:0] v_11108;
  function [7:0] mux_11108(input [0:0] sel);
    case (sel) 0: mux_11108 = 8'h0; 1: mux_11108 = vout_peek_921;
    endcase
  endfunction
  wire [7:0] v_11109;
  function [7:0] mux_11109(input [0:0] sel);
    case (sel) 0: mux_11109 = 8'h0; 1: mux_11109 = vout_peek_913;
    endcase
  endfunction
  wire [7:0] v_11110;
  function [7:0] mux_11110(input [0:0] sel);
    case (sel) 0: mux_11110 = 8'h0; 1: mux_11110 = v_11111;
    endcase
  endfunction
  reg [7:0] v_11111 = 8'h0;
  wire [7:0] v_11112;
  wire [7:0] v_11113;
  function [7:0] mux_11113(input [0:0] sel);
    case (sel) 0: mux_11113 = 8'h0; 1: mux_11113 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11114;
  wire [7:0] v_11115;
  wire [7:0] v_11116;
  function [7:0] mux_11116(input [0:0] sel);
    case (sel) 0: mux_11116 = 8'h0; 1: mux_11116 = vout_peek_907;
    endcase
  endfunction
  wire [7:0] v_11117;
  function [7:0] mux_11117(input [0:0] sel);
    case (sel) 0: mux_11117 = 8'h0; 1: mux_11117 = vout_peek_899;
    endcase
  endfunction
  wire [7:0] v_11118;
  function [7:0] mux_11118(input [0:0] sel);
    case (sel) 0: mux_11118 = 8'h0; 1: mux_11118 = v_11119;
    endcase
  endfunction
  reg [7:0] v_11119 = 8'h0;
  wire [7:0] v_11120;
  wire [7:0] v_11121;
  function [7:0] mux_11121(input [0:0] sel);
    case (sel) 0: mux_11121 = 8'h0; 1: mux_11121 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11122;
  wire [7:0] v_11123;
  wire [7:0] v_11124;
  function [7:0] mux_11124(input [0:0] sel);
    case (sel) 0: mux_11124 = 8'h0; 1: mux_11124 = v_11125;
    endcase
  endfunction
  reg [7:0] v_11125 = 8'h0;
  wire [7:0] v_11126;
  wire [7:0] v_11127;
  function [7:0] mux_11127(input [0:0] sel);
    case (sel) 0: mux_11127 = 8'h0; 1: mux_11127 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11128;
  wire [7:0] v_11129;
  wire [7:0] v_11130;
  function [7:0] mux_11130(input [0:0] sel);
    case (sel) 0: mux_11130 = 8'h0; 1: mux_11130 = v_11131;
    endcase
  endfunction
  reg [7:0] v_11131 = 8'h0;
  wire [7:0] v_11132;
  wire [7:0] v_11133;
  function [7:0] mux_11133(input [0:0] sel);
    case (sel) 0: mux_11133 = 8'h0; 1: mux_11133 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11134;
  wire [7:0] v_11135;
  wire [7:0] v_11136;
  function [7:0] mux_11136(input [0:0] sel);
    case (sel) 0: mux_11136 = 8'h0; 1: mux_11136 = v_11137;
    endcase
  endfunction
  reg [7:0] v_11137 = 8'h0;
  wire [7:0] v_11138;
  wire [7:0] v_11139;
  function [7:0] mux_11139(input [0:0] sel);
    case (sel) 0: mux_11139 = 8'h0; 1: mux_11139 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11140;
  wire [7:0] v_11141;
  wire [7:0] v_11142;
  function [7:0] mux_11142(input [0:0] sel);
    case (sel) 0: mux_11142 = 8'h0; 1: mux_11142 = v_11143;
    endcase
  endfunction
  reg [7:0] v_11143 = 8'h0;
  wire [7:0] v_11144;
  wire [7:0] v_11145;
  function [7:0] mux_11145(input [0:0] sel);
    case (sel) 0: mux_11145 = 8'h0; 1: mux_11145 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11146;
  wire [7:0] v_11147;
  wire [7:0] v_11148;
  function [7:0] mux_11148(input [0:0] sel);
    case (sel) 0: mux_11148 = 8'h0; 1: mux_11148 = vout_peek_893;
    endcase
  endfunction
  wire [7:0] v_11149;
  function [7:0] mux_11149(input [0:0] sel);
    case (sel) 0: mux_11149 = 8'h0; 1: mux_11149 = vout_peek_885;
    endcase
  endfunction
  wire [7:0] v_11150;
  function [7:0] mux_11150(input [0:0] sel);
    case (sel) 0: mux_11150 = 8'h0; 1: mux_11150 = v_11151;
    endcase
  endfunction
  reg [7:0] v_11151 = 8'h0;
  wire [7:0] v_11152;
  wire [7:0] v_11153;
  function [7:0] mux_11153(input [0:0] sel);
    case (sel) 0: mux_11153 = 8'h0; 1: mux_11153 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11154;
  wire [7:0] v_11155;
  wire [7:0] v_11156;
  function [7:0] mux_11156(input [0:0] sel);
    case (sel) 0: mux_11156 = 8'h0; 1: mux_11156 = vout_peek_879;
    endcase
  endfunction
  wire [7:0] v_11157;
  function [7:0] mux_11157(input [0:0] sel);
    case (sel) 0: mux_11157 = 8'h0; 1: mux_11157 = vout_peek_871;
    endcase
  endfunction
  wire [7:0] v_11158;
  function [7:0] mux_11158(input [0:0] sel);
    case (sel) 0: mux_11158 = 8'h0; 1: mux_11158 = v_11159;
    endcase
  endfunction
  reg [7:0] v_11159 = 8'h0;
  wire [7:0] v_11160;
  wire [7:0] v_11161;
  function [7:0] mux_11161(input [0:0] sel);
    case (sel) 0: mux_11161 = 8'h0; 1: mux_11161 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11162;
  wire [7:0] v_11163;
  wire [7:0] v_11164;
  function [7:0] mux_11164(input [0:0] sel);
    case (sel) 0: mux_11164 = 8'h0; 1: mux_11164 = v_11165;
    endcase
  endfunction
  reg [7:0] v_11165 = 8'h0;
  wire [7:0] v_11166;
  wire [7:0] v_11167;
  function [7:0] mux_11167(input [0:0] sel);
    case (sel) 0: mux_11167 = 8'h0; 1: mux_11167 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11168;
  wire [7:0] v_11169;
  wire [7:0] v_11170;
  function [7:0] mux_11170(input [0:0] sel);
    case (sel) 0: mux_11170 = 8'h0; 1: mux_11170 = vout_peek_865;
    endcase
  endfunction
  wire [7:0] v_11171;
  function [7:0] mux_11171(input [0:0] sel);
    case (sel) 0: mux_11171 = 8'h0; 1: mux_11171 = vout_peek_857;
    endcase
  endfunction
  wire [7:0] v_11172;
  function [7:0] mux_11172(input [0:0] sel);
    case (sel) 0: mux_11172 = 8'h0; 1: mux_11172 = v_11173;
    endcase
  endfunction
  reg [7:0] v_11173 = 8'h0;
  wire [7:0] v_11174;
  wire [7:0] v_11175;
  function [7:0] mux_11175(input [0:0] sel);
    case (sel) 0: mux_11175 = 8'h0; 1: mux_11175 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11176;
  wire [7:0] v_11177;
  wire [7:0] v_11178;
  function [7:0] mux_11178(input [0:0] sel);
    case (sel) 0: mux_11178 = 8'h0; 1: mux_11178 = vout_peek_851;
    endcase
  endfunction
  wire [7:0] v_11179;
  function [7:0] mux_11179(input [0:0] sel);
    case (sel) 0: mux_11179 = 8'h0; 1: mux_11179 = vout_peek_843;
    endcase
  endfunction
  wire [7:0] v_11180;
  function [7:0] mux_11180(input [0:0] sel);
    case (sel) 0: mux_11180 = 8'h0; 1: mux_11180 = v_11181;
    endcase
  endfunction
  reg [7:0] v_11181 = 8'h0;
  wire [7:0] v_11182;
  wire [7:0] v_11183;
  function [7:0] mux_11183(input [0:0] sel);
    case (sel) 0: mux_11183 = 8'h0; 1: mux_11183 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11184;
  wire [7:0] v_11185;
  wire [7:0] v_11186;
  function [7:0] mux_11186(input [0:0] sel);
    case (sel) 0: mux_11186 = 8'h0; 1: mux_11186 = v_11187;
    endcase
  endfunction
  reg [7:0] v_11187 = 8'h0;
  wire [7:0] v_11188;
  wire [7:0] v_11189;
  function [7:0] mux_11189(input [0:0] sel);
    case (sel) 0: mux_11189 = 8'h0; 1: mux_11189 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11190;
  wire [7:0] v_11191;
  wire [7:0] v_11192;
  function [7:0] mux_11192(input [0:0] sel);
    case (sel) 0: mux_11192 = 8'h0; 1: mux_11192 = v_11193;
    endcase
  endfunction
  reg [7:0] v_11193 = 8'h0;
  wire [7:0] v_11194;
  wire [7:0] v_11195;
  function [7:0] mux_11195(input [0:0] sel);
    case (sel) 0: mux_11195 = 8'h0; 1: mux_11195 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11196;
  wire [7:0] v_11197;
  wire [7:0] v_11198;
  function [7:0] mux_11198(input [0:0] sel);
    case (sel) 0: mux_11198 = 8'h0; 1: mux_11198 = vout_peek_837;
    endcase
  endfunction
  wire [7:0] v_11199;
  function [7:0] mux_11199(input [0:0] sel);
    case (sel) 0: mux_11199 = 8'h0; 1: mux_11199 = vout_peek_829;
    endcase
  endfunction
  wire [7:0] v_11200;
  function [7:0] mux_11200(input [0:0] sel);
    case (sel) 0: mux_11200 = 8'h0; 1: mux_11200 = v_11201;
    endcase
  endfunction
  reg [7:0] v_11201 = 8'h0;
  wire [7:0] v_11202;
  wire [7:0] v_11203;
  function [7:0] mux_11203(input [0:0] sel);
    case (sel) 0: mux_11203 = 8'h0; 1: mux_11203 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11204;
  wire [7:0] v_11205;
  wire [7:0] v_11206;
  function [7:0] mux_11206(input [0:0] sel);
    case (sel) 0: mux_11206 = 8'h0; 1: mux_11206 = vout_peek_823;
    endcase
  endfunction
  wire [7:0] v_11207;
  function [7:0] mux_11207(input [0:0] sel);
    case (sel) 0: mux_11207 = 8'h0; 1: mux_11207 = vout_peek_815;
    endcase
  endfunction
  wire [7:0] v_11208;
  function [7:0] mux_11208(input [0:0] sel);
    case (sel) 0: mux_11208 = 8'h0; 1: mux_11208 = v_11209;
    endcase
  endfunction
  reg [7:0] v_11209 = 8'h0;
  wire [7:0] v_11210;
  wire [7:0] v_11211;
  function [7:0] mux_11211(input [0:0] sel);
    case (sel) 0: mux_11211 = 8'h0; 1: mux_11211 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11212;
  wire [7:0] v_11213;
  wire [7:0] v_11214;
  function [7:0] mux_11214(input [0:0] sel);
    case (sel) 0: mux_11214 = 8'h0; 1: mux_11214 = v_11215;
    endcase
  endfunction
  reg [7:0] v_11215 = 8'h0;
  wire [7:0] v_11216;
  wire [7:0] v_11217;
  function [7:0] mux_11217(input [0:0] sel);
    case (sel) 0: mux_11217 = 8'h0; 1: mux_11217 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11218;
  wire [7:0] v_11219;
  wire [7:0] v_11220;
  function [7:0] mux_11220(input [0:0] sel);
    case (sel) 0: mux_11220 = 8'h0; 1: mux_11220 = vout_peek_809;
    endcase
  endfunction
  wire [7:0] v_11221;
  function [7:0] mux_11221(input [0:0] sel);
    case (sel) 0: mux_11221 = 8'h0; 1: mux_11221 = vout_peek_801;
    endcase
  endfunction
  wire [7:0] v_11222;
  function [7:0] mux_11222(input [0:0] sel);
    case (sel) 0: mux_11222 = 8'h0; 1: mux_11222 = v_11223;
    endcase
  endfunction
  reg [7:0] v_11223 = 8'h0;
  wire [7:0] v_11224;
  wire [7:0] v_11225;
  function [7:0] mux_11225(input [0:0] sel);
    case (sel) 0: mux_11225 = 8'h0; 1: mux_11225 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11226;
  wire [7:0] v_11227;
  wire [7:0] v_11228;
  function [7:0] mux_11228(input [0:0] sel);
    case (sel) 0: mux_11228 = 8'h0; 1: mux_11228 = vout_peek_795;
    endcase
  endfunction
  wire [7:0] v_11229;
  function [7:0] mux_11229(input [0:0] sel);
    case (sel) 0: mux_11229 = 8'h0; 1: mux_11229 = vout_peek_787;
    endcase
  endfunction
  wire [7:0] v_11230;
  function [7:0] mux_11230(input [0:0] sel);
    case (sel) 0: mux_11230 = 8'h0; 1: mux_11230 = v_11231;
    endcase
  endfunction
  reg [7:0] v_11231 = 8'h0;
  wire [7:0] v_11232;
  wire [7:0] v_11233;
  function [7:0] mux_11233(input [0:0] sel);
    case (sel) 0: mux_11233 = 8'h0; 1: mux_11233 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11234;
  wire [7:0] v_11235;
  wire [7:0] v_11236;
  function [7:0] mux_11236(input [0:0] sel);
    case (sel) 0: mux_11236 = 8'h0; 1: mux_11236 = v_11237;
    endcase
  endfunction
  reg [7:0] v_11237 = 8'h0;
  wire [7:0] v_11238;
  wire [7:0] v_11239;
  function [7:0] mux_11239(input [0:0] sel);
    case (sel) 0: mux_11239 = 8'h0; 1: mux_11239 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11240;
  wire [7:0] v_11241;
  wire [7:0] v_11242;
  function [7:0] mux_11242(input [0:0] sel);
    case (sel) 0: mux_11242 = 8'h0; 1: mux_11242 = v_11243;
    endcase
  endfunction
  reg [7:0] v_11243 = 8'h0;
  wire [7:0] v_11244;
  wire [7:0] v_11245;
  function [7:0] mux_11245(input [0:0] sel);
    case (sel) 0: mux_11245 = 8'h0; 1: mux_11245 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11246;
  wire [7:0] v_11247;
  wire [7:0] v_11248;
  function [7:0] mux_11248(input [0:0] sel);
    case (sel) 0: mux_11248 = 8'h0; 1: mux_11248 = v_11249;
    endcase
  endfunction
  reg [7:0] v_11249 = 8'h0;
  wire [7:0] v_11250;
  wire [7:0] v_11251;
  function [7:0] mux_11251(input [0:0] sel);
    case (sel) 0: mux_11251 = 8'h0; 1: mux_11251 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11252;
  wire [7:0] v_11253;
  wire [7:0] v_11254;
  function [7:0] mux_11254(input [0:0] sel);
    case (sel) 0: mux_11254 = 8'h0; 1: mux_11254 = vout_peek_781;
    endcase
  endfunction
  wire [7:0] v_11255;
  function [7:0] mux_11255(input [0:0] sel);
    case (sel) 0: mux_11255 = 8'h0; 1: mux_11255 = vout_peek_773;
    endcase
  endfunction
  wire [7:0] v_11256;
  function [7:0] mux_11256(input [0:0] sel);
    case (sel) 0: mux_11256 = 8'h0; 1: mux_11256 = v_11257;
    endcase
  endfunction
  reg [7:0] v_11257 = 8'h0;
  wire [7:0] v_11258;
  wire [7:0] v_11259;
  function [7:0] mux_11259(input [0:0] sel);
    case (sel) 0: mux_11259 = 8'h0; 1: mux_11259 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11260;
  wire [7:0] v_11261;
  wire [7:0] v_11262;
  function [7:0] mux_11262(input [0:0] sel);
    case (sel) 0: mux_11262 = 8'h0; 1: mux_11262 = vout_peek_767;
    endcase
  endfunction
  wire [7:0] v_11263;
  function [7:0] mux_11263(input [0:0] sel);
    case (sel) 0: mux_11263 = 8'h0; 1: mux_11263 = vout_peek_759;
    endcase
  endfunction
  wire [7:0] v_11264;
  function [7:0] mux_11264(input [0:0] sel);
    case (sel) 0: mux_11264 = 8'h0; 1: mux_11264 = v_11265;
    endcase
  endfunction
  reg [7:0] v_11265 = 8'h0;
  wire [7:0] v_11266;
  wire [7:0] v_11267;
  function [7:0] mux_11267(input [0:0] sel);
    case (sel) 0: mux_11267 = 8'h0; 1: mux_11267 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11268;
  wire [7:0] v_11269;
  wire [7:0] v_11270;
  function [7:0] mux_11270(input [0:0] sel);
    case (sel) 0: mux_11270 = 8'h0; 1: mux_11270 = v_11271;
    endcase
  endfunction
  reg [7:0] v_11271 = 8'h0;
  wire [7:0] v_11272;
  wire [7:0] v_11273;
  function [7:0] mux_11273(input [0:0] sel);
    case (sel) 0: mux_11273 = 8'h0; 1: mux_11273 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11274;
  wire [7:0] v_11275;
  wire [7:0] v_11276;
  function [7:0] mux_11276(input [0:0] sel);
    case (sel) 0: mux_11276 = 8'h0; 1: mux_11276 = vout_peek_753;
    endcase
  endfunction
  wire [7:0] v_11277;
  function [7:0] mux_11277(input [0:0] sel);
    case (sel) 0: mux_11277 = 8'h0; 1: mux_11277 = vout_peek_745;
    endcase
  endfunction
  wire [7:0] v_11278;
  function [7:0] mux_11278(input [0:0] sel);
    case (sel) 0: mux_11278 = 8'h0; 1: mux_11278 = v_11279;
    endcase
  endfunction
  reg [7:0] v_11279 = 8'h0;
  wire [7:0] v_11280;
  wire [7:0] v_11281;
  function [7:0] mux_11281(input [0:0] sel);
    case (sel) 0: mux_11281 = 8'h0; 1: mux_11281 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11282;
  wire [7:0] v_11283;
  wire [7:0] v_11284;
  function [7:0] mux_11284(input [0:0] sel);
    case (sel) 0: mux_11284 = 8'h0; 1: mux_11284 = vout_peek_739;
    endcase
  endfunction
  wire [7:0] v_11285;
  function [7:0] mux_11285(input [0:0] sel);
    case (sel) 0: mux_11285 = 8'h0; 1: mux_11285 = vout_peek_731;
    endcase
  endfunction
  wire [7:0] v_11286;
  function [7:0] mux_11286(input [0:0] sel);
    case (sel) 0: mux_11286 = 8'h0; 1: mux_11286 = v_11287;
    endcase
  endfunction
  reg [7:0] v_11287 = 8'h0;
  wire [7:0] v_11288;
  wire [7:0] v_11289;
  function [7:0] mux_11289(input [0:0] sel);
    case (sel) 0: mux_11289 = 8'h0; 1: mux_11289 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11290;
  wire [7:0] v_11291;
  wire [7:0] v_11292;
  function [7:0] mux_11292(input [0:0] sel);
    case (sel) 0: mux_11292 = 8'h0; 1: mux_11292 = v_11293;
    endcase
  endfunction
  reg [7:0] v_11293 = 8'h0;
  wire [7:0] v_11294;
  wire [7:0] v_11295;
  function [7:0] mux_11295(input [0:0] sel);
    case (sel) 0: mux_11295 = 8'h0; 1: mux_11295 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11296;
  wire [7:0] v_11297;
  wire [7:0] v_11298;
  function [7:0] mux_11298(input [0:0] sel);
    case (sel) 0: mux_11298 = 8'h0; 1: mux_11298 = v_11299;
    endcase
  endfunction
  reg [7:0] v_11299 = 8'h0;
  wire [7:0] v_11300;
  wire [7:0] v_11301;
  function [7:0] mux_11301(input [0:0] sel);
    case (sel) 0: mux_11301 = 8'h0; 1: mux_11301 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11302;
  wire [7:0] v_11303;
  wire [7:0] v_11304;
  function [7:0] mux_11304(input [0:0] sel);
    case (sel) 0: mux_11304 = 8'h0; 1: mux_11304 = vout_peek_725;
    endcase
  endfunction
  wire [7:0] v_11305;
  function [7:0] mux_11305(input [0:0] sel);
    case (sel) 0: mux_11305 = 8'h0; 1: mux_11305 = vout_peek_717;
    endcase
  endfunction
  wire [7:0] v_11306;
  function [7:0] mux_11306(input [0:0] sel);
    case (sel) 0: mux_11306 = 8'h0; 1: mux_11306 = v_11307;
    endcase
  endfunction
  reg [7:0] v_11307 = 8'h0;
  wire [7:0] v_11308;
  wire [7:0] v_11309;
  function [7:0] mux_11309(input [0:0] sel);
    case (sel) 0: mux_11309 = 8'h0; 1: mux_11309 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11310;
  wire [7:0] v_11311;
  wire [7:0] v_11312;
  function [7:0] mux_11312(input [0:0] sel);
    case (sel) 0: mux_11312 = 8'h0; 1: mux_11312 = vout_peek_711;
    endcase
  endfunction
  wire [7:0] v_11313;
  function [7:0] mux_11313(input [0:0] sel);
    case (sel) 0: mux_11313 = 8'h0; 1: mux_11313 = vout_peek_703;
    endcase
  endfunction
  wire [7:0] v_11314;
  function [7:0] mux_11314(input [0:0] sel);
    case (sel) 0: mux_11314 = 8'h0; 1: mux_11314 = v_11315;
    endcase
  endfunction
  reg [7:0] v_11315 = 8'h0;
  wire [7:0] v_11316;
  wire [7:0] v_11317;
  function [7:0] mux_11317(input [0:0] sel);
    case (sel) 0: mux_11317 = 8'h0; 1: mux_11317 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11318;
  wire [7:0] v_11319;
  wire [7:0] v_11320;
  function [7:0] mux_11320(input [0:0] sel);
    case (sel) 0: mux_11320 = 8'h0; 1: mux_11320 = v_11321;
    endcase
  endfunction
  reg [7:0] v_11321 = 8'h0;
  wire [7:0] v_11322;
  wire [7:0] v_11323;
  function [7:0] mux_11323(input [0:0] sel);
    case (sel) 0: mux_11323 = 8'h0; 1: mux_11323 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11324;
  wire [7:0] v_11325;
  wire [7:0] v_11326;
  function [7:0] mux_11326(input [0:0] sel);
    case (sel) 0: mux_11326 = 8'h0; 1: mux_11326 = vout_peek_697;
    endcase
  endfunction
  wire [7:0] v_11327;
  function [7:0] mux_11327(input [0:0] sel);
    case (sel) 0: mux_11327 = 8'h0; 1: mux_11327 = vout_peek_689;
    endcase
  endfunction
  wire [7:0] v_11328;
  function [7:0] mux_11328(input [0:0] sel);
    case (sel) 0: mux_11328 = 8'h0; 1: mux_11328 = v_11329;
    endcase
  endfunction
  reg [7:0] v_11329 = 8'h0;
  wire [7:0] v_11330;
  wire [7:0] v_11331;
  function [7:0] mux_11331(input [0:0] sel);
    case (sel) 0: mux_11331 = 8'h0; 1: mux_11331 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11332;
  wire [7:0] v_11333;
  wire [7:0] v_11334;
  function [7:0] mux_11334(input [0:0] sel);
    case (sel) 0: mux_11334 = 8'h0; 1: mux_11334 = vout_peek_683;
    endcase
  endfunction
  wire [7:0] v_11335;
  function [7:0] mux_11335(input [0:0] sel);
    case (sel) 0: mux_11335 = 8'h0; 1: mux_11335 = vout_peek_675;
    endcase
  endfunction
  wire [7:0] v_11336;
  function [7:0] mux_11336(input [0:0] sel);
    case (sel) 0: mux_11336 = 8'h0; 1: mux_11336 = v_11337;
    endcase
  endfunction
  reg [7:0] v_11337 = 8'h0;
  wire [7:0] v_11338;
  wire [7:0] v_11339;
  function [7:0] mux_11339(input [0:0] sel);
    case (sel) 0: mux_11339 = 8'h0; 1: mux_11339 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11340;
  wire [7:0] v_11341;
  wire [7:0] v_11342;
  function [7:0] mux_11342(input [0:0] sel);
    case (sel) 0: mux_11342 = 8'h0; 1: mux_11342 = v_11343;
    endcase
  endfunction
  reg [7:0] v_11343 = 8'h0;
  wire [7:0] v_11344;
  wire [7:0] v_11345;
  function [7:0] mux_11345(input [0:0] sel);
    case (sel) 0: mux_11345 = 8'h0; 1: mux_11345 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11346;
  wire [7:0] v_11347;
  wire [7:0] v_11348;
  function [7:0] mux_11348(input [0:0] sel);
    case (sel) 0: mux_11348 = 8'h0; 1: mux_11348 = v_11349;
    endcase
  endfunction
  reg [7:0] v_11349 = 8'h0;
  wire [7:0] v_11350;
  wire [7:0] v_11351;
  function [7:0] mux_11351(input [0:0] sel);
    case (sel) 0: mux_11351 = 8'h0; 1: mux_11351 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11352;
  wire [7:0] v_11353;
  wire [7:0] v_11354;
  function [7:0] mux_11354(input [0:0] sel);
    case (sel) 0: mux_11354 = 8'h0; 1: mux_11354 = v_11355;
    endcase
  endfunction
  reg [7:0] v_11355 = 8'h0;
  wire [7:0] v_11356;
  wire [7:0] v_11357;
  function [7:0] mux_11357(input [0:0] sel);
    case (sel) 0: mux_11357 = 8'h0; 1: mux_11357 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11358;
  wire [7:0] v_11359;
  wire [7:0] v_11360;
  function [7:0] mux_11360(input [0:0] sel);
    case (sel) 0: mux_11360 = 8'h0; 1: mux_11360 = v_11361;
    endcase
  endfunction
  reg [7:0] v_11361 = 8'h0;
  wire [7:0] v_11362;
  wire [7:0] v_11363;
  function [7:0] mux_11363(input [0:0] sel);
    case (sel) 0: mux_11363 = 8'h0; 1: mux_11363 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11364;
  wire [7:0] v_11365;
  wire [7:0] v_11366;
  function [7:0] mux_11366(input [0:0] sel);
    case (sel) 0: mux_11366 = 8'h0; 1: mux_11366 = v_11367;
    endcase
  endfunction
  reg [7:0] v_11367 = 8'h0;
  wire [7:0] v_11368;
  wire [7:0] v_11369;
  function [7:0] mux_11369(input [0:0] sel);
    case (sel) 0: mux_11369 = 8'h0; 1: mux_11369 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11370;
  wire [7:0] v_11371;
  wire [7:0] v_11372;
  function [7:0] mux_11372(input [0:0] sel);
    case (sel) 0: mux_11372 = 8'h0; 1: mux_11372 = vout_peek_669;
    endcase
  endfunction
  wire [7:0] v_11373;
  function [7:0] mux_11373(input [0:0] sel);
    case (sel) 0: mux_11373 = 8'h0; 1: mux_11373 = vout_peek_661;
    endcase
  endfunction
  wire [7:0] v_11374;
  function [7:0] mux_11374(input [0:0] sel);
    case (sel) 0: mux_11374 = 8'h0; 1: mux_11374 = v_11375;
    endcase
  endfunction
  reg [7:0] v_11375 = 8'h0;
  wire [7:0] v_11376;
  wire [7:0] v_11377;
  function [7:0] mux_11377(input [0:0] sel);
    case (sel) 0: mux_11377 = 8'h0; 1: mux_11377 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11378;
  wire [7:0] v_11379;
  wire [7:0] v_11380;
  function [7:0] mux_11380(input [0:0] sel);
    case (sel) 0: mux_11380 = 8'h0; 1: mux_11380 = vout_peek_655;
    endcase
  endfunction
  wire [7:0] v_11381;
  function [7:0] mux_11381(input [0:0] sel);
    case (sel) 0: mux_11381 = 8'h0; 1: mux_11381 = vout_peek_647;
    endcase
  endfunction
  wire [7:0] v_11382;
  function [7:0] mux_11382(input [0:0] sel);
    case (sel) 0: mux_11382 = 8'h0; 1: mux_11382 = v_11383;
    endcase
  endfunction
  reg [7:0] v_11383 = 8'h0;
  wire [7:0] v_11384;
  wire [7:0] v_11385;
  function [7:0] mux_11385(input [0:0] sel);
    case (sel) 0: mux_11385 = 8'h0; 1: mux_11385 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11386;
  wire [7:0] v_11387;
  wire [7:0] v_11388;
  function [7:0] mux_11388(input [0:0] sel);
    case (sel) 0: mux_11388 = 8'h0; 1: mux_11388 = v_11389;
    endcase
  endfunction
  reg [7:0] v_11389 = 8'h0;
  wire [7:0] v_11390;
  wire [7:0] v_11391;
  function [7:0] mux_11391(input [0:0] sel);
    case (sel) 0: mux_11391 = 8'h0; 1: mux_11391 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11392;
  wire [7:0] v_11393;
  wire [7:0] v_11394;
  function [7:0] mux_11394(input [0:0] sel);
    case (sel) 0: mux_11394 = 8'h0; 1: mux_11394 = vout_peek_641;
    endcase
  endfunction
  wire [7:0] v_11395;
  function [7:0] mux_11395(input [0:0] sel);
    case (sel) 0: mux_11395 = 8'h0; 1: mux_11395 = vout_peek_633;
    endcase
  endfunction
  wire [7:0] v_11396;
  function [7:0] mux_11396(input [0:0] sel);
    case (sel) 0: mux_11396 = 8'h0; 1: mux_11396 = v_11397;
    endcase
  endfunction
  reg [7:0] v_11397 = 8'h0;
  wire [7:0] v_11398;
  wire [7:0] v_11399;
  function [7:0] mux_11399(input [0:0] sel);
    case (sel) 0: mux_11399 = 8'h0; 1: mux_11399 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11400;
  wire [7:0] v_11401;
  wire [7:0] v_11402;
  function [7:0] mux_11402(input [0:0] sel);
    case (sel) 0: mux_11402 = 8'h0; 1: mux_11402 = vout_peek_627;
    endcase
  endfunction
  wire [7:0] v_11403;
  function [7:0] mux_11403(input [0:0] sel);
    case (sel) 0: mux_11403 = 8'h0; 1: mux_11403 = vout_peek_619;
    endcase
  endfunction
  wire [7:0] v_11404;
  function [7:0] mux_11404(input [0:0] sel);
    case (sel) 0: mux_11404 = 8'h0; 1: mux_11404 = v_11405;
    endcase
  endfunction
  reg [7:0] v_11405 = 8'h0;
  wire [7:0] v_11406;
  wire [7:0] v_11407;
  function [7:0] mux_11407(input [0:0] sel);
    case (sel) 0: mux_11407 = 8'h0; 1: mux_11407 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11408;
  wire [7:0] v_11409;
  wire [7:0] v_11410;
  function [7:0] mux_11410(input [0:0] sel);
    case (sel) 0: mux_11410 = 8'h0; 1: mux_11410 = v_11411;
    endcase
  endfunction
  reg [7:0] v_11411 = 8'h0;
  wire [7:0] v_11412;
  wire [7:0] v_11413;
  function [7:0] mux_11413(input [0:0] sel);
    case (sel) 0: mux_11413 = 8'h0; 1: mux_11413 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11414;
  wire [7:0] v_11415;
  wire [7:0] v_11416;
  function [7:0] mux_11416(input [0:0] sel);
    case (sel) 0: mux_11416 = 8'h0; 1: mux_11416 = v_11417;
    endcase
  endfunction
  reg [7:0] v_11417 = 8'h0;
  wire [7:0] v_11418;
  wire [7:0] v_11419;
  function [7:0] mux_11419(input [0:0] sel);
    case (sel) 0: mux_11419 = 8'h0; 1: mux_11419 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11420;
  wire [7:0] v_11421;
  wire [7:0] v_11422;
  function [7:0] mux_11422(input [0:0] sel);
    case (sel) 0: mux_11422 = 8'h0; 1: mux_11422 = vout_peek_613;
    endcase
  endfunction
  wire [7:0] v_11423;
  function [7:0] mux_11423(input [0:0] sel);
    case (sel) 0: mux_11423 = 8'h0; 1: mux_11423 = vout_peek_605;
    endcase
  endfunction
  wire [7:0] v_11424;
  function [7:0] mux_11424(input [0:0] sel);
    case (sel) 0: mux_11424 = 8'h0; 1: mux_11424 = v_11425;
    endcase
  endfunction
  reg [7:0] v_11425 = 8'h0;
  wire [7:0] v_11426;
  wire [7:0] v_11427;
  function [7:0] mux_11427(input [0:0] sel);
    case (sel) 0: mux_11427 = 8'h0; 1: mux_11427 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11428;
  wire [7:0] v_11429;
  wire [7:0] v_11430;
  function [7:0] mux_11430(input [0:0] sel);
    case (sel) 0: mux_11430 = 8'h0; 1: mux_11430 = vout_peek_599;
    endcase
  endfunction
  wire [7:0] v_11431;
  function [7:0] mux_11431(input [0:0] sel);
    case (sel) 0: mux_11431 = 8'h0; 1: mux_11431 = vout_peek_591;
    endcase
  endfunction
  wire [7:0] v_11432;
  function [7:0] mux_11432(input [0:0] sel);
    case (sel) 0: mux_11432 = 8'h0; 1: mux_11432 = v_11433;
    endcase
  endfunction
  reg [7:0] v_11433 = 8'h0;
  wire [7:0] v_11434;
  wire [7:0] v_11435;
  function [7:0] mux_11435(input [0:0] sel);
    case (sel) 0: mux_11435 = 8'h0; 1: mux_11435 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11436;
  wire [7:0] v_11437;
  wire [7:0] v_11438;
  function [7:0] mux_11438(input [0:0] sel);
    case (sel) 0: mux_11438 = 8'h0; 1: mux_11438 = v_11439;
    endcase
  endfunction
  reg [7:0] v_11439 = 8'h0;
  wire [7:0] v_11440;
  wire [7:0] v_11441;
  function [7:0] mux_11441(input [0:0] sel);
    case (sel) 0: mux_11441 = 8'h0; 1: mux_11441 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11442;
  wire [7:0] v_11443;
  wire [7:0] v_11444;
  function [7:0] mux_11444(input [0:0] sel);
    case (sel) 0: mux_11444 = 8'h0; 1: mux_11444 = vout_peek_585;
    endcase
  endfunction
  wire [7:0] v_11445;
  function [7:0] mux_11445(input [0:0] sel);
    case (sel) 0: mux_11445 = 8'h0; 1: mux_11445 = vout_peek_577;
    endcase
  endfunction
  wire [7:0] v_11446;
  function [7:0] mux_11446(input [0:0] sel);
    case (sel) 0: mux_11446 = 8'h0; 1: mux_11446 = v_11447;
    endcase
  endfunction
  reg [7:0] v_11447 = 8'h0;
  wire [7:0] v_11448;
  wire [7:0] v_11449;
  function [7:0] mux_11449(input [0:0] sel);
    case (sel) 0: mux_11449 = 8'h0; 1: mux_11449 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11450;
  wire [7:0] v_11451;
  wire [7:0] v_11452;
  function [7:0] mux_11452(input [0:0] sel);
    case (sel) 0: mux_11452 = 8'h0; 1: mux_11452 = vout_peek_571;
    endcase
  endfunction
  wire [7:0] v_11453;
  function [7:0] mux_11453(input [0:0] sel);
    case (sel) 0: mux_11453 = 8'h0; 1: mux_11453 = vout_peek_563;
    endcase
  endfunction
  wire [7:0] v_11454;
  function [7:0] mux_11454(input [0:0] sel);
    case (sel) 0: mux_11454 = 8'h0; 1: mux_11454 = v_11455;
    endcase
  endfunction
  reg [7:0] v_11455 = 8'h0;
  wire [7:0] v_11456;
  wire [7:0] v_11457;
  function [7:0] mux_11457(input [0:0] sel);
    case (sel) 0: mux_11457 = 8'h0; 1: mux_11457 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11458;
  wire [7:0] v_11459;
  wire [7:0] v_11460;
  function [7:0] mux_11460(input [0:0] sel);
    case (sel) 0: mux_11460 = 8'h0; 1: mux_11460 = v_11461;
    endcase
  endfunction
  reg [7:0] v_11461 = 8'h0;
  wire [7:0] v_11462;
  wire [7:0] v_11463;
  function [7:0] mux_11463(input [0:0] sel);
    case (sel) 0: mux_11463 = 8'h0; 1: mux_11463 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11464;
  wire [7:0] v_11465;
  wire [7:0] v_11466;
  function [7:0] mux_11466(input [0:0] sel);
    case (sel) 0: mux_11466 = 8'h0; 1: mux_11466 = v_11467;
    endcase
  endfunction
  reg [7:0] v_11467 = 8'h0;
  wire [7:0] v_11468;
  wire [7:0] v_11469;
  function [7:0] mux_11469(input [0:0] sel);
    case (sel) 0: mux_11469 = 8'h0; 1: mux_11469 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11470;
  wire [7:0] v_11471;
  wire [7:0] v_11472;
  function [7:0] mux_11472(input [0:0] sel);
    case (sel) 0: mux_11472 = 8'h0; 1: mux_11472 = v_11473;
    endcase
  endfunction
  reg [7:0] v_11473 = 8'h0;
  wire [7:0] v_11474;
  wire [7:0] v_11475;
  function [7:0] mux_11475(input [0:0] sel);
    case (sel) 0: mux_11475 = 8'h0; 1: mux_11475 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11476;
  wire [7:0] v_11477;
  wire [7:0] v_11478;
  function [7:0] mux_11478(input [0:0] sel);
    case (sel) 0: mux_11478 = 8'h0; 1: mux_11478 = vout_peek_557;
    endcase
  endfunction
  wire [7:0] v_11479;
  function [7:0] mux_11479(input [0:0] sel);
    case (sel) 0: mux_11479 = 8'h0; 1: mux_11479 = vout_peek_549;
    endcase
  endfunction
  wire [7:0] v_11480;
  function [7:0] mux_11480(input [0:0] sel);
    case (sel) 0: mux_11480 = 8'h0; 1: mux_11480 = v_11481;
    endcase
  endfunction
  reg [7:0] v_11481 = 8'h0;
  wire [7:0] v_11482;
  wire [7:0] v_11483;
  function [7:0] mux_11483(input [0:0] sel);
    case (sel) 0: mux_11483 = 8'h0; 1: mux_11483 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11484;
  wire [7:0] v_11485;
  wire [7:0] v_11486;
  function [7:0] mux_11486(input [0:0] sel);
    case (sel) 0: mux_11486 = 8'h0; 1: mux_11486 = vout_peek_543;
    endcase
  endfunction
  wire [7:0] v_11487;
  function [7:0] mux_11487(input [0:0] sel);
    case (sel) 0: mux_11487 = 8'h0; 1: mux_11487 = vout_peek_535;
    endcase
  endfunction
  wire [7:0] v_11488;
  function [7:0] mux_11488(input [0:0] sel);
    case (sel) 0: mux_11488 = 8'h0; 1: mux_11488 = v_11489;
    endcase
  endfunction
  reg [7:0] v_11489 = 8'h0;
  wire [7:0] v_11490;
  wire [7:0] v_11491;
  function [7:0] mux_11491(input [0:0] sel);
    case (sel) 0: mux_11491 = 8'h0; 1: mux_11491 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11492;
  wire [7:0] v_11493;
  wire [7:0] v_11494;
  function [7:0] mux_11494(input [0:0] sel);
    case (sel) 0: mux_11494 = 8'h0; 1: mux_11494 = v_11495;
    endcase
  endfunction
  reg [7:0] v_11495 = 8'h0;
  wire [7:0] v_11496;
  wire [7:0] v_11497;
  function [7:0] mux_11497(input [0:0] sel);
    case (sel) 0: mux_11497 = 8'h0; 1: mux_11497 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11498;
  wire [7:0] v_11499;
  wire [7:0] v_11500;
  function [7:0] mux_11500(input [0:0] sel);
    case (sel) 0: mux_11500 = 8'h0; 1: mux_11500 = vout_peek_529;
    endcase
  endfunction
  wire [7:0] v_11501;
  function [7:0] mux_11501(input [0:0] sel);
    case (sel) 0: mux_11501 = 8'h0; 1: mux_11501 = vout_peek_521;
    endcase
  endfunction
  wire [7:0] v_11502;
  function [7:0] mux_11502(input [0:0] sel);
    case (sel) 0: mux_11502 = 8'h0; 1: mux_11502 = v_11503;
    endcase
  endfunction
  reg [7:0] v_11503 = 8'h0;
  wire [7:0] v_11504;
  wire [7:0] v_11505;
  function [7:0] mux_11505(input [0:0] sel);
    case (sel) 0: mux_11505 = 8'h0; 1: mux_11505 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11506;
  wire [7:0] v_11507;
  wire [7:0] v_11508;
  function [7:0] mux_11508(input [0:0] sel);
    case (sel) 0: mux_11508 = 8'h0; 1: mux_11508 = vout_peek_515;
    endcase
  endfunction
  wire [7:0] v_11509;
  function [7:0] mux_11509(input [0:0] sel);
    case (sel) 0: mux_11509 = 8'h0; 1: mux_11509 = vout_peek_507;
    endcase
  endfunction
  wire [7:0] v_11510;
  function [7:0] mux_11510(input [0:0] sel);
    case (sel) 0: mux_11510 = 8'h0; 1: mux_11510 = v_11511;
    endcase
  endfunction
  reg [7:0] v_11511 = 8'h0;
  wire [7:0] v_11512;
  wire [7:0] v_11513;
  function [7:0] mux_11513(input [0:0] sel);
    case (sel) 0: mux_11513 = 8'h0; 1: mux_11513 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11514;
  wire [7:0] v_11515;
  wire [7:0] v_11516;
  function [7:0] mux_11516(input [0:0] sel);
    case (sel) 0: mux_11516 = 8'h0; 1: mux_11516 = v_11517;
    endcase
  endfunction
  reg [7:0] v_11517 = 8'h0;
  wire [7:0] v_11518;
  wire [7:0] v_11519;
  function [7:0] mux_11519(input [0:0] sel);
    case (sel) 0: mux_11519 = 8'h0; 1: mux_11519 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11520;
  wire [7:0] v_11521;
  wire [7:0] v_11522;
  function [7:0] mux_11522(input [0:0] sel);
    case (sel) 0: mux_11522 = 8'h0; 1: mux_11522 = v_11523;
    endcase
  endfunction
  reg [7:0] v_11523 = 8'h0;
  wire [7:0] v_11524;
  wire [7:0] v_11525;
  function [7:0] mux_11525(input [0:0] sel);
    case (sel) 0: mux_11525 = 8'h0; 1: mux_11525 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11526;
  wire [7:0] v_11527;
  wire [7:0] v_11528;
  function [7:0] mux_11528(input [0:0] sel);
    case (sel) 0: mux_11528 = 8'h0; 1: mux_11528 = vout_peek_501;
    endcase
  endfunction
  wire [7:0] v_11529;
  function [7:0] mux_11529(input [0:0] sel);
    case (sel) 0: mux_11529 = 8'h0; 1: mux_11529 = vout_peek_493;
    endcase
  endfunction
  wire [7:0] v_11530;
  function [7:0] mux_11530(input [0:0] sel);
    case (sel) 0: mux_11530 = 8'h0; 1: mux_11530 = v_11531;
    endcase
  endfunction
  reg [7:0] v_11531 = 8'h0;
  wire [7:0] v_11532;
  wire [7:0] v_11533;
  function [7:0] mux_11533(input [0:0] sel);
    case (sel) 0: mux_11533 = 8'h0; 1: mux_11533 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11534;
  wire [7:0] v_11535;
  wire [7:0] v_11536;
  function [7:0] mux_11536(input [0:0] sel);
    case (sel) 0: mux_11536 = 8'h0; 1: mux_11536 = vout_peek_487;
    endcase
  endfunction
  wire [7:0] v_11537;
  function [7:0] mux_11537(input [0:0] sel);
    case (sel) 0: mux_11537 = 8'h0; 1: mux_11537 = vout_peek_479;
    endcase
  endfunction
  wire [7:0] v_11538;
  function [7:0] mux_11538(input [0:0] sel);
    case (sel) 0: mux_11538 = 8'h0; 1: mux_11538 = v_11539;
    endcase
  endfunction
  reg [7:0] v_11539 = 8'h0;
  wire [7:0] v_11540;
  wire [7:0] v_11541;
  function [7:0] mux_11541(input [0:0] sel);
    case (sel) 0: mux_11541 = 8'h0; 1: mux_11541 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11542;
  wire [7:0] v_11543;
  wire [7:0] v_11544;
  function [7:0] mux_11544(input [0:0] sel);
    case (sel) 0: mux_11544 = 8'h0; 1: mux_11544 = v_11545;
    endcase
  endfunction
  reg [7:0] v_11545 = 8'h0;
  wire [7:0] v_11546;
  wire [7:0] v_11547;
  function [7:0] mux_11547(input [0:0] sel);
    case (sel) 0: mux_11547 = 8'h0; 1: mux_11547 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11548;
  wire [7:0] v_11549;
  wire [7:0] v_11550;
  function [7:0] mux_11550(input [0:0] sel);
    case (sel) 0: mux_11550 = 8'h0; 1: mux_11550 = vout_peek_473;
    endcase
  endfunction
  wire [7:0] v_11551;
  function [7:0] mux_11551(input [0:0] sel);
    case (sel) 0: mux_11551 = 8'h0; 1: mux_11551 = vout_peek_465;
    endcase
  endfunction
  wire [7:0] v_11552;
  function [7:0] mux_11552(input [0:0] sel);
    case (sel) 0: mux_11552 = 8'h0; 1: mux_11552 = v_11553;
    endcase
  endfunction
  reg [7:0] v_11553 = 8'h0;
  wire [7:0] v_11554;
  wire [7:0] v_11555;
  function [7:0] mux_11555(input [0:0] sel);
    case (sel) 0: mux_11555 = 8'h0; 1: mux_11555 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11556;
  wire [7:0] v_11557;
  wire [7:0] v_11558;
  function [7:0] mux_11558(input [0:0] sel);
    case (sel) 0: mux_11558 = 8'h0; 1: mux_11558 = vout_peek_459;
    endcase
  endfunction
  wire [7:0] v_11559;
  function [7:0] mux_11559(input [0:0] sel);
    case (sel) 0: mux_11559 = 8'h0; 1: mux_11559 = vout_peek_451;
    endcase
  endfunction
  wire [7:0] v_11560;
  function [7:0] mux_11560(input [0:0] sel);
    case (sel) 0: mux_11560 = 8'h0; 1: mux_11560 = v_11561;
    endcase
  endfunction
  reg [7:0] v_11561 = 8'h0;
  wire [7:0] v_11562;
  wire [7:0] v_11563;
  function [7:0] mux_11563(input [0:0] sel);
    case (sel) 0: mux_11563 = 8'h0; 1: mux_11563 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11564;
  wire [7:0] v_11565;
  wire [7:0] v_11566;
  function [7:0] mux_11566(input [0:0] sel);
    case (sel) 0: mux_11566 = 8'h0; 1: mux_11566 = v_11567;
    endcase
  endfunction
  reg [7:0] v_11567 = 8'h0;
  wire [7:0] v_11568;
  wire [7:0] v_11569;
  function [7:0] mux_11569(input [0:0] sel);
    case (sel) 0: mux_11569 = 8'h0; 1: mux_11569 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11570;
  wire [7:0] v_11571;
  wire [7:0] v_11572;
  function [7:0] mux_11572(input [0:0] sel);
    case (sel) 0: mux_11572 = 8'h0; 1: mux_11572 = v_11573;
    endcase
  endfunction
  reg [7:0] v_11573 = 8'h0;
  wire [7:0] v_11574;
  wire [7:0] v_11575;
  function [7:0] mux_11575(input [0:0] sel);
    case (sel) 0: mux_11575 = 8'h0; 1: mux_11575 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11576;
  wire [7:0] v_11577;
  wire [7:0] v_11578;
  function [7:0] mux_11578(input [0:0] sel);
    case (sel) 0: mux_11578 = 8'h0; 1: mux_11578 = v_11579;
    endcase
  endfunction
  reg [7:0] v_11579 = 8'h0;
  wire [7:0] v_11580;
  wire [7:0] v_11581;
  function [7:0] mux_11581(input [0:0] sel);
    case (sel) 0: mux_11581 = 8'h0; 1: mux_11581 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11582;
  wire [7:0] v_11583;
  wire [7:0] v_11584;
  function [7:0] mux_11584(input [0:0] sel);
    case (sel) 0: mux_11584 = 8'h0; 1: mux_11584 = v_11585;
    endcase
  endfunction
  reg [7:0] v_11585 = 8'h0;
  wire [7:0] v_11586;
  wire [7:0] v_11587;
  function [7:0] mux_11587(input [0:0] sel);
    case (sel) 0: mux_11587 = 8'h0; 1: mux_11587 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11588;
  wire [7:0] v_11589;
  wire [7:0] v_11590;
  function [7:0] mux_11590(input [0:0] sel);
    case (sel) 0: mux_11590 = 8'h0; 1: mux_11590 = vout_peek_445;
    endcase
  endfunction
  wire [7:0] v_11591;
  function [7:0] mux_11591(input [0:0] sel);
    case (sel) 0: mux_11591 = 8'h0; 1: mux_11591 = vout_peek_437;
    endcase
  endfunction
  wire [7:0] v_11592;
  function [7:0] mux_11592(input [0:0] sel);
    case (sel) 0: mux_11592 = 8'h0; 1: mux_11592 = v_11593;
    endcase
  endfunction
  reg [7:0] v_11593 = 8'h0;
  wire [7:0] v_11594;
  wire [7:0] v_11595;
  function [7:0] mux_11595(input [0:0] sel);
    case (sel) 0: mux_11595 = 8'h0; 1: mux_11595 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11596;
  wire [7:0] v_11597;
  wire [7:0] v_11598;
  function [7:0] mux_11598(input [0:0] sel);
    case (sel) 0: mux_11598 = 8'h0; 1: mux_11598 = vout_peek_431;
    endcase
  endfunction
  wire [7:0] v_11599;
  function [7:0] mux_11599(input [0:0] sel);
    case (sel) 0: mux_11599 = 8'h0; 1: mux_11599 = vout_peek_423;
    endcase
  endfunction
  wire [7:0] v_11600;
  function [7:0] mux_11600(input [0:0] sel);
    case (sel) 0: mux_11600 = 8'h0; 1: mux_11600 = v_11601;
    endcase
  endfunction
  reg [7:0] v_11601 = 8'h0;
  wire [7:0] v_11602;
  wire [7:0] v_11603;
  function [7:0] mux_11603(input [0:0] sel);
    case (sel) 0: mux_11603 = 8'h0; 1: mux_11603 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11604;
  wire [7:0] v_11605;
  wire [7:0] v_11606;
  function [7:0] mux_11606(input [0:0] sel);
    case (sel) 0: mux_11606 = 8'h0; 1: mux_11606 = v_11607;
    endcase
  endfunction
  reg [7:0] v_11607 = 8'h0;
  wire [7:0] v_11608;
  wire [7:0] v_11609;
  function [7:0] mux_11609(input [0:0] sel);
    case (sel) 0: mux_11609 = 8'h0; 1: mux_11609 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11610;
  wire [7:0] v_11611;
  wire [7:0] v_11612;
  function [7:0] mux_11612(input [0:0] sel);
    case (sel) 0: mux_11612 = 8'h0; 1: mux_11612 = vout_peek_417;
    endcase
  endfunction
  wire [7:0] v_11613;
  function [7:0] mux_11613(input [0:0] sel);
    case (sel) 0: mux_11613 = 8'h0; 1: mux_11613 = vout_peek_409;
    endcase
  endfunction
  wire [7:0] v_11614;
  function [7:0] mux_11614(input [0:0] sel);
    case (sel) 0: mux_11614 = 8'h0; 1: mux_11614 = v_11615;
    endcase
  endfunction
  reg [7:0] v_11615 = 8'h0;
  wire [7:0] v_11616;
  wire [7:0] v_11617;
  function [7:0] mux_11617(input [0:0] sel);
    case (sel) 0: mux_11617 = 8'h0; 1: mux_11617 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11618;
  wire [7:0] v_11619;
  wire [7:0] v_11620;
  function [7:0] mux_11620(input [0:0] sel);
    case (sel) 0: mux_11620 = 8'h0; 1: mux_11620 = vout_peek_403;
    endcase
  endfunction
  wire [7:0] v_11621;
  function [7:0] mux_11621(input [0:0] sel);
    case (sel) 0: mux_11621 = 8'h0; 1: mux_11621 = vout_peek_395;
    endcase
  endfunction
  wire [7:0] v_11622;
  function [7:0] mux_11622(input [0:0] sel);
    case (sel) 0: mux_11622 = 8'h0; 1: mux_11622 = v_11623;
    endcase
  endfunction
  reg [7:0] v_11623 = 8'h0;
  wire [7:0] v_11624;
  wire [7:0] v_11625;
  function [7:0] mux_11625(input [0:0] sel);
    case (sel) 0: mux_11625 = 8'h0; 1: mux_11625 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11626;
  wire [7:0] v_11627;
  wire [7:0] v_11628;
  function [7:0] mux_11628(input [0:0] sel);
    case (sel) 0: mux_11628 = 8'h0; 1: mux_11628 = v_11629;
    endcase
  endfunction
  reg [7:0] v_11629 = 8'h0;
  wire [7:0] v_11630;
  wire [7:0] v_11631;
  function [7:0] mux_11631(input [0:0] sel);
    case (sel) 0: mux_11631 = 8'h0; 1: mux_11631 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11632;
  wire [7:0] v_11633;
  wire [7:0] v_11634;
  function [7:0] mux_11634(input [0:0] sel);
    case (sel) 0: mux_11634 = 8'h0; 1: mux_11634 = v_11635;
    endcase
  endfunction
  reg [7:0] v_11635 = 8'h0;
  wire [7:0] v_11636;
  wire [7:0] v_11637;
  function [7:0] mux_11637(input [0:0] sel);
    case (sel) 0: mux_11637 = 8'h0; 1: mux_11637 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11638;
  wire [7:0] v_11639;
  wire [7:0] v_11640;
  function [7:0] mux_11640(input [0:0] sel);
    case (sel) 0: mux_11640 = 8'h0; 1: mux_11640 = vout_peek_389;
    endcase
  endfunction
  wire [7:0] v_11641;
  function [7:0] mux_11641(input [0:0] sel);
    case (sel) 0: mux_11641 = 8'h0; 1: mux_11641 = vout_peek_381;
    endcase
  endfunction
  wire [7:0] v_11642;
  function [7:0] mux_11642(input [0:0] sel);
    case (sel) 0: mux_11642 = 8'h0; 1: mux_11642 = v_11643;
    endcase
  endfunction
  reg [7:0] v_11643 = 8'h0;
  wire [7:0] v_11644;
  wire [7:0] v_11645;
  function [7:0] mux_11645(input [0:0] sel);
    case (sel) 0: mux_11645 = 8'h0; 1: mux_11645 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11646;
  wire [7:0] v_11647;
  wire [7:0] v_11648;
  function [7:0] mux_11648(input [0:0] sel);
    case (sel) 0: mux_11648 = 8'h0; 1: mux_11648 = vout_peek_375;
    endcase
  endfunction
  wire [7:0] v_11649;
  function [7:0] mux_11649(input [0:0] sel);
    case (sel) 0: mux_11649 = 8'h0; 1: mux_11649 = vout_peek_367;
    endcase
  endfunction
  wire [7:0] v_11650;
  function [7:0] mux_11650(input [0:0] sel);
    case (sel) 0: mux_11650 = 8'h0; 1: mux_11650 = v_11651;
    endcase
  endfunction
  reg [7:0] v_11651 = 8'h0;
  wire [7:0] v_11652;
  wire [7:0] v_11653;
  function [7:0] mux_11653(input [0:0] sel);
    case (sel) 0: mux_11653 = 8'h0; 1: mux_11653 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11654;
  wire [7:0] v_11655;
  wire [7:0] v_11656;
  function [7:0] mux_11656(input [0:0] sel);
    case (sel) 0: mux_11656 = 8'h0; 1: mux_11656 = v_11657;
    endcase
  endfunction
  reg [7:0] v_11657 = 8'h0;
  wire [7:0] v_11658;
  wire [7:0] v_11659;
  function [7:0] mux_11659(input [0:0] sel);
    case (sel) 0: mux_11659 = 8'h0; 1: mux_11659 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11660;
  wire [7:0] v_11661;
  wire [7:0] v_11662;
  function [7:0] mux_11662(input [0:0] sel);
    case (sel) 0: mux_11662 = 8'h0; 1: mux_11662 = vout_peek_361;
    endcase
  endfunction
  wire [7:0] v_11663;
  function [7:0] mux_11663(input [0:0] sel);
    case (sel) 0: mux_11663 = 8'h0; 1: mux_11663 = vout_peek_353;
    endcase
  endfunction
  wire [7:0] v_11664;
  function [7:0] mux_11664(input [0:0] sel);
    case (sel) 0: mux_11664 = 8'h0; 1: mux_11664 = v_11665;
    endcase
  endfunction
  reg [7:0] v_11665 = 8'h0;
  wire [7:0] v_11666;
  wire [7:0] v_11667;
  function [7:0] mux_11667(input [0:0] sel);
    case (sel) 0: mux_11667 = 8'h0; 1: mux_11667 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11668;
  wire [7:0] v_11669;
  wire [7:0] v_11670;
  function [7:0] mux_11670(input [0:0] sel);
    case (sel) 0: mux_11670 = 8'h0; 1: mux_11670 = vout_peek_347;
    endcase
  endfunction
  wire [7:0] v_11671;
  function [7:0] mux_11671(input [0:0] sel);
    case (sel) 0: mux_11671 = 8'h0; 1: mux_11671 = vout_peek_339;
    endcase
  endfunction
  wire [7:0] v_11672;
  function [7:0] mux_11672(input [0:0] sel);
    case (sel) 0: mux_11672 = 8'h0; 1: mux_11672 = v_11673;
    endcase
  endfunction
  reg [7:0] v_11673 = 8'h0;
  wire [7:0] v_11674;
  wire [7:0] v_11675;
  function [7:0] mux_11675(input [0:0] sel);
    case (sel) 0: mux_11675 = 8'h0; 1: mux_11675 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11676;
  wire [7:0] v_11677;
  wire [7:0] v_11678;
  function [7:0] mux_11678(input [0:0] sel);
    case (sel) 0: mux_11678 = 8'h0; 1: mux_11678 = v_11679;
    endcase
  endfunction
  reg [7:0] v_11679 = 8'h0;
  wire [7:0] v_11680;
  wire [7:0] v_11681;
  function [7:0] mux_11681(input [0:0] sel);
    case (sel) 0: mux_11681 = 8'h0; 1: mux_11681 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11682;
  wire [7:0] v_11683;
  wire [7:0] v_11684;
  function [7:0] mux_11684(input [0:0] sel);
    case (sel) 0: mux_11684 = 8'h0; 1: mux_11684 = v_11685;
    endcase
  endfunction
  reg [7:0] v_11685 = 8'h0;
  wire [7:0] v_11686;
  wire [7:0] v_11687;
  function [7:0] mux_11687(input [0:0] sel);
    case (sel) 0: mux_11687 = 8'h0; 1: mux_11687 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11688;
  wire [7:0] v_11689;
  wire [7:0] v_11690;
  function [7:0] mux_11690(input [0:0] sel);
    case (sel) 0: mux_11690 = 8'h0; 1: mux_11690 = v_11691;
    endcase
  endfunction
  reg [7:0] v_11691 = 8'h0;
  wire [7:0] v_11692;
  wire [7:0] v_11693;
  function [7:0] mux_11693(input [0:0] sel);
    case (sel) 0: mux_11693 = 8'h0; 1: mux_11693 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11694;
  wire [7:0] v_11695;
  wire [7:0] v_11696;
  function [7:0] mux_11696(input [0:0] sel);
    case (sel) 0: mux_11696 = 8'h0; 1: mux_11696 = vout_peek_333;
    endcase
  endfunction
  wire [7:0] v_11697;
  function [7:0] mux_11697(input [0:0] sel);
    case (sel) 0: mux_11697 = 8'h0; 1: mux_11697 = vout_peek_325;
    endcase
  endfunction
  wire [7:0] v_11698;
  function [7:0] mux_11698(input [0:0] sel);
    case (sel) 0: mux_11698 = 8'h0; 1: mux_11698 = v_11699;
    endcase
  endfunction
  reg [7:0] v_11699 = 8'h0;
  wire [7:0] v_11700;
  wire [7:0] v_11701;
  function [7:0] mux_11701(input [0:0] sel);
    case (sel) 0: mux_11701 = 8'h0; 1: mux_11701 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11702;
  wire [7:0] v_11703;
  wire [7:0] v_11704;
  function [7:0] mux_11704(input [0:0] sel);
    case (sel) 0: mux_11704 = 8'h0; 1: mux_11704 = vout_peek_319;
    endcase
  endfunction
  wire [7:0] v_11705;
  function [7:0] mux_11705(input [0:0] sel);
    case (sel) 0: mux_11705 = 8'h0; 1: mux_11705 = vout_peek_311;
    endcase
  endfunction
  wire [7:0] v_11706;
  function [7:0] mux_11706(input [0:0] sel);
    case (sel) 0: mux_11706 = 8'h0; 1: mux_11706 = v_11707;
    endcase
  endfunction
  reg [7:0] v_11707 = 8'h0;
  wire [7:0] v_11708;
  wire [7:0] v_11709;
  function [7:0] mux_11709(input [0:0] sel);
    case (sel) 0: mux_11709 = 8'h0; 1: mux_11709 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11710;
  wire [7:0] v_11711;
  wire [7:0] v_11712;
  function [7:0] mux_11712(input [0:0] sel);
    case (sel) 0: mux_11712 = 8'h0; 1: mux_11712 = v_11713;
    endcase
  endfunction
  reg [7:0] v_11713 = 8'h0;
  wire [7:0] v_11714;
  wire [7:0] v_11715;
  function [7:0] mux_11715(input [0:0] sel);
    case (sel) 0: mux_11715 = 8'h0; 1: mux_11715 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11716;
  wire [7:0] v_11717;
  wire [7:0] v_11718;
  function [7:0] mux_11718(input [0:0] sel);
    case (sel) 0: mux_11718 = 8'h0; 1: mux_11718 = vout_peek_305;
    endcase
  endfunction
  wire [7:0] v_11719;
  function [7:0] mux_11719(input [0:0] sel);
    case (sel) 0: mux_11719 = 8'h0; 1: mux_11719 = vout_peek_297;
    endcase
  endfunction
  wire [7:0] v_11720;
  function [7:0] mux_11720(input [0:0] sel);
    case (sel) 0: mux_11720 = 8'h0; 1: mux_11720 = v_11721;
    endcase
  endfunction
  reg [7:0] v_11721 = 8'h0;
  wire [7:0] v_11722;
  wire [7:0] v_11723;
  function [7:0] mux_11723(input [0:0] sel);
    case (sel) 0: mux_11723 = 8'h0; 1: mux_11723 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11724;
  wire [7:0] v_11725;
  wire [7:0] v_11726;
  function [7:0] mux_11726(input [0:0] sel);
    case (sel) 0: mux_11726 = 8'h0; 1: mux_11726 = vout_peek_291;
    endcase
  endfunction
  wire [7:0] v_11727;
  function [7:0] mux_11727(input [0:0] sel);
    case (sel) 0: mux_11727 = 8'h0; 1: mux_11727 = vout_peek_283;
    endcase
  endfunction
  wire [7:0] v_11728;
  function [7:0] mux_11728(input [0:0] sel);
    case (sel) 0: mux_11728 = 8'h0; 1: mux_11728 = v_11729;
    endcase
  endfunction
  reg [7:0] v_11729 = 8'h0;
  wire [7:0] v_11730;
  wire [7:0] v_11731;
  function [7:0] mux_11731(input [0:0] sel);
    case (sel) 0: mux_11731 = 8'h0; 1: mux_11731 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11732;
  wire [7:0] v_11733;
  wire [7:0] v_11734;
  function [7:0] mux_11734(input [0:0] sel);
    case (sel) 0: mux_11734 = 8'h0; 1: mux_11734 = v_11735;
    endcase
  endfunction
  reg [7:0] v_11735 = 8'h0;
  wire [7:0] v_11736;
  wire [7:0] v_11737;
  function [7:0] mux_11737(input [0:0] sel);
    case (sel) 0: mux_11737 = 8'h0; 1: mux_11737 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11738;
  wire [7:0] v_11739;
  wire [7:0] v_11740;
  function [7:0] mux_11740(input [0:0] sel);
    case (sel) 0: mux_11740 = 8'h0; 1: mux_11740 = v_11741;
    endcase
  endfunction
  reg [7:0] v_11741 = 8'h0;
  wire [7:0] v_11742;
  wire [7:0] v_11743;
  function [7:0] mux_11743(input [0:0] sel);
    case (sel) 0: mux_11743 = 8'h0; 1: mux_11743 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11744;
  wire [7:0] v_11745;
  wire [7:0] v_11746;
  function [7:0] mux_11746(input [0:0] sel);
    case (sel) 0: mux_11746 = 8'h0; 1: mux_11746 = vout_peek_277;
    endcase
  endfunction
  wire [7:0] v_11747;
  function [7:0] mux_11747(input [0:0] sel);
    case (sel) 0: mux_11747 = 8'h0; 1: mux_11747 = vout_peek_269;
    endcase
  endfunction
  wire [7:0] v_11748;
  function [7:0] mux_11748(input [0:0] sel);
    case (sel) 0: mux_11748 = 8'h0; 1: mux_11748 = v_11749;
    endcase
  endfunction
  reg [7:0] v_11749 = 8'h0;
  wire [7:0] v_11750;
  wire [7:0] v_11751;
  function [7:0] mux_11751(input [0:0] sel);
    case (sel) 0: mux_11751 = 8'h0; 1: mux_11751 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11752;
  wire [7:0] v_11753;
  wire [7:0] v_11754;
  function [7:0] mux_11754(input [0:0] sel);
    case (sel) 0: mux_11754 = 8'h0; 1: mux_11754 = vout_peek_263;
    endcase
  endfunction
  wire [7:0] v_11755;
  function [7:0] mux_11755(input [0:0] sel);
    case (sel) 0: mux_11755 = 8'h0; 1: mux_11755 = vout_peek_255;
    endcase
  endfunction
  wire [7:0] v_11756;
  function [7:0] mux_11756(input [0:0] sel);
    case (sel) 0: mux_11756 = 8'h0; 1: mux_11756 = v_11757;
    endcase
  endfunction
  reg [7:0] v_11757 = 8'h0;
  wire [7:0] v_11758;
  wire [7:0] v_11759;
  function [7:0] mux_11759(input [0:0] sel);
    case (sel) 0: mux_11759 = 8'h0; 1: mux_11759 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11760;
  wire [7:0] v_11761;
  wire [7:0] v_11762;
  function [7:0] mux_11762(input [0:0] sel);
    case (sel) 0: mux_11762 = 8'h0; 1: mux_11762 = v_11763;
    endcase
  endfunction
  reg [7:0] v_11763 = 8'h0;
  wire [7:0] v_11764;
  wire [7:0] v_11765;
  function [7:0] mux_11765(input [0:0] sel);
    case (sel) 0: mux_11765 = 8'h0; 1: mux_11765 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11766;
  wire [7:0] v_11767;
  wire [7:0] v_11768;
  function [7:0] mux_11768(input [0:0] sel);
    case (sel) 0: mux_11768 = 8'h0; 1: mux_11768 = vout_peek_249;
    endcase
  endfunction
  wire [7:0] v_11769;
  function [7:0] mux_11769(input [0:0] sel);
    case (sel) 0: mux_11769 = 8'h0; 1: mux_11769 = vout_peek_241;
    endcase
  endfunction
  wire [7:0] v_11770;
  function [7:0] mux_11770(input [0:0] sel);
    case (sel) 0: mux_11770 = 8'h0; 1: mux_11770 = v_11771;
    endcase
  endfunction
  reg [7:0] v_11771 = 8'h0;
  wire [7:0] v_11772;
  wire [7:0] v_11773;
  function [7:0] mux_11773(input [0:0] sel);
    case (sel) 0: mux_11773 = 8'h0; 1: mux_11773 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11774;
  wire [7:0] v_11775;
  wire [7:0] v_11776;
  function [7:0] mux_11776(input [0:0] sel);
    case (sel) 0: mux_11776 = 8'h0; 1: mux_11776 = vout_peek_235;
    endcase
  endfunction
  wire [7:0] v_11777;
  function [7:0] mux_11777(input [0:0] sel);
    case (sel) 0: mux_11777 = 8'h0; 1: mux_11777 = vout_peek_227;
    endcase
  endfunction
  wire [7:0] v_11778;
  function [7:0] mux_11778(input [0:0] sel);
    case (sel) 0: mux_11778 = 8'h0; 1: mux_11778 = v_11779;
    endcase
  endfunction
  reg [7:0] v_11779 = 8'h0;
  wire [7:0] v_11780;
  wire [7:0] v_11781;
  function [7:0] mux_11781(input [0:0] sel);
    case (sel) 0: mux_11781 = 8'h0; 1: mux_11781 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11782;
  wire [7:0] v_11783;
  wire [7:0] v_11784;
  function [7:0] mux_11784(input [0:0] sel);
    case (sel) 0: mux_11784 = 8'h0; 1: mux_11784 = v_11785;
    endcase
  endfunction
  reg [7:0] v_11785 = 8'h0;
  wire [7:0] v_11786;
  wire [7:0] v_11787;
  function [7:0] mux_11787(input [0:0] sel);
    case (sel) 0: mux_11787 = 8'h0; 1: mux_11787 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11788;
  wire [7:0] v_11789;
  wire [7:0] v_11790;
  function [7:0] mux_11790(input [0:0] sel);
    case (sel) 0: mux_11790 = 8'h0; 1: mux_11790 = v_11791;
    endcase
  endfunction
  reg [7:0] v_11791 = 8'h0;
  wire [7:0] v_11792;
  wire [7:0] v_11793;
  function [7:0] mux_11793(input [0:0] sel);
    case (sel) 0: mux_11793 = 8'h0; 1: mux_11793 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11794;
  wire [7:0] v_11795;
  wire [7:0] v_11796;
  function [7:0] mux_11796(input [0:0] sel);
    case (sel) 0: mux_11796 = 8'h0; 1: mux_11796 = v_11797;
    endcase
  endfunction
  reg [7:0] v_11797 = 8'h0;
  wire [7:0] v_11798;
  wire [7:0] v_11799;
  function [7:0] mux_11799(input [0:0] sel);
    case (sel) 0: mux_11799 = 8'h0; 1: mux_11799 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11800;
  wire [7:0] v_11801;
  wire [7:0] v_11802;
  function [7:0] mux_11802(input [0:0] sel);
    case (sel) 0: mux_11802 = 8'h0; 1: mux_11802 = v_11803;
    endcase
  endfunction
  reg [7:0] v_11803 = 8'h0;
  wire [7:0] v_11804;
  wire [7:0] v_11805;
  function [7:0] mux_11805(input [0:0] sel);
    case (sel) 0: mux_11805 = 8'h0; 1: mux_11805 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11806;
  wire [7:0] v_11807;
  wire [7:0] v_11808;
  function [7:0] mux_11808(input [0:0] sel);
    case (sel) 0: mux_11808 = 8'h0; 1: mux_11808 = v_11809;
    endcase
  endfunction
  reg [7:0] v_11809 = 8'h0;
  wire [7:0] v_11810;
  wire [7:0] v_11811;
  function [7:0] mux_11811(input [0:0] sel);
    case (sel) 0: mux_11811 = 8'h0; 1: mux_11811 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11812;
  wire [7:0] v_11813;
  wire [7:0] v_11814;
  function [7:0] mux_11814(input [0:0] sel);
    case (sel) 0: mux_11814 = 8'h0; 1: mux_11814 = v_11815;
    endcase
  endfunction
  reg [7:0] v_11815 = 8'h0;
  wire [7:0] v_11816;
  wire [7:0] v_11817;
  function [7:0] mux_11817(input [0:0] sel);
    case (sel) 0: mux_11817 = 8'h0; 1: mux_11817 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11818;
  wire [7:0] v_11819;
  wire [7:0] v_11820;
  function [7:0] mux_11820(input [0:0] sel);
    case (sel) 0: mux_11820 = 8'h0; 1: mux_11820 = v_11821;
    endcase
  endfunction
  reg [7:0] v_11821 = 8'h0;
  wire [7:0] v_11822;
  wire [7:0] v_11823;
  function [7:0] mux_11823(input [0:0] sel);
    case (sel) 0: mux_11823 = 8'h0; 1: mux_11823 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11824;
  wire [7:0] v_11825;
  wire [7:0] v_11826;
  function [7:0] mux_11826(input [0:0] sel);
    case (sel) 0: mux_11826 = 8'h0; 1: mux_11826 = vout_peek_221;
    endcase
  endfunction
  wire [7:0] v_11827;
  function [7:0] mux_11827(input [0:0] sel);
    case (sel) 0: mux_11827 = 8'h0; 1: mux_11827 = vout_peek_213;
    endcase
  endfunction
  wire [7:0] v_11828;
  function [7:0] mux_11828(input [0:0] sel);
    case (sel) 0: mux_11828 = 8'h0; 1: mux_11828 = v_11829;
    endcase
  endfunction
  reg [7:0] v_11829 = 8'h0;
  wire [7:0] v_11830;
  wire [7:0] v_11831;
  function [7:0] mux_11831(input [0:0] sel);
    case (sel) 0: mux_11831 = 8'h0; 1: mux_11831 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11832;
  wire [7:0] v_11833;
  wire [7:0] v_11834;
  function [7:0] mux_11834(input [0:0] sel);
    case (sel) 0: mux_11834 = 8'h0; 1: mux_11834 = vout_peek_207;
    endcase
  endfunction
  wire [7:0] v_11835;
  function [7:0] mux_11835(input [0:0] sel);
    case (sel) 0: mux_11835 = 8'h0; 1: mux_11835 = vout_peek_199;
    endcase
  endfunction
  wire [7:0] v_11836;
  function [7:0] mux_11836(input [0:0] sel);
    case (sel) 0: mux_11836 = 8'h0; 1: mux_11836 = v_11837;
    endcase
  endfunction
  reg [7:0] v_11837 = 8'h0;
  wire [7:0] v_11838;
  wire [7:0] v_11839;
  function [7:0] mux_11839(input [0:0] sel);
    case (sel) 0: mux_11839 = 8'h0; 1: mux_11839 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11840;
  wire [7:0] v_11841;
  wire [7:0] v_11842;
  function [7:0] mux_11842(input [0:0] sel);
    case (sel) 0: mux_11842 = 8'h0; 1: mux_11842 = v_11843;
    endcase
  endfunction
  reg [7:0] v_11843 = 8'h0;
  wire [7:0] v_11844;
  wire [7:0] v_11845;
  function [7:0] mux_11845(input [0:0] sel);
    case (sel) 0: mux_11845 = 8'h0; 1: mux_11845 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11846;
  wire [7:0] v_11847;
  wire [7:0] v_11848;
  function [7:0] mux_11848(input [0:0] sel);
    case (sel) 0: mux_11848 = 8'h0; 1: mux_11848 = vout_peek_193;
    endcase
  endfunction
  wire [7:0] v_11849;
  function [7:0] mux_11849(input [0:0] sel);
    case (sel) 0: mux_11849 = 8'h0; 1: mux_11849 = vout_peek_185;
    endcase
  endfunction
  wire [7:0] v_11850;
  function [7:0] mux_11850(input [0:0] sel);
    case (sel) 0: mux_11850 = 8'h0; 1: mux_11850 = v_11851;
    endcase
  endfunction
  reg [7:0] v_11851 = 8'h0;
  wire [7:0] v_11852;
  wire [7:0] v_11853;
  function [7:0] mux_11853(input [0:0] sel);
    case (sel) 0: mux_11853 = 8'h0; 1: mux_11853 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11854;
  wire [7:0] v_11855;
  wire [7:0] v_11856;
  function [7:0] mux_11856(input [0:0] sel);
    case (sel) 0: mux_11856 = 8'h0; 1: mux_11856 = vout_peek_179;
    endcase
  endfunction
  wire [7:0] v_11857;
  function [7:0] mux_11857(input [0:0] sel);
    case (sel) 0: mux_11857 = 8'h0; 1: mux_11857 = vout_peek_171;
    endcase
  endfunction
  wire [7:0] v_11858;
  function [7:0] mux_11858(input [0:0] sel);
    case (sel) 0: mux_11858 = 8'h0; 1: mux_11858 = v_11859;
    endcase
  endfunction
  reg [7:0] v_11859 = 8'h0;
  wire [7:0] v_11860;
  wire [7:0] v_11861;
  function [7:0] mux_11861(input [0:0] sel);
    case (sel) 0: mux_11861 = 8'h0; 1: mux_11861 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11862;
  wire [7:0] v_11863;
  wire [7:0] v_11864;
  function [7:0] mux_11864(input [0:0] sel);
    case (sel) 0: mux_11864 = 8'h0; 1: mux_11864 = v_11865;
    endcase
  endfunction
  reg [7:0] v_11865 = 8'h0;
  wire [7:0] v_11866;
  wire [7:0] v_11867;
  function [7:0] mux_11867(input [0:0] sel);
    case (sel) 0: mux_11867 = 8'h0; 1: mux_11867 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11868;
  wire [7:0] v_11869;
  wire [7:0] v_11870;
  function [7:0] mux_11870(input [0:0] sel);
    case (sel) 0: mux_11870 = 8'h0; 1: mux_11870 = v_11871;
    endcase
  endfunction
  reg [7:0] v_11871 = 8'h0;
  wire [7:0] v_11872;
  wire [7:0] v_11873;
  function [7:0] mux_11873(input [0:0] sel);
    case (sel) 0: mux_11873 = 8'h0; 1: mux_11873 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11874;
  wire [7:0] v_11875;
  wire [7:0] v_11876;
  function [7:0] mux_11876(input [0:0] sel);
    case (sel) 0: mux_11876 = 8'h0; 1: mux_11876 = vout_peek_165;
    endcase
  endfunction
  wire [7:0] v_11877;
  function [7:0] mux_11877(input [0:0] sel);
    case (sel) 0: mux_11877 = 8'h0; 1: mux_11877 = vout_peek_157;
    endcase
  endfunction
  wire [7:0] v_11878;
  function [7:0] mux_11878(input [0:0] sel);
    case (sel) 0: mux_11878 = 8'h0; 1: mux_11878 = v_11879;
    endcase
  endfunction
  reg [7:0] v_11879 = 8'h0;
  wire [7:0] v_11880;
  wire [7:0] v_11881;
  function [7:0] mux_11881(input [0:0] sel);
    case (sel) 0: mux_11881 = 8'h0; 1: mux_11881 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11882;
  wire [7:0] v_11883;
  wire [7:0] v_11884;
  function [7:0] mux_11884(input [0:0] sel);
    case (sel) 0: mux_11884 = 8'h0; 1: mux_11884 = vout_peek_151;
    endcase
  endfunction
  wire [7:0] v_11885;
  function [7:0] mux_11885(input [0:0] sel);
    case (sel) 0: mux_11885 = 8'h0; 1: mux_11885 = vout_peek_143;
    endcase
  endfunction
  wire [7:0] v_11886;
  function [7:0] mux_11886(input [0:0] sel);
    case (sel) 0: mux_11886 = 8'h0; 1: mux_11886 = v_11887;
    endcase
  endfunction
  reg [7:0] v_11887 = 8'h0;
  wire [7:0] v_11888;
  wire [7:0] v_11889;
  function [7:0] mux_11889(input [0:0] sel);
    case (sel) 0: mux_11889 = 8'h0; 1: mux_11889 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11890;
  wire [7:0] v_11891;
  wire [7:0] v_11892;
  function [7:0] mux_11892(input [0:0] sel);
    case (sel) 0: mux_11892 = 8'h0; 1: mux_11892 = v_11893;
    endcase
  endfunction
  reg [7:0] v_11893 = 8'h0;
  wire [7:0] v_11894;
  wire [7:0] v_11895;
  function [7:0] mux_11895(input [0:0] sel);
    case (sel) 0: mux_11895 = 8'h0; 1: mux_11895 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11896;
  wire [7:0] v_11897;
  wire [7:0] v_11898;
  function [7:0] mux_11898(input [0:0] sel);
    case (sel) 0: mux_11898 = 8'h0; 1: mux_11898 = vout_peek_137;
    endcase
  endfunction
  wire [7:0] v_11899;
  function [7:0] mux_11899(input [0:0] sel);
    case (sel) 0: mux_11899 = 8'h0; 1: mux_11899 = vout_peek_129;
    endcase
  endfunction
  wire [7:0] v_11900;
  function [7:0] mux_11900(input [0:0] sel);
    case (sel) 0: mux_11900 = 8'h0; 1: mux_11900 = v_11901;
    endcase
  endfunction
  reg [7:0] v_11901 = 8'h0;
  wire [7:0] v_11902;
  wire [7:0] v_11903;
  function [7:0] mux_11903(input [0:0] sel);
    case (sel) 0: mux_11903 = 8'h0; 1: mux_11903 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11904;
  wire [7:0] v_11905;
  wire [7:0] v_11906;
  function [7:0] mux_11906(input [0:0] sel);
    case (sel) 0: mux_11906 = 8'h0; 1: mux_11906 = vout_peek_123;
    endcase
  endfunction
  wire [7:0] v_11907;
  function [7:0] mux_11907(input [0:0] sel);
    case (sel) 0: mux_11907 = 8'h0; 1: mux_11907 = vout_peek_115;
    endcase
  endfunction
  wire [7:0] v_11908;
  function [7:0] mux_11908(input [0:0] sel);
    case (sel) 0: mux_11908 = 8'h0; 1: mux_11908 = v_11909;
    endcase
  endfunction
  reg [7:0] v_11909 = 8'h0;
  wire [7:0] v_11910;
  wire [7:0] v_11911;
  function [7:0] mux_11911(input [0:0] sel);
    case (sel) 0: mux_11911 = 8'h0; 1: mux_11911 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11912;
  wire [7:0] v_11913;
  wire [7:0] v_11914;
  function [7:0] mux_11914(input [0:0] sel);
    case (sel) 0: mux_11914 = 8'h0; 1: mux_11914 = v_11915;
    endcase
  endfunction
  reg [7:0] v_11915 = 8'h0;
  wire [7:0] v_11916;
  wire [7:0] v_11917;
  function [7:0] mux_11917(input [0:0] sel);
    case (sel) 0: mux_11917 = 8'h0; 1: mux_11917 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11918;
  wire [7:0] v_11919;
  wire [7:0] v_11920;
  function [7:0] mux_11920(input [0:0] sel);
    case (sel) 0: mux_11920 = 8'h0; 1: mux_11920 = v_11921;
    endcase
  endfunction
  reg [7:0] v_11921 = 8'h0;
  wire [7:0] v_11922;
  wire [7:0] v_11923;
  function [7:0] mux_11923(input [0:0] sel);
    case (sel) 0: mux_11923 = 8'h0; 1: mux_11923 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11924;
  wire [7:0] v_11925;
  wire [7:0] v_11926;
  function [7:0] mux_11926(input [0:0] sel);
    case (sel) 0: mux_11926 = 8'h0; 1: mux_11926 = v_11927;
    endcase
  endfunction
  reg [7:0] v_11927 = 8'h0;
  wire [7:0] v_11928;
  wire [7:0] v_11929;
  function [7:0] mux_11929(input [0:0] sel);
    case (sel) 0: mux_11929 = 8'h0; 1: mux_11929 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11930;
  wire [7:0] v_11931;
  wire [7:0] v_11932;
  function [7:0] mux_11932(input [0:0] sel);
    case (sel) 0: mux_11932 = 8'h0; 1: mux_11932 = vout_peek_109;
    endcase
  endfunction
  wire [7:0] v_11933;
  function [7:0] mux_11933(input [0:0] sel);
    case (sel) 0: mux_11933 = 8'h0; 1: mux_11933 = vout_peek_101;
    endcase
  endfunction
  wire [7:0] v_11934;
  function [7:0] mux_11934(input [0:0] sel);
    case (sel) 0: mux_11934 = 8'h0; 1: mux_11934 = v_11935;
    endcase
  endfunction
  reg [7:0] v_11935 = 8'h0;
  wire [7:0] v_11936;
  wire [7:0] v_11937;
  function [7:0] mux_11937(input [0:0] sel);
    case (sel) 0: mux_11937 = 8'h0; 1: mux_11937 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11938;
  wire [7:0] v_11939;
  wire [7:0] v_11940;
  function [7:0] mux_11940(input [0:0] sel);
    case (sel) 0: mux_11940 = 8'h0; 1: mux_11940 = vout_peek_95;
    endcase
  endfunction
  wire [7:0] v_11941;
  function [7:0] mux_11941(input [0:0] sel);
    case (sel) 0: mux_11941 = 8'h0; 1: mux_11941 = vout_peek_87;
    endcase
  endfunction
  wire [7:0] v_11942;
  function [7:0] mux_11942(input [0:0] sel);
    case (sel) 0: mux_11942 = 8'h0; 1: mux_11942 = v_11943;
    endcase
  endfunction
  reg [7:0] v_11943 = 8'h0;
  wire [7:0] v_11944;
  wire [7:0] v_11945;
  function [7:0] mux_11945(input [0:0] sel);
    case (sel) 0: mux_11945 = 8'h0; 1: mux_11945 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11946;
  wire [7:0] v_11947;
  wire [7:0] v_11948;
  function [7:0] mux_11948(input [0:0] sel);
    case (sel) 0: mux_11948 = 8'h0; 1: mux_11948 = v_11949;
    endcase
  endfunction
  reg [7:0] v_11949 = 8'h0;
  wire [7:0] v_11950;
  wire [7:0] v_11951;
  function [7:0] mux_11951(input [0:0] sel);
    case (sel) 0: mux_11951 = 8'h0; 1: mux_11951 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11952;
  wire [7:0] v_11953;
  wire [7:0] v_11954;
  function [7:0] mux_11954(input [0:0] sel);
    case (sel) 0: mux_11954 = 8'h0; 1: mux_11954 = vout_peek_81;
    endcase
  endfunction
  wire [7:0] v_11955;
  function [7:0] mux_11955(input [0:0] sel);
    case (sel) 0: mux_11955 = 8'h0; 1: mux_11955 = vout_peek_73;
    endcase
  endfunction
  wire [7:0] v_11956;
  function [7:0] mux_11956(input [0:0] sel);
    case (sel) 0: mux_11956 = 8'h0; 1: mux_11956 = v_11957;
    endcase
  endfunction
  reg [7:0] v_11957 = 8'h0;
  wire [7:0] v_11958;
  wire [7:0] v_11959;
  function [7:0] mux_11959(input [0:0] sel);
    case (sel) 0: mux_11959 = 8'h0; 1: mux_11959 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11960;
  wire [7:0] v_11961;
  wire [7:0] v_11962;
  function [7:0] mux_11962(input [0:0] sel);
    case (sel) 0: mux_11962 = 8'h0; 1: mux_11962 = vout_peek_67;
    endcase
  endfunction
  wire [7:0] v_11963;
  function [7:0] mux_11963(input [0:0] sel);
    case (sel) 0: mux_11963 = 8'h0; 1: mux_11963 = vout_peek_59;
    endcase
  endfunction
  wire [7:0] v_11964;
  function [7:0] mux_11964(input [0:0] sel);
    case (sel) 0: mux_11964 = 8'h0; 1: mux_11964 = v_11965;
    endcase
  endfunction
  reg [7:0] v_11965 = 8'h0;
  wire [7:0] v_11966;
  wire [7:0] v_11967;
  function [7:0] mux_11967(input [0:0] sel);
    case (sel) 0: mux_11967 = 8'h0; 1: mux_11967 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11968;
  wire [7:0] v_11969;
  wire [7:0] v_11970;
  function [7:0] mux_11970(input [0:0] sel);
    case (sel) 0: mux_11970 = 8'h0; 1: mux_11970 = v_11971;
    endcase
  endfunction
  reg [7:0] v_11971 = 8'h0;
  wire [7:0] v_11972;
  wire [7:0] v_11973;
  function [7:0] mux_11973(input [0:0] sel);
    case (sel) 0: mux_11973 = 8'h0; 1: mux_11973 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11974;
  wire [7:0] v_11975;
  wire [7:0] v_11976;
  function [7:0] mux_11976(input [0:0] sel);
    case (sel) 0: mux_11976 = 8'h0; 1: mux_11976 = v_11977;
    endcase
  endfunction
  reg [7:0] v_11977 = 8'h0;
  wire [7:0] v_11978;
  wire [7:0] v_11979;
  function [7:0] mux_11979(input [0:0] sel);
    case (sel) 0: mux_11979 = 8'h0; 1: mux_11979 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11980;
  wire [7:0] v_11981;
  wire [7:0] v_11982;
  function [7:0] mux_11982(input [0:0] sel);
    case (sel) 0: mux_11982 = 8'h0; 1: mux_11982 = vout_peek_53;
    endcase
  endfunction
  wire [7:0] v_11983;
  function [7:0] mux_11983(input [0:0] sel);
    case (sel) 0: mux_11983 = 8'h0; 1: mux_11983 = vout_peek_45;
    endcase
  endfunction
  wire [7:0] v_11984;
  function [7:0] mux_11984(input [0:0] sel);
    case (sel) 0: mux_11984 = 8'h0; 1: mux_11984 = v_11985;
    endcase
  endfunction
  reg [7:0] v_11985 = 8'h0;
  wire [7:0] v_11986;
  wire [7:0] v_11987;
  function [7:0] mux_11987(input [0:0] sel);
    case (sel) 0: mux_11987 = 8'h0; 1: mux_11987 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11988;
  wire [7:0] v_11989;
  wire [7:0] v_11990;
  function [7:0] mux_11990(input [0:0] sel);
    case (sel) 0: mux_11990 = 8'h0; 1: mux_11990 = vout_peek_39;
    endcase
  endfunction
  wire [7:0] v_11991;
  function [7:0] mux_11991(input [0:0] sel);
    case (sel) 0: mux_11991 = 8'h0; 1: mux_11991 = vout_peek_31;
    endcase
  endfunction
  wire [7:0] v_11992;
  function [7:0] mux_11992(input [0:0] sel);
    case (sel) 0: mux_11992 = 8'h0; 1: mux_11992 = v_11993;
    endcase
  endfunction
  reg [7:0] v_11993 = 8'h0;
  wire [7:0] v_11994;
  wire [7:0] v_11995;
  function [7:0] mux_11995(input [0:0] sel);
    case (sel) 0: mux_11995 = 8'h0; 1: mux_11995 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_11996;
  wire [7:0] v_11997;
  wire [7:0] v_11998;
  function [7:0] mux_11998(input [0:0] sel);
    case (sel) 0: mux_11998 = 8'h0; 1: mux_11998 = v_11999;
    endcase
  endfunction
  reg [7:0] v_11999 = 8'h0;
  wire [7:0] v_12000;
  wire [7:0] v_12001;
  function [7:0] mux_12001(input [0:0] sel);
    case (sel) 0: mux_12001 = 8'h0; 1: mux_12001 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12002;
  wire [7:0] v_12003;
  wire [7:0] v_12004;
  function [7:0] mux_12004(input [0:0] sel);
    case (sel) 0: mux_12004 = 8'h0; 1: mux_12004 = vout_peek_25;
    endcase
  endfunction
  wire [7:0] v_12005;
  function [7:0] mux_12005(input [0:0] sel);
    case (sel) 0: mux_12005 = 8'h0; 1: mux_12005 = vout_peek_17;
    endcase
  endfunction
  wire [7:0] v_12006;
  function [7:0] mux_12006(input [0:0] sel);
    case (sel) 0: mux_12006 = 8'h0; 1: mux_12006 = v_12007;
    endcase
  endfunction
  reg [7:0] v_12007 = 8'h0;
  wire [7:0] v_12008;
  wire [7:0] v_12009;
  function [7:0] mux_12009(input [0:0] sel);
    case (sel) 0: mux_12009 = 8'h0; 1: mux_12009 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12010;
  wire [7:0] v_12011;
  wire [7:0] v_12012;
  function [7:0] mux_12012(input [0:0] sel);
    case (sel) 0: mux_12012 = 8'h0; 1: mux_12012 = vout_peek_11;
    endcase
  endfunction
  wire [7:0] v_12013;
  function [7:0] mux_12013(input [0:0] sel);
    case (sel) 0: mux_12013 = 8'h0; 1: mux_12013 = vout_peek_3;
    endcase
  endfunction
  wire [7:0] v_12014;
  function [7:0] mux_12014(input [0:0] sel);
    case (sel) 0: mux_12014 = 8'h0; 1: mux_12014 = v_12015;
    endcase
  endfunction
  reg [7:0] v_12015 = 8'h0;
  wire [7:0] v_12016;
  wire [7:0] v_12017;
  function [7:0] mux_12017(input [0:0] sel);
    case (sel) 0: mux_12017 = 8'h0; 1: mux_12017 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12018;
  wire [7:0] v_12019;
  wire [7:0] v_12020;
  function [7:0] mux_12020(input [0:0] sel);
    case (sel) 0: mux_12020 = 8'h0; 1: mux_12020 = v_12021;
    endcase
  endfunction
  reg [7:0] v_12021 = 8'h0;
  wire [7:0] v_12022;
  wire [7:0] v_12023;
  function [7:0] mux_12023(input [0:0] sel);
    case (sel) 0: mux_12023 = 8'h0; 1: mux_12023 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12024;
  wire [7:0] v_12025;
  wire [7:0] v_12026;
  function [7:0] mux_12026(input [0:0] sel);
    case (sel) 0: mux_12026 = 8'h0; 1: mux_12026 = v_12027;
    endcase
  endfunction
  reg [7:0] v_12027 = 8'h0;
  wire [7:0] v_12028;
  wire [7:0] v_12029;
  function [7:0] mux_12029(input [0:0] sel);
    case (sel) 0: mux_12029 = 8'h0; 1: mux_12029 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12030;
  wire [7:0] v_12031;
  wire [7:0] v_12032;
  function [7:0] mux_12032(input [0:0] sel);
    case (sel) 0: mux_12032 = 8'h0; 1: mux_12032 = v_12033;
    endcase
  endfunction
  reg [7:0] v_12033 = 8'h0;
  wire [7:0] v_12034;
  wire [7:0] v_12035;
  function [7:0] mux_12035(input [0:0] sel);
    case (sel) 0: mux_12035 = 8'h0; 1: mux_12035 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12036;
  wire [7:0] v_12037;
  wire [7:0] v_12038;
  function [7:0] mux_12038(input [0:0] sel);
    case (sel) 0: mux_12038 = 8'h0; 1: mux_12038 = vout_peek_2797;
    endcase
  endfunction
  wire [7:0] v_12039;
  function [7:0] mux_12039(input [0:0] sel);
    case (sel) 0: mux_12039 = 8'h0; 1: mux_12039 = vout_peek_2789;
    endcase
  endfunction
  wire [7:0] v_12040;
  function [7:0] mux_12040(input [0:0] sel);
    case (sel) 0: mux_12040 = 8'h0; 1: mux_12040 = v_12041;
    endcase
  endfunction
  reg [7:0] v_12041 = 8'h0;
  wire [7:0] v_12042;
  wire [7:0] v_12043;
  function [7:0] mux_12043(input [0:0] sel);
    case (sel) 0: mux_12043 = 8'h0; 1: mux_12043 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12044;
  wire [7:0] v_12045;
  wire [7:0] v_12046;
  function [7:0] mux_12046(input [0:0] sel);
    case (sel) 0: mux_12046 = 8'h0; 1: mux_12046 = vout_peek_2783;
    endcase
  endfunction
  wire [7:0] v_12047;
  function [7:0] mux_12047(input [0:0] sel);
    case (sel) 0: mux_12047 = 8'h0; 1: mux_12047 = vout_peek_2775;
    endcase
  endfunction
  wire [7:0] v_12048;
  function [7:0] mux_12048(input [0:0] sel);
    case (sel) 0: mux_12048 = 8'h0; 1: mux_12048 = v_12049;
    endcase
  endfunction
  reg [7:0] v_12049 = 8'h0;
  wire [7:0] v_12050;
  wire [7:0] v_12051;
  function [7:0] mux_12051(input [0:0] sel);
    case (sel) 0: mux_12051 = 8'h0; 1: mux_12051 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12052;
  wire [7:0] v_12053;
  wire [7:0] v_12054;
  function [7:0] mux_12054(input [0:0] sel);
    case (sel) 0: mux_12054 = 8'h0; 1: mux_12054 = v_12055;
    endcase
  endfunction
  reg [7:0] v_12055 = 8'h0;
  wire [7:0] v_12056;
  wire [7:0] v_12057;
  function [7:0] mux_12057(input [0:0] sel);
    case (sel) 0: mux_12057 = 8'h0; 1: mux_12057 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12058;
  wire [7:0] v_12059;
  wire [7:0] v_12060;
  function [7:0] mux_12060(input [0:0] sel);
    case (sel) 0: mux_12060 = 8'h0; 1: mux_12060 = vout_peek_2769;
    endcase
  endfunction
  wire [7:0] v_12061;
  function [7:0] mux_12061(input [0:0] sel);
    case (sel) 0: mux_12061 = 8'h0; 1: mux_12061 = vout_peek_2761;
    endcase
  endfunction
  wire [7:0] v_12062;
  function [7:0] mux_12062(input [0:0] sel);
    case (sel) 0: mux_12062 = 8'h0; 1: mux_12062 = v_12063;
    endcase
  endfunction
  reg [7:0] v_12063 = 8'h0;
  wire [7:0] v_12064;
  wire [7:0] v_12065;
  function [7:0] mux_12065(input [0:0] sel);
    case (sel) 0: mux_12065 = 8'h0; 1: mux_12065 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12066;
  wire [7:0] v_12067;
  wire [7:0] v_12068;
  function [7:0] mux_12068(input [0:0] sel);
    case (sel) 0: mux_12068 = 8'h0; 1: mux_12068 = vout_peek_2755;
    endcase
  endfunction
  wire [7:0] v_12069;
  function [7:0] mux_12069(input [0:0] sel);
    case (sel) 0: mux_12069 = 8'h0; 1: mux_12069 = vout_peek_2747;
    endcase
  endfunction
  wire [7:0] v_12070;
  function [7:0] mux_12070(input [0:0] sel);
    case (sel) 0: mux_12070 = 8'h0; 1: mux_12070 = v_12071;
    endcase
  endfunction
  reg [7:0] v_12071 = 8'h0;
  wire [7:0] v_12072;
  wire [7:0] v_12073;
  function [7:0] mux_12073(input [0:0] sel);
    case (sel) 0: mux_12073 = 8'h0; 1: mux_12073 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12074;
  wire [7:0] v_12075;
  wire [7:0] v_12076;
  function [7:0] mux_12076(input [0:0] sel);
    case (sel) 0: mux_12076 = 8'h0; 1: mux_12076 = v_12077;
    endcase
  endfunction
  reg [7:0] v_12077 = 8'h0;
  wire [7:0] v_12078;
  wire [7:0] v_12079;
  function [7:0] mux_12079(input [0:0] sel);
    case (sel) 0: mux_12079 = 8'h0; 1: mux_12079 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12080;
  wire [7:0] v_12081;
  wire [7:0] v_12082;
  function [7:0] mux_12082(input [0:0] sel);
    case (sel) 0: mux_12082 = 8'h0; 1: mux_12082 = v_12083;
    endcase
  endfunction
  reg [7:0] v_12083 = 8'h0;
  wire [7:0] v_12084;
  wire [7:0] v_12085;
  function [7:0] mux_12085(input [0:0] sel);
    case (sel) 0: mux_12085 = 8'h0; 1: mux_12085 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12086;
  wire [7:0] v_12087;
  wire [7:0] v_12088;
  function [7:0] mux_12088(input [0:0] sel);
    case (sel) 0: mux_12088 = 8'h0; 1: mux_12088 = vout_peek_2741;
    endcase
  endfunction
  wire [7:0] v_12089;
  function [7:0] mux_12089(input [0:0] sel);
    case (sel) 0: mux_12089 = 8'h0; 1: mux_12089 = vout_peek_2733;
    endcase
  endfunction
  wire [7:0] v_12090;
  function [7:0] mux_12090(input [0:0] sel);
    case (sel) 0: mux_12090 = 8'h0; 1: mux_12090 = v_12091;
    endcase
  endfunction
  reg [7:0] v_12091 = 8'h0;
  wire [7:0] v_12092;
  wire [7:0] v_12093;
  function [7:0] mux_12093(input [0:0] sel);
    case (sel) 0: mux_12093 = 8'h0; 1: mux_12093 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12094;
  wire [7:0] v_12095;
  wire [7:0] v_12096;
  function [7:0] mux_12096(input [0:0] sel);
    case (sel) 0: mux_12096 = 8'h0; 1: mux_12096 = vout_peek_2727;
    endcase
  endfunction
  wire [7:0] v_12097;
  function [7:0] mux_12097(input [0:0] sel);
    case (sel) 0: mux_12097 = 8'h0; 1: mux_12097 = vout_peek_2719;
    endcase
  endfunction
  wire [7:0] v_12098;
  function [7:0] mux_12098(input [0:0] sel);
    case (sel) 0: mux_12098 = 8'h0; 1: mux_12098 = v_12099;
    endcase
  endfunction
  reg [7:0] v_12099 = 8'h0;
  wire [7:0] v_12100;
  wire [7:0] v_12101;
  function [7:0] mux_12101(input [0:0] sel);
    case (sel) 0: mux_12101 = 8'h0; 1: mux_12101 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12102;
  wire [7:0] v_12103;
  wire [7:0] v_12104;
  function [7:0] mux_12104(input [0:0] sel);
    case (sel) 0: mux_12104 = 8'h0; 1: mux_12104 = v_12105;
    endcase
  endfunction
  reg [7:0] v_12105 = 8'h0;
  wire [7:0] v_12106;
  wire [7:0] v_12107;
  function [7:0] mux_12107(input [0:0] sel);
    case (sel) 0: mux_12107 = 8'h0; 1: mux_12107 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12108;
  wire [7:0] v_12109;
  wire [7:0] v_12110;
  function [7:0] mux_12110(input [0:0] sel);
    case (sel) 0: mux_12110 = 8'h0; 1: mux_12110 = vout_peek_2713;
    endcase
  endfunction
  wire [7:0] v_12111;
  function [7:0] mux_12111(input [0:0] sel);
    case (sel) 0: mux_12111 = 8'h0; 1: mux_12111 = vout_peek_2705;
    endcase
  endfunction
  wire [7:0] v_12112;
  function [7:0] mux_12112(input [0:0] sel);
    case (sel) 0: mux_12112 = 8'h0; 1: mux_12112 = v_12113;
    endcase
  endfunction
  reg [7:0] v_12113 = 8'h0;
  wire [7:0] v_12114;
  wire [7:0] v_12115;
  function [7:0] mux_12115(input [0:0] sel);
    case (sel) 0: mux_12115 = 8'h0; 1: mux_12115 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12116;
  wire [7:0] v_12117;
  wire [7:0] v_12118;
  function [7:0] mux_12118(input [0:0] sel);
    case (sel) 0: mux_12118 = 8'h0; 1: mux_12118 = vout_peek_2699;
    endcase
  endfunction
  wire [7:0] v_12119;
  function [7:0] mux_12119(input [0:0] sel);
    case (sel) 0: mux_12119 = 8'h0; 1: mux_12119 = vout_peek_2691;
    endcase
  endfunction
  wire [7:0] v_12120;
  function [7:0] mux_12120(input [0:0] sel);
    case (sel) 0: mux_12120 = 8'h0; 1: mux_12120 = v_12121;
    endcase
  endfunction
  reg [7:0] v_12121 = 8'h0;
  wire [7:0] v_12122;
  wire [7:0] v_12123;
  function [7:0] mux_12123(input [0:0] sel);
    case (sel) 0: mux_12123 = 8'h0; 1: mux_12123 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12124;
  wire [7:0] v_12125;
  wire [7:0] v_12126;
  function [7:0] mux_12126(input [0:0] sel);
    case (sel) 0: mux_12126 = 8'h0; 1: mux_12126 = v_12127;
    endcase
  endfunction
  reg [7:0] v_12127 = 8'h0;
  wire [7:0] v_12128;
  wire [7:0] v_12129;
  function [7:0] mux_12129(input [0:0] sel);
    case (sel) 0: mux_12129 = 8'h0; 1: mux_12129 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12130;
  wire [7:0] v_12131;
  wire [7:0] v_12132;
  function [7:0] mux_12132(input [0:0] sel);
    case (sel) 0: mux_12132 = 8'h0; 1: mux_12132 = v_12133;
    endcase
  endfunction
  reg [7:0] v_12133 = 8'h0;
  wire [7:0] v_12134;
  wire [7:0] v_12135;
  function [7:0] mux_12135(input [0:0] sel);
    case (sel) 0: mux_12135 = 8'h0; 1: mux_12135 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12136;
  wire [7:0] v_12137;
  wire [7:0] v_12138;
  function [7:0] mux_12138(input [0:0] sel);
    case (sel) 0: mux_12138 = 8'h0; 1: mux_12138 = v_12139;
    endcase
  endfunction
  reg [7:0] v_12139 = 8'h0;
  wire [7:0] v_12140;
  wire [7:0] v_12141;
  function [7:0] mux_12141(input [0:0] sel);
    case (sel) 0: mux_12141 = 8'h0; 1: mux_12141 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12142;
  wire [7:0] v_12143;
  wire [7:0] v_12144;
  function [7:0] mux_12144(input [0:0] sel);
    case (sel) 0: mux_12144 = 8'h0; 1: mux_12144 = v_12145;
    endcase
  endfunction
  reg [7:0] v_12145 = 8'h0;
  wire [7:0] v_12146;
  wire [7:0] v_12147;
  function [7:0] mux_12147(input [0:0] sel);
    case (sel) 0: mux_12147 = 8'h0; 1: mux_12147 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12148;
  wire [7:0] v_12149;
  wire [7:0] v_12150;
  function [7:0] mux_12150(input [0:0] sel);
    case (sel) 0: mux_12150 = 8'h0; 1: mux_12150 = vout_peek_2685;
    endcase
  endfunction
  wire [7:0] v_12151;
  function [7:0] mux_12151(input [0:0] sel);
    case (sel) 0: mux_12151 = 8'h0; 1: mux_12151 = vout_peek_2677;
    endcase
  endfunction
  wire [7:0] v_12152;
  function [7:0] mux_12152(input [0:0] sel);
    case (sel) 0: mux_12152 = 8'h0; 1: mux_12152 = v_12153;
    endcase
  endfunction
  reg [7:0] v_12153 = 8'h0;
  wire [7:0] v_12154;
  wire [7:0] v_12155;
  function [7:0] mux_12155(input [0:0] sel);
    case (sel) 0: mux_12155 = 8'h0; 1: mux_12155 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12156;
  wire [7:0] v_12157;
  wire [7:0] v_12158;
  function [7:0] mux_12158(input [0:0] sel);
    case (sel) 0: mux_12158 = 8'h0; 1: mux_12158 = vout_peek_2671;
    endcase
  endfunction
  wire [7:0] v_12159;
  function [7:0] mux_12159(input [0:0] sel);
    case (sel) 0: mux_12159 = 8'h0; 1: mux_12159 = vout_peek_2663;
    endcase
  endfunction
  wire [7:0] v_12160;
  function [7:0] mux_12160(input [0:0] sel);
    case (sel) 0: mux_12160 = 8'h0; 1: mux_12160 = v_12161;
    endcase
  endfunction
  reg [7:0] v_12161 = 8'h0;
  wire [7:0] v_12162;
  wire [7:0] v_12163;
  function [7:0] mux_12163(input [0:0] sel);
    case (sel) 0: mux_12163 = 8'h0; 1: mux_12163 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12164;
  wire [7:0] v_12165;
  wire [7:0] v_12166;
  function [7:0] mux_12166(input [0:0] sel);
    case (sel) 0: mux_12166 = 8'h0; 1: mux_12166 = v_12167;
    endcase
  endfunction
  reg [7:0] v_12167 = 8'h0;
  wire [7:0] v_12168;
  wire [7:0] v_12169;
  function [7:0] mux_12169(input [0:0] sel);
    case (sel) 0: mux_12169 = 8'h0; 1: mux_12169 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12170;
  wire [7:0] v_12171;
  wire [7:0] v_12172;
  function [7:0] mux_12172(input [0:0] sel);
    case (sel) 0: mux_12172 = 8'h0; 1: mux_12172 = vout_peek_2657;
    endcase
  endfunction
  wire [7:0] v_12173;
  function [7:0] mux_12173(input [0:0] sel);
    case (sel) 0: mux_12173 = 8'h0; 1: mux_12173 = vout_peek_2649;
    endcase
  endfunction
  wire [7:0] v_12174;
  function [7:0] mux_12174(input [0:0] sel);
    case (sel) 0: mux_12174 = 8'h0; 1: mux_12174 = v_12175;
    endcase
  endfunction
  reg [7:0] v_12175 = 8'h0;
  wire [7:0] v_12176;
  wire [7:0] v_12177;
  function [7:0] mux_12177(input [0:0] sel);
    case (sel) 0: mux_12177 = 8'h0; 1: mux_12177 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12178;
  wire [7:0] v_12179;
  wire [7:0] v_12180;
  function [7:0] mux_12180(input [0:0] sel);
    case (sel) 0: mux_12180 = 8'h0; 1: mux_12180 = vout_peek_2643;
    endcase
  endfunction
  wire [7:0] v_12181;
  function [7:0] mux_12181(input [0:0] sel);
    case (sel) 0: mux_12181 = 8'h0; 1: mux_12181 = vout_peek_2635;
    endcase
  endfunction
  wire [7:0] v_12182;
  function [7:0] mux_12182(input [0:0] sel);
    case (sel) 0: mux_12182 = 8'h0; 1: mux_12182 = v_12183;
    endcase
  endfunction
  reg [7:0] v_12183 = 8'h0;
  wire [7:0] v_12184;
  wire [7:0] v_12185;
  function [7:0] mux_12185(input [0:0] sel);
    case (sel) 0: mux_12185 = 8'h0; 1: mux_12185 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12186;
  wire [7:0] v_12187;
  wire [7:0] v_12188;
  function [7:0] mux_12188(input [0:0] sel);
    case (sel) 0: mux_12188 = 8'h0; 1: mux_12188 = v_12189;
    endcase
  endfunction
  reg [7:0] v_12189 = 8'h0;
  wire [7:0] v_12190;
  wire [7:0] v_12191;
  function [7:0] mux_12191(input [0:0] sel);
    case (sel) 0: mux_12191 = 8'h0; 1: mux_12191 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12192;
  wire [7:0] v_12193;
  wire [7:0] v_12194;
  function [7:0] mux_12194(input [0:0] sel);
    case (sel) 0: mux_12194 = 8'h0; 1: mux_12194 = v_12195;
    endcase
  endfunction
  reg [7:0] v_12195 = 8'h0;
  wire [7:0] v_12196;
  wire [7:0] v_12197;
  function [7:0] mux_12197(input [0:0] sel);
    case (sel) 0: mux_12197 = 8'h0; 1: mux_12197 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12198;
  wire [7:0] v_12199;
  wire [7:0] v_12200;
  function [7:0] mux_12200(input [0:0] sel);
    case (sel) 0: mux_12200 = 8'h0; 1: mux_12200 = vout_peek_2629;
    endcase
  endfunction
  wire [7:0] v_12201;
  function [7:0] mux_12201(input [0:0] sel);
    case (sel) 0: mux_12201 = 8'h0; 1: mux_12201 = vout_peek_2621;
    endcase
  endfunction
  wire [7:0] v_12202;
  function [7:0] mux_12202(input [0:0] sel);
    case (sel) 0: mux_12202 = 8'h0; 1: mux_12202 = v_12203;
    endcase
  endfunction
  reg [7:0] v_12203 = 8'h0;
  wire [7:0] v_12204;
  wire [7:0] v_12205;
  function [7:0] mux_12205(input [0:0] sel);
    case (sel) 0: mux_12205 = 8'h0; 1: mux_12205 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12206;
  wire [7:0] v_12207;
  wire [7:0] v_12208;
  function [7:0] mux_12208(input [0:0] sel);
    case (sel) 0: mux_12208 = 8'h0; 1: mux_12208 = vout_peek_2615;
    endcase
  endfunction
  wire [7:0] v_12209;
  function [7:0] mux_12209(input [0:0] sel);
    case (sel) 0: mux_12209 = 8'h0; 1: mux_12209 = vout_peek_2607;
    endcase
  endfunction
  wire [7:0] v_12210;
  function [7:0] mux_12210(input [0:0] sel);
    case (sel) 0: mux_12210 = 8'h0; 1: mux_12210 = v_12211;
    endcase
  endfunction
  reg [7:0] v_12211 = 8'h0;
  wire [7:0] v_12212;
  wire [7:0] v_12213;
  function [7:0] mux_12213(input [0:0] sel);
    case (sel) 0: mux_12213 = 8'h0; 1: mux_12213 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12214;
  wire [7:0] v_12215;
  wire [7:0] v_12216;
  function [7:0] mux_12216(input [0:0] sel);
    case (sel) 0: mux_12216 = 8'h0; 1: mux_12216 = v_12217;
    endcase
  endfunction
  reg [7:0] v_12217 = 8'h0;
  wire [7:0] v_12218;
  wire [7:0] v_12219;
  function [7:0] mux_12219(input [0:0] sel);
    case (sel) 0: mux_12219 = 8'h0; 1: mux_12219 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12220;
  wire [7:0] v_12221;
  wire [7:0] v_12222;
  function [7:0] mux_12222(input [0:0] sel);
    case (sel) 0: mux_12222 = 8'h0; 1: mux_12222 = vout_peek_2601;
    endcase
  endfunction
  wire [7:0] v_12223;
  function [7:0] mux_12223(input [0:0] sel);
    case (sel) 0: mux_12223 = 8'h0; 1: mux_12223 = vout_peek_2593;
    endcase
  endfunction
  wire [7:0] v_12224;
  function [7:0] mux_12224(input [0:0] sel);
    case (sel) 0: mux_12224 = 8'h0; 1: mux_12224 = v_12225;
    endcase
  endfunction
  reg [7:0] v_12225 = 8'h0;
  wire [7:0] v_12226;
  wire [7:0] v_12227;
  function [7:0] mux_12227(input [0:0] sel);
    case (sel) 0: mux_12227 = 8'h0; 1: mux_12227 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12228;
  wire [7:0] v_12229;
  wire [7:0] v_12230;
  function [7:0] mux_12230(input [0:0] sel);
    case (sel) 0: mux_12230 = 8'h0; 1: mux_12230 = vout_peek_2587;
    endcase
  endfunction
  wire [7:0] v_12231;
  function [7:0] mux_12231(input [0:0] sel);
    case (sel) 0: mux_12231 = 8'h0; 1: mux_12231 = vout_peek_2579;
    endcase
  endfunction
  wire [7:0] v_12232;
  function [7:0] mux_12232(input [0:0] sel);
    case (sel) 0: mux_12232 = 8'h0; 1: mux_12232 = v_12233;
    endcase
  endfunction
  reg [7:0] v_12233 = 8'h0;
  wire [7:0] v_12234;
  wire [7:0] v_12235;
  function [7:0] mux_12235(input [0:0] sel);
    case (sel) 0: mux_12235 = 8'h0; 1: mux_12235 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12236;
  wire [7:0] v_12237;
  wire [7:0] v_12238;
  function [7:0] mux_12238(input [0:0] sel);
    case (sel) 0: mux_12238 = 8'h0; 1: mux_12238 = v_12239;
    endcase
  endfunction
  reg [7:0] v_12239 = 8'h0;
  wire [7:0] v_12240;
  wire [7:0] v_12241;
  function [7:0] mux_12241(input [0:0] sel);
    case (sel) 0: mux_12241 = 8'h0; 1: mux_12241 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12242;
  wire [7:0] v_12243;
  wire [7:0] v_12244;
  function [7:0] mux_12244(input [0:0] sel);
    case (sel) 0: mux_12244 = 8'h0; 1: mux_12244 = v_12245;
    endcase
  endfunction
  reg [7:0] v_12245 = 8'h0;
  wire [7:0] v_12246;
  wire [7:0] v_12247;
  function [7:0] mux_12247(input [0:0] sel);
    case (sel) 0: mux_12247 = 8'h0; 1: mux_12247 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12248;
  wire [7:0] v_12249;
  wire [7:0] v_12250;
  function [7:0] mux_12250(input [0:0] sel);
    case (sel) 0: mux_12250 = 8'h0; 1: mux_12250 = v_12251;
    endcase
  endfunction
  reg [7:0] v_12251 = 8'h0;
  wire [7:0] v_12252;
  wire [7:0] v_12253;
  function [7:0] mux_12253(input [0:0] sel);
    case (sel) 0: mux_12253 = 8'h0; 1: mux_12253 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12254;
  wire [7:0] v_12255;
  wire [7:0] v_12256;
  function [7:0] mux_12256(input [0:0] sel);
    case (sel) 0: mux_12256 = 8'h0; 1: mux_12256 = vout_peek_2573;
    endcase
  endfunction
  wire [7:0] v_12257;
  function [7:0] mux_12257(input [0:0] sel);
    case (sel) 0: mux_12257 = 8'h0; 1: mux_12257 = vout_peek_2565;
    endcase
  endfunction
  wire [7:0] v_12258;
  function [7:0] mux_12258(input [0:0] sel);
    case (sel) 0: mux_12258 = 8'h0; 1: mux_12258 = v_12259;
    endcase
  endfunction
  reg [7:0] v_12259 = 8'h0;
  wire [7:0] v_12260;
  wire [7:0] v_12261;
  function [7:0] mux_12261(input [0:0] sel);
    case (sel) 0: mux_12261 = 8'h0; 1: mux_12261 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12262;
  wire [7:0] v_12263;
  wire [7:0] v_12264;
  function [7:0] mux_12264(input [0:0] sel);
    case (sel) 0: mux_12264 = 8'h0; 1: mux_12264 = vout_peek_2559;
    endcase
  endfunction
  wire [7:0] v_12265;
  function [7:0] mux_12265(input [0:0] sel);
    case (sel) 0: mux_12265 = 8'h0; 1: mux_12265 = vout_peek_2551;
    endcase
  endfunction
  wire [7:0] v_12266;
  function [7:0] mux_12266(input [0:0] sel);
    case (sel) 0: mux_12266 = 8'h0; 1: mux_12266 = v_12267;
    endcase
  endfunction
  reg [7:0] v_12267 = 8'h0;
  wire [7:0] v_12268;
  wire [7:0] v_12269;
  function [7:0] mux_12269(input [0:0] sel);
    case (sel) 0: mux_12269 = 8'h0; 1: mux_12269 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12270;
  wire [7:0] v_12271;
  wire [7:0] v_12272;
  function [7:0] mux_12272(input [0:0] sel);
    case (sel) 0: mux_12272 = 8'h0; 1: mux_12272 = v_12273;
    endcase
  endfunction
  reg [7:0] v_12273 = 8'h0;
  wire [7:0] v_12274;
  wire [7:0] v_12275;
  function [7:0] mux_12275(input [0:0] sel);
    case (sel) 0: mux_12275 = 8'h0; 1: mux_12275 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12276;
  wire [7:0] v_12277;
  wire [7:0] v_12278;
  function [7:0] mux_12278(input [0:0] sel);
    case (sel) 0: mux_12278 = 8'h0; 1: mux_12278 = vout_peek_2545;
    endcase
  endfunction
  wire [7:0] v_12279;
  function [7:0] mux_12279(input [0:0] sel);
    case (sel) 0: mux_12279 = 8'h0; 1: mux_12279 = vout_peek_2537;
    endcase
  endfunction
  wire [7:0] v_12280;
  function [7:0] mux_12280(input [0:0] sel);
    case (sel) 0: mux_12280 = 8'h0; 1: mux_12280 = v_12281;
    endcase
  endfunction
  reg [7:0] v_12281 = 8'h0;
  wire [7:0] v_12282;
  wire [7:0] v_12283;
  function [7:0] mux_12283(input [0:0] sel);
    case (sel) 0: mux_12283 = 8'h0; 1: mux_12283 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12284;
  wire [7:0] v_12285;
  wire [7:0] v_12286;
  function [7:0] mux_12286(input [0:0] sel);
    case (sel) 0: mux_12286 = 8'h0; 1: mux_12286 = vout_peek_2531;
    endcase
  endfunction
  wire [7:0] v_12287;
  function [7:0] mux_12287(input [0:0] sel);
    case (sel) 0: mux_12287 = 8'h0; 1: mux_12287 = vout_peek_2523;
    endcase
  endfunction
  wire [7:0] v_12288;
  function [7:0] mux_12288(input [0:0] sel);
    case (sel) 0: mux_12288 = 8'h0; 1: mux_12288 = v_12289;
    endcase
  endfunction
  reg [7:0] v_12289 = 8'h0;
  wire [7:0] v_12290;
  wire [7:0] v_12291;
  function [7:0] mux_12291(input [0:0] sel);
    case (sel) 0: mux_12291 = 8'h0; 1: mux_12291 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12292;
  wire [7:0] v_12293;
  wire [7:0] v_12294;
  function [7:0] mux_12294(input [0:0] sel);
    case (sel) 0: mux_12294 = 8'h0; 1: mux_12294 = v_12295;
    endcase
  endfunction
  reg [7:0] v_12295 = 8'h0;
  wire [7:0] v_12296;
  wire [7:0] v_12297;
  function [7:0] mux_12297(input [0:0] sel);
    case (sel) 0: mux_12297 = 8'h0; 1: mux_12297 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12298;
  wire [7:0] v_12299;
  wire [7:0] v_12300;
  function [7:0] mux_12300(input [0:0] sel);
    case (sel) 0: mux_12300 = 8'h0; 1: mux_12300 = v_12301;
    endcase
  endfunction
  reg [7:0] v_12301 = 8'h0;
  wire [7:0] v_12302;
  wire [7:0] v_12303;
  function [7:0] mux_12303(input [0:0] sel);
    case (sel) 0: mux_12303 = 8'h0; 1: mux_12303 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12304;
  wire [7:0] v_12305;
  wire [7:0] v_12306;
  function [7:0] mux_12306(input [0:0] sel);
    case (sel) 0: mux_12306 = 8'h0; 1: mux_12306 = vout_peek_2517;
    endcase
  endfunction
  wire [7:0] v_12307;
  function [7:0] mux_12307(input [0:0] sel);
    case (sel) 0: mux_12307 = 8'h0; 1: mux_12307 = vout_peek_2509;
    endcase
  endfunction
  wire [7:0] v_12308;
  function [7:0] mux_12308(input [0:0] sel);
    case (sel) 0: mux_12308 = 8'h0; 1: mux_12308 = v_12309;
    endcase
  endfunction
  reg [7:0] v_12309 = 8'h0;
  wire [7:0] v_12310;
  wire [7:0] v_12311;
  function [7:0] mux_12311(input [0:0] sel);
    case (sel) 0: mux_12311 = 8'h0; 1: mux_12311 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12312;
  wire [7:0] v_12313;
  wire [7:0] v_12314;
  function [7:0] mux_12314(input [0:0] sel);
    case (sel) 0: mux_12314 = 8'h0; 1: mux_12314 = vout_peek_2503;
    endcase
  endfunction
  wire [7:0] v_12315;
  function [7:0] mux_12315(input [0:0] sel);
    case (sel) 0: mux_12315 = 8'h0; 1: mux_12315 = vout_peek_2495;
    endcase
  endfunction
  wire [7:0] v_12316;
  function [7:0] mux_12316(input [0:0] sel);
    case (sel) 0: mux_12316 = 8'h0; 1: mux_12316 = v_12317;
    endcase
  endfunction
  reg [7:0] v_12317 = 8'h0;
  wire [7:0] v_12318;
  wire [7:0] v_12319;
  function [7:0] mux_12319(input [0:0] sel);
    case (sel) 0: mux_12319 = 8'h0; 1: mux_12319 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12320;
  wire [7:0] v_12321;
  wire [7:0] v_12322;
  function [7:0] mux_12322(input [0:0] sel);
    case (sel) 0: mux_12322 = 8'h0; 1: mux_12322 = v_12323;
    endcase
  endfunction
  reg [7:0] v_12323 = 8'h0;
  wire [7:0] v_12324;
  wire [7:0] v_12325;
  function [7:0] mux_12325(input [0:0] sel);
    case (sel) 0: mux_12325 = 8'h0; 1: mux_12325 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12326;
  wire [7:0] v_12327;
  wire [7:0] v_12328;
  function [7:0] mux_12328(input [0:0] sel);
    case (sel) 0: mux_12328 = 8'h0; 1: mux_12328 = vout_peek_2489;
    endcase
  endfunction
  wire [7:0] v_12329;
  function [7:0] mux_12329(input [0:0] sel);
    case (sel) 0: mux_12329 = 8'h0; 1: mux_12329 = vout_peek_2481;
    endcase
  endfunction
  wire [7:0] v_12330;
  function [7:0] mux_12330(input [0:0] sel);
    case (sel) 0: mux_12330 = 8'h0; 1: mux_12330 = v_12331;
    endcase
  endfunction
  reg [7:0] v_12331 = 8'h0;
  wire [7:0] v_12332;
  wire [7:0] v_12333;
  function [7:0] mux_12333(input [0:0] sel);
    case (sel) 0: mux_12333 = 8'h0; 1: mux_12333 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12334;
  wire [7:0] v_12335;
  wire [7:0] v_12336;
  function [7:0] mux_12336(input [0:0] sel);
    case (sel) 0: mux_12336 = 8'h0; 1: mux_12336 = vout_peek_2475;
    endcase
  endfunction
  wire [7:0] v_12337;
  function [7:0] mux_12337(input [0:0] sel);
    case (sel) 0: mux_12337 = 8'h0; 1: mux_12337 = vout_peek_2467;
    endcase
  endfunction
  wire [7:0] v_12338;
  function [7:0] mux_12338(input [0:0] sel);
    case (sel) 0: mux_12338 = 8'h0; 1: mux_12338 = v_12339;
    endcase
  endfunction
  reg [7:0] v_12339 = 8'h0;
  wire [7:0] v_12340;
  wire [7:0] v_12341;
  function [7:0] mux_12341(input [0:0] sel);
    case (sel) 0: mux_12341 = 8'h0; 1: mux_12341 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12342;
  wire [7:0] v_12343;
  wire [7:0] v_12344;
  function [7:0] mux_12344(input [0:0] sel);
    case (sel) 0: mux_12344 = 8'h0; 1: mux_12344 = v_12345;
    endcase
  endfunction
  reg [7:0] v_12345 = 8'h0;
  wire [7:0] v_12346;
  wire [7:0] v_12347;
  function [7:0] mux_12347(input [0:0] sel);
    case (sel) 0: mux_12347 = 8'h0; 1: mux_12347 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12348;
  wire [7:0] v_12349;
  wire [7:0] v_12350;
  function [7:0] mux_12350(input [0:0] sel);
    case (sel) 0: mux_12350 = 8'h0; 1: mux_12350 = v_12351;
    endcase
  endfunction
  reg [7:0] v_12351 = 8'h0;
  wire [7:0] v_12352;
  wire [7:0] v_12353;
  function [7:0] mux_12353(input [0:0] sel);
    case (sel) 0: mux_12353 = 8'h0; 1: mux_12353 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12354;
  wire [7:0] v_12355;
  wire [7:0] v_12356;
  function [7:0] mux_12356(input [0:0] sel);
    case (sel) 0: mux_12356 = 8'h0; 1: mux_12356 = v_12357;
    endcase
  endfunction
  reg [7:0] v_12357 = 8'h0;
  wire [7:0] v_12358;
  wire [7:0] v_12359;
  function [7:0] mux_12359(input [0:0] sel);
    case (sel) 0: mux_12359 = 8'h0; 1: mux_12359 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12360;
  wire [7:0] v_12361;
  wire [7:0] v_12362;
  function [7:0] mux_12362(input [0:0] sel);
    case (sel) 0: mux_12362 = 8'h0; 1: mux_12362 = v_12363;
    endcase
  endfunction
  reg [7:0] v_12363 = 8'h0;
  wire [7:0] v_12364;
  wire [7:0] v_12365;
  function [7:0] mux_12365(input [0:0] sel);
    case (sel) 0: mux_12365 = 8'h0; 1: mux_12365 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12366;
  wire [7:0] v_12367;
  wire [7:0] v_12368;
  function [7:0] mux_12368(input [0:0] sel);
    case (sel) 0: mux_12368 = 8'h0; 1: mux_12368 = v_12369;
    endcase
  endfunction
  reg [7:0] v_12369 = 8'h0;
  wire [7:0] v_12370;
  wire [7:0] v_12371;
  function [7:0] mux_12371(input [0:0] sel);
    case (sel) 0: mux_12371 = 8'h0; 1: mux_12371 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12372;
  wire [7:0] v_12373;
  wire [7:0] v_12374;
  function [7:0] mux_12374(input [0:0] sel);
    case (sel) 0: mux_12374 = 8'h0; 1: mux_12374 = vout_peek_2461;
    endcase
  endfunction
  wire [7:0] v_12375;
  function [7:0] mux_12375(input [0:0] sel);
    case (sel) 0: mux_12375 = 8'h0; 1: mux_12375 = vout_peek_2453;
    endcase
  endfunction
  wire [7:0] v_12376;
  function [7:0] mux_12376(input [0:0] sel);
    case (sel) 0: mux_12376 = 8'h0; 1: mux_12376 = v_12377;
    endcase
  endfunction
  reg [7:0] v_12377 = 8'h0;
  wire [7:0] v_12378;
  wire [7:0] v_12379;
  function [7:0] mux_12379(input [0:0] sel);
    case (sel) 0: mux_12379 = 8'h0; 1: mux_12379 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12380;
  wire [7:0] v_12381;
  wire [7:0] v_12382;
  function [7:0] mux_12382(input [0:0] sel);
    case (sel) 0: mux_12382 = 8'h0; 1: mux_12382 = vout_peek_2447;
    endcase
  endfunction
  wire [7:0] v_12383;
  function [7:0] mux_12383(input [0:0] sel);
    case (sel) 0: mux_12383 = 8'h0; 1: mux_12383 = vout_peek_2439;
    endcase
  endfunction
  wire [7:0] v_12384;
  function [7:0] mux_12384(input [0:0] sel);
    case (sel) 0: mux_12384 = 8'h0; 1: mux_12384 = v_12385;
    endcase
  endfunction
  reg [7:0] v_12385 = 8'h0;
  wire [7:0] v_12386;
  wire [7:0] v_12387;
  function [7:0] mux_12387(input [0:0] sel);
    case (sel) 0: mux_12387 = 8'h0; 1: mux_12387 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12388;
  wire [7:0] v_12389;
  wire [7:0] v_12390;
  function [7:0] mux_12390(input [0:0] sel);
    case (sel) 0: mux_12390 = 8'h0; 1: mux_12390 = v_12391;
    endcase
  endfunction
  reg [7:0] v_12391 = 8'h0;
  wire [7:0] v_12392;
  wire [7:0] v_12393;
  function [7:0] mux_12393(input [0:0] sel);
    case (sel) 0: mux_12393 = 8'h0; 1: mux_12393 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12394;
  wire [7:0] v_12395;
  wire [7:0] v_12396;
  function [7:0] mux_12396(input [0:0] sel);
    case (sel) 0: mux_12396 = 8'h0; 1: mux_12396 = vout_peek_2433;
    endcase
  endfunction
  wire [7:0] v_12397;
  function [7:0] mux_12397(input [0:0] sel);
    case (sel) 0: mux_12397 = 8'h0; 1: mux_12397 = vout_peek_2425;
    endcase
  endfunction
  wire [7:0] v_12398;
  function [7:0] mux_12398(input [0:0] sel);
    case (sel) 0: mux_12398 = 8'h0; 1: mux_12398 = v_12399;
    endcase
  endfunction
  reg [7:0] v_12399 = 8'h0;
  wire [7:0] v_12400;
  wire [7:0] v_12401;
  function [7:0] mux_12401(input [0:0] sel);
    case (sel) 0: mux_12401 = 8'h0; 1: mux_12401 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12402;
  wire [7:0] v_12403;
  wire [7:0] v_12404;
  function [7:0] mux_12404(input [0:0] sel);
    case (sel) 0: mux_12404 = 8'h0; 1: mux_12404 = vout_peek_2419;
    endcase
  endfunction
  wire [7:0] v_12405;
  function [7:0] mux_12405(input [0:0] sel);
    case (sel) 0: mux_12405 = 8'h0; 1: mux_12405 = vout_peek_2411;
    endcase
  endfunction
  wire [7:0] v_12406;
  function [7:0] mux_12406(input [0:0] sel);
    case (sel) 0: mux_12406 = 8'h0; 1: mux_12406 = v_12407;
    endcase
  endfunction
  reg [7:0] v_12407 = 8'h0;
  wire [7:0] v_12408;
  wire [7:0] v_12409;
  function [7:0] mux_12409(input [0:0] sel);
    case (sel) 0: mux_12409 = 8'h0; 1: mux_12409 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12410;
  wire [7:0] v_12411;
  wire [7:0] v_12412;
  function [7:0] mux_12412(input [0:0] sel);
    case (sel) 0: mux_12412 = 8'h0; 1: mux_12412 = v_12413;
    endcase
  endfunction
  reg [7:0] v_12413 = 8'h0;
  wire [7:0] v_12414;
  wire [7:0] v_12415;
  function [7:0] mux_12415(input [0:0] sel);
    case (sel) 0: mux_12415 = 8'h0; 1: mux_12415 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12416;
  wire [7:0] v_12417;
  wire [7:0] v_12418;
  function [7:0] mux_12418(input [0:0] sel);
    case (sel) 0: mux_12418 = 8'h0; 1: mux_12418 = v_12419;
    endcase
  endfunction
  reg [7:0] v_12419 = 8'h0;
  wire [7:0] v_12420;
  wire [7:0] v_12421;
  function [7:0] mux_12421(input [0:0] sel);
    case (sel) 0: mux_12421 = 8'h0; 1: mux_12421 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12422;
  wire [7:0] v_12423;
  wire [7:0] v_12424;
  function [7:0] mux_12424(input [0:0] sel);
    case (sel) 0: mux_12424 = 8'h0; 1: mux_12424 = vout_peek_2405;
    endcase
  endfunction
  wire [7:0] v_12425;
  function [7:0] mux_12425(input [0:0] sel);
    case (sel) 0: mux_12425 = 8'h0; 1: mux_12425 = vout_peek_2397;
    endcase
  endfunction
  wire [7:0] v_12426;
  function [7:0] mux_12426(input [0:0] sel);
    case (sel) 0: mux_12426 = 8'h0; 1: mux_12426 = v_12427;
    endcase
  endfunction
  reg [7:0] v_12427 = 8'h0;
  wire [7:0] v_12428;
  wire [7:0] v_12429;
  function [7:0] mux_12429(input [0:0] sel);
    case (sel) 0: mux_12429 = 8'h0; 1: mux_12429 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12430;
  wire [7:0] v_12431;
  wire [7:0] v_12432;
  function [7:0] mux_12432(input [0:0] sel);
    case (sel) 0: mux_12432 = 8'h0; 1: mux_12432 = vout_peek_2391;
    endcase
  endfunction
  wire [7:0] v_12433;
  function [7:0] mux_12433(input [0:0] sel);
    case (sel) 0: mux_12433 = 8'h0; 1: mux_12433 = vout_peek_2383;
    endcase
  endfunction
  wire [7:0] v_12434;
  function [7:0] mux_12434(input [0:0] sel);
    case (sel) 0: mux_12434 = 8'h0; 1: mux_12434 = v_12435;
    endcase
  endfunction
  reg [7:0] v_12435 = 8'h0;
  wire [7:0] v_12436;
  wire [7:0] v_12437;
  function [7:0] mux_12437(input [0:0] sel);
    case (sel) 0: mux_12437 = 8'h0; 1: mux_12437 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12438;
  wire [7:0] v_12439;
  wire [7:0] v_12440;
  function [7:0] mux_12440(input [0:0] sel);
    case (sel) 0: mux_12440 = 8'h0; 1: mux_12440 = v_12441;
    endcase
  endfunction
  reg [7:0] v_12441 = 8'h0;
  wire [7:0] v_12442;
  wire [7:0] v_12443;
  function [7:0] mux_12443(input [0:0] sel);
    case (sel) 0: mux_12443 = 8'h0; 1: mux_12443 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12444;
  wire [7:0] v_12445;
  wire [7:0] v_12446;
  function [7:0] mux_12446(input [0:0] sel);
    case (sel) 0: mux_12446 = 8'h0; 1: mux_12446 = vout_peek_2377;
    endcase
  endfunction
  wire [7:0] v_12447;
  function [7:0] mux_12447(input [0:0] sel);
    case (sel) 0: mux_12447 = 8'h0; 1: mux_12447 = vout_peek_2369;
    endcase
  endfunction
  wire [7:0] v_12448;
  function [7:0] mux_12448(input [0:0] sel);
    case (sel) 0: mux_12448 = 8'h0; 1: mux_12448 = v_12449;
    endcase
  endfunction
  reg [7:0] v_12449 = 8'h0;
  wire [7:0] v_12450;
  wire [7:0] v_12451;
  function [7:0] mux_12451(input [0:0] sel);
    case (sel) 0: mux_12451 = 8'h0; 1: mux_12451 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12452;
  wire [7:0] v_12453;
  wire [7:0] v_12454;
  function [7:0] mux_12454(input [0:0] sel);
    case (sel) 0: mux_12454 = 8'h0; 1: mux_12454 = vout_peek_2363;
    endcase
  endfunction
  wire [7:0] v_12455;
  function [7:0] mux_12455(input [0:0] sel);
    case (sel) 0: mux_12455 = 8'h0; 1: mux_12455 = vout_peek_2355;
    endcase
  endfunction
  wire [7:0] v_12456;
  function [7:0] mux_12456(input [0:0] sel);
    case (sel) 0: mux_12456 = 8'h0; 1: mux_12456 = v_12457;
    endcase
  endfunction
  reg [7:0] v_12457 = 8'h0;
  wire [7:0] v_12458;
  wire [7:0] v_12459;
  function [7:0] mux_12459(input [0:0] sel);
    case (sel) 0: mux_12459 = 8'h0; 1: mux_12459 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12460;
  wire [7:0] v_12461;
  wire [7:0] v_12462;
  function [7:0] mux_12462(input [0:0] sel);
    case (sel) 0: mux_12462 = 8'h0; 1: mux_12462 = v_12463;
    endcase
  endfunction
  reg [7:0] v_12463 = 8'h0;
  wire [7:0] v_12464;
  wire [7:0] v_12465;
  function [7:0] mux_12465(input [0:0] sel);
    case (sel) 0: mux_12465 = 8'h0; 1: mux_12465 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12466;
  wire [7:0] v_12467;
  wire [7:0] v_12468;
  function [7:0] mux_12468(input [0:0] sel);
    case (sel) 0: mux_12468 = 8'h0; 1: mux_12468 = v_12469;
    endcase
  endfunction
  reg [7:0] v_12469 = 8'h0;
  wire [7:0] v_12470;
  wire [7:0] v_12471;
  function [7:0] mux_12471(input [0:0] sel);
    case (sel) 0: mux_12471 = 8'h0; 1: mux_12471 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12472;
  wire [7:0] v_12473;
  wire [7:0] v_12474;
  function [7:0] mux_12474(input [0:0] sel);
    case (sel) 0: mux_12474 = 8'h0; 1: mux_12474 = v_12475;
    endcase
  endfunction
  reg [7:0] v_12475 = 8'h0;
  wire [7:0] v_12476;
  wire [7:0] v_12477;
  function [7:0] mux_12477(input [0:0] sel);
    case (sel) 0: mux_12477 = 8'h0; 1: mux_12477 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12478;
  wire [7:0] v_12479;
  wire [7:0] v_12480;
  function [7:0] mux_12480(input [0:0] sel);
    case (sel) 0: mux_12480 = 8'h0; 1: mux_12480 = vout_peek_2349;
    endcase
  endfunction
  wire [7:0] v_12481;
  function [7:0] mux_12481(input [0:0] sel);
    case (sel) 0: mux_12481 = 8'h0; 1: mux_12481 = vout_peek_2341;
    endcase
  endfunction
  wire [7:0] v_12482;
  function [7:0] mux_12482(input [0:0] sel);
    case (sel) 0: mux_12482 = 8'h0; 1: mux_12482 = v_12483;
    endcase
  endfunction
  reg [7:0] v_12483 = 8'h0;
  wire [7:0] v_12484;
  wire [7:0] v_12485;
  function [7:0] mux_12485(input [0:0] sel);
    case (sel) 0: mux_12485 = 8'h0; 1: mux_12485 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12486;
  wire [7:0] v_12487;
  wire [7:0] v_12488;
  function [7:0] mux_12488(input [0:0] sel);
    case (sel) 0: mux_12488 = 8'h0; 1: mux_12488 = vout_peek_2335;
    endcase
  endfunction
  wire [7:0] v_12489;
  function [7:0] mux_12489(input [0:0] sel);
    case (sel) 0: mux_12489 = 8'h0; 1: mux_12489 = vout_peek_2327;
    endcase
  endfunction
  wire [7:0] v_12490;
  function [7:0] mux_12490(input [0:0] sel);
    case (sel) 0: mux_12490 = 8'h0; 1: mux_12490 = v_12491;
    endcase
  endfunction
  reg [7:0] v_12491 = 8'h0;
  wire [7:0] v_12492;
  wire [7:0] v_12493;
  function [7:0] mux_12493(input [0:0] sel);
    case (sel) 0: mux_12493 = 8'h0; 1: mux_12493 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12494;
  wire [7:0] v_12495;
  wire [7:0] v_12496;
  function [7:0] mux_12496(input [0:0] sel);
    case (sel) 0: mux_12496 = 8'h0; 1: mux_12496 = v_12497;
    endcase
  endfunction
  reg [7:0] v_12497 = 8'h0;
  wire [7:0] v_12498;
  wire [7:0] v_12499;
  function [7:0] mux_12499(input [0:0] sel);
    case (sel) 0: mux_12499 = 8'h0; 1: mux_12499 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12500;
  wire [7:0] v_12501;
  wire [7:0] v_12502;
  function [7:0] mux_12502(input [0:0] sel);
    case (sel) 0: mux_12502 = 8'h0; 1: mux_12502 = vout_peek_2321;
    endcase
  endfunction
  wire [7:0] v_12503;
  function [7:0] mux_12503(input [0:0] sel);
    case (sel) 0: mux_12503 = 8'h0; 1: mux_12503 = vout_peek_2313;
    endcase
  endfunction
  wire [7:0] v_12504;
  function [7:0] mux_12504(input [0:0] sel);
    case (sel) 0: mux_12504 = 8'h0; 1: mux_12504 = v_12505;
    endcase
  endfunction
  reg [7:0] v_12505 = 8'h0;
  wire [7:0] v_12506;
  wire [7:0] v_12507;
  function [7:0] mux_12507(input [0:0] sel);
    case (sel) 0: mux_12507 = 8'h0; 1: mux_12507 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12508;
  wire [7:0] v_12509;
  wire [7:0] v_12510;
  function [7:0] mux_12510(input [0:0] sel);
    case (sel) 0: mux_12510 = 8'h0; 1: mux_12510 = vout_peek_2307;
    endcase
  endfunction
  wire [7:0] v_12511;
  function [7:0] mux_12511(input [0:0] sel);
    case (sel) 0: mux_12511 = 8'h0; 1: mux_12511 = vout_peek_2299;
    endcase
  endfunction
  wire [7:0] v_12512;
  function [7:0] mux_12512(input [0:0] sel);
    case (sel) 0: mux_12512 = 8'h0; 1: mux_12512 = v_12513;
    endcase
  endfunction
  reg [7:0] v_12513 = 8'h0;
  wire [7:0] v_12514;
  wire [7:0] v_12515;
  function [7:0] mux_12515(input [0:0] sel);
    case (sel) 0: mux_12515 = 8'h0; 1: mux_12515 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12516;
  wire [7:0] v_12517;
  wire [7:0] v_12518;
  function [7:0] mux_12518(input [0:0] sel);
    case (sel) 0: mux_12518 = 8'h0; 1: mux_12518 = v_12519;
    endcase
  endfunction
  reg [7:0] v_12519 = 8'h0;
  wire [7:0] v_12520;
  wire [7:0] v_12521;
  function [7:0] mux_12521(input [0:0] sel);
    case (sel) 0: mux_12521 = 8'h0; 1: mux_12521 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12522;
  wire [7:0] v_12523;
  wire [7:0] v_12524;
  function [7:0] mux_12524(input [0:0] sel);
    case (sel) 0: mux_12524 = 8'h0; 1: mux_12524 = v_12525;
    endcase
  endfunction
  reg [7:0] v_12525 = 8'h0;
  wire [7:0] v_12526;
  wire [7:0] v_12527;
  function [7:0] mux_12527(input [0:0] sel);
    case (sel) 0: mux_12527 = 8'h0; 1: mux_12527 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12528;
  wire [7:0] v_12529;
  wire [7:0] v_12530;
  function [7:0] mux_12530(input [0:0] sel);
    case (sel) 0: mux_12530 = 8'h0; 1: mux_12530 = vout_peek_2293;
    endcase
  endfunction
  wire [7:0] v_12531;
  function [7:0] mux_12531(input [0:0] sel);
    case (sel) 0: mux_12531 = 8'h0; 1: mux_12531 = vout_peek_2285;
    endcase
  endfunction
  wire [7:0] v_12532;
  function [7:0] mux_12532(input [0:0] sel);
    case (sel) 0: mux_12532 = 8'h0; 1: mux_12532 = v_12533;
    endcase
  endfunction
  reg [7:0] v_12533 = 8'h0;
  wire [7:0] v_12534;
  wire [7:0] v_12535;
  function [7:0] mux_12535(input [0:0] sel);
    case (sel) 0: mux_12535 = 8'h0; 1: mux_12535 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12536;
  wire [7:0] v_12537;
  wire [7:0] v_12538;
  function [7:0] mux_12538(input [0:0] sel);
    case (sel) 0: mux_12538 = 8'h0; 1: mux_12538 = vout_peek_2279;
    endcase
  endfunction
  wire [7:0] v_12539;
  function [7:0] mux_12539(input [0:0] sel);
    case (sel) 0: mux_12539 = 8'h0; 1: mux_12539 = vout_peek_2271;
    endcase
  endfunction
  wire [7:0] v_12540;
  function [7:0] mux_12540(input [0:0] sel);
    case (sel) 0: mux_12540 = 8'h0; 1: mux_12540 = v_12541;
    endcase
  endfunction
  reg [7:0] v_12541 = 8'h0;
  wire [7:0] v_12542;
  wire [7:0] v_12543;
  function [7:0] mux_12543(input [0:0] sel);
    case (sel) 0: mux_12543 = 8'h0; 1: mux_12543 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12544;
  wire [7:0] v_12545;
  wire [7:0] v_12546;
  function [7:0] mux_12546(input [0:0] sel);
    case (sel) 0: mux_12546 = 8'h0; 1: mux_12546 = v_12547;
    endcase
  endfunction
  reg [7:0] v_12547 = 8'h0;
  wire [7:0] v_12548;
  wire [7:0] v_12549;
  function [7:0] mux_12549(input [0:0] sel);
    case (sel) 0: mux_12549 = 8'h0; 1: mux_12549 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12550;
  wire [7:0] v_12551;
  wire [7:0] v_12552;
  function [7:0] mux_12552(input [0:0] sel);
    case (sel) 0: mux_12552 = 8'h0; 1: mux_12552 = vout_peek_2265;
    endcase
  endfunction
  wire [7:0] v_12553;
  function [7:0] mux_12553(input [0:0] sel);
    case (sel) 0: mux_12553 = 8'h0; 1: mux_12553 = vout_peek_2257;
    endcase
  endfunction
  wire [7:0] v_12554;
  function [7:0] mux_12554(input [0:0] sel);
    case (sel) 0: mux_12554 = 8'h0; 1: mux_12554 = v_12555;
    endcase
  endfunction
  reg [7:0] v_12555 = 8'h0;
  wire [7:0] v_12556;
  wire [7:0] v_12557;
  function [7:0] mux_12557(input [0:0] sel);
    case (sel) 0: mux_12557 = 8'h0; 1: mux_12557 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12558;
  wire [7:0] v_12559;
  wire [7:0] v_12560;
  function [7:0] mux_12560(input [0:0] sel);
    case (sel) 0: mux_12560 = 8'h0; 1: mux_12560 = vout_peek_2251;
    endcase
  endfunction
  wire [7:0] v_12561;
  function [7:0] mux_12561(input [0:0] sel);
    case (sel) 0: mux_12561 = 8'h0; 1: mux_12561 = vout_peek_2243;
    endcase
  endfunction
  wire [7:0] v_12562;
  function [7:0] mux_12562(input [0:0] sel);
    case (sel) 0: mux_12562 = 8'h0; 1: mux_12562 = v_12563;
    endcase
  endfunction
  reg [7:0] v_12563 = 8'h0;
  wire [7:0] v_12564;
  wire [7:0] v_12565;
  function [7:0] mux_12565(input [0:0] sel);
    case (sel) 0: mux_12565 = 8'h0; 1: mux_12565 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12566;
  wire [7:0] v_12567;
  wire [7:0] v_12568;
  function [7:0] mux_12568(input [0:0] sel);
    case (sel) 0: mux_12568 = 8'h0; 1: mux_12568 = v_12569;
    endcase
  endfunction
  reg [7:0] v_12569 = 8'h0;
  wire [7:0] v_12570;
  wire [7:0] v_12571;
  function [7:0] mux_12571(input [0:0] sel);
    case (sel) 0: mux_12571 = 8'h0; 1: mux_12571 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12572;
  wire [7:0] v_12573;
  wire [7:0] v_12574;
  function [7:0] mux_12574(input [0:0] sel);
    case (sel) 0: mux_12574 = 8'h0; 1: mux_12574 = v_12575;
    endcase
  endfunction
  reg [7:0] v_12575 = 8'h0;
  wire [7:0] v_12576;
  wire [7:0] v_12577;
  function [7:0] mux_12577(input [0:0] sel);
    case (sel) 0: mux_12577 = 8'h0; 1: mux_12577 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12578;
  wire [7:0] v_12579;
  wire [7:0] v_12580;
  function [7:0] mux_12580(input [0:0] sel);
    case (sel) 0: mux_12580 = 8'h0; 1: mux_12580 = v_12581;
    endcase
  endfunction
  reg [7:0] v_12581 = 8'h0;
  wire [7:0] v_12582;
  wire [7:0] v_12583;
  function [7:0] mux_12583(input [0:0] sel);
    case (sel) 0: mux_12583 = 8'h0; 1: mux_12583 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12584;
  wire [7:0] v_12585;
  wire [7:0] v_12586;
  function [7:0] mux_12586(input [0:0] sel);
    case (sel) 0: mux_12586 = 8'h0; 1: mux_12586 = v_12587;
    endcase
  endfunction
  reg [7:0] v_12587 = 8'h0;
  wire [7:0] v_12588;
  wire [7:0] v_12589;
  function [7:0] mux_12589(input [0:0] sel);
    case (sel) 0: mux_12589 = 8'h0; 1: mux_12589 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12590;
  wire [7:0] v_12591;
  wire [7:0] v_12592;
  function [7:0] mux_12592(input [0:0] sel);
    case (sel) 0: mux_12592 = 8'h0; 1: mux_12592 = vout_peek_2237;
    endcase
  endfunction
  wire [7:0] v_12593;
  function [7:0] mux_12593(input [0:0] sel);
    case (sel) 0: mux_12593 = 8'h0; 1: mux_12593 = vout_peek_2229;
    endcase
  endfunction
  wire [7:0] v_12594;
  function [7:0] mux_12594(input [0:0] sel);
    case (sel) 0: mux_12594 = 8'h0; 1: mux_12594 = v_12595;
    endcase
  endfunction
  reg [7:0] v_12595 = 8'h0;
  wire [7:0] v_12596;
  wire [7:0] v_12597;
  function [7:0] mux_12597(input [0:0] sel);
    case (sel) 0: mux_12597 = 8'h0; 1: mux_12597 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12598;
  wire [7:0] v_12599;
  wire [7:0] v_12600;
  function [7:0] mux_12600(input [0:0] sel);
    case (sel) 0: mux_12600 = 8'h0; 1: mux_12600 = vout_peek_2223;
    endcase
  endfunction
  wire [7:0] v_12601;
  function [7:0] mux_12601(input [0:0] sel);
    case (sel) 0: mux_12601 = 8'h0; 1: mux_12601 = vout_peek_2215;
    endcase
  endfunction
  wire [7:0] v_12602;
  function [7:0] mux_12602(input [0:0] sel);
    case (sel) 0: mux_12602 = 8'h0; 1: mux_12602 = v_12603;
    endcase
  endfunction
  reg [7:0] v_12603 = 8'h0;
  wire [7:0] v_12604;
  wire [7:0] v_12605;
  function [7:0] mux_12605(input [0:0] sel);
    case (sel) 0: mux_12605 = 8'h0; 1: mux_12605 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12606;
  wire [7:0] v_12607;
  wire [7:0] v_12608;
  function [7:0] mux_12608(input [0:0] sel);
    case (sel) 0: mux_12608 = 8'h0; 1: mux_12608 = v_12609;
    endcase
  endfunction
  reg [7:0] v_12609 = 8'h0;
  wire [7:0] v_12610;
  wire [7:0] v_12611;
  function [7:0] mux_12611(input [0:0] sel);
    case (sel) 0: mux_12611 = 8'h0; 1: mux_12611 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12612;
  wire [7:0] v_12613;
  wire [7:0] v_12614;
  function [7:0] mux_12614(input [0:0] sel);
    case (sel) 0: mux_12614 = 8'h0; 1: mux_12614 = vout_peek_2209;
    endcase
  endfunction
  wire [7:0] v_12615;
  function [7:0] mux_12615(input [0:0] sel);
    case (sel) 0: mux_12615 = 8'h0; 1: mux_12615 = vout_peek_2201;
    endcase
  endfunction
  wire [7:0] v_12616;
  function [7:0] mux_12616(input [0:0] sel);
    case (sel) 0: mux_12616 = 8'h0; 1: mux_12616 = v_12617;
    endcase
  endfunction
  reg [7:0] v_12617 = 8'h0;
  wire [7:0] v_12618;
  wire [7:0] v_12619;
  function [7:0] mux_12619(input [0:0] sel);
    case (sel) 0: mux_12619 = 8'h0; 1: mux_12619 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12620;
  wire [7:0] v_12621;
  wire [7:0] v_12622;
  function [7:0] mux_12622(input [0:0] sel);
    case (sel) 0: mux_12622 = 8'h0; 1: mux_12622 = vout_peek_2195;
    endcase
  endfunction
  wire [7:0] v_12623;
  function [7:0] mux_12623(input [0:0] sel);
    case (sel) 0: mux_12623 = 8'h0; 1: mux_12623 = vout_peek_2187;
    endcase
  endfunction
  wire [7:0] v_12624;
  function [7:0] mux_12624(input [0:0] sel);
    case (sel) 0: mux_12624 = 8'h0; 1: mux_12624 = v_12625;
    endcase
  endfunction
  reg [7:0] v_12625 = 8'h0;
  wire [7:0] v_12626;
  wire [7:0] v_12627;
  function [7:0] mux_12627(input [0:0] sel);
    case (sel) 0: mux_12627 = 8'h0; 1: mux_12627 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12628;
  wire [7:0] v_12629;
  wire [7:0] v_12630;
  function [7:0] mux_12630(input [0:0] sel);
    case (sel) 0: mux_12630 = 8'h0; 1: mux_12630 = v_12631;
    endcase
  endfunction
  reg [7:0] v_12631 = 8'h0;
  wire [7:0] v_12632;
  wire [7:0] v_12633;
  function [7:0] mux_12633(input [0:0] sel);
    case (sel) 0: mux_12633 = 8'h0; 1: mux_12633 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12634;
  wire [7:0] v_12635;
  wire [7:0] v_12636;
  function [7:0] mux_12636(input [0:0] sel);
    case (sel) 0: mux_12636 = 8'h0; 1: mux_12636 = v_12637;
    endcase
  endfunction
  reg [7:0] v_12637 = 8'h0;
  wire [7:0] v_12638;
  wire [7:0] v_12639;
  function [7:0] mux_12639(input [0:0] sel);
    case (sel) 0: mux_12639 = 8'h0; 1: mux_12639 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12640;
  wire [7:0] v_12641;
  wire [7:0] v_12642;
  function [7:0] mux_12642(input [0:0] sel);
    case (sel) 0: mux_12642 = 8'h0; 1: mux_12642 = vout_peek_2181;
    endcase
  endfunction
  wire [7:0] v_12643;
  function [7:0] mux_12643(input [0:0] sel);
    case (sel) 0: mux_12643 = 8'h0; 1: mux_12643 = vout_peek_2173;
    endcase
  endfunction
  wire [7:0] v_12644;
  function [7:0] mux_12644(input [0:0] sel);
    case (sel) 0: mux_12644 = 8'h0; 1: mux_12644 = v_12645;
    endcase
  endfunction
  reg [7:0] v_12645 = 8'h0;
  wire [7:0] v_12646;
  wire [7:0] v_12647;
  function [7:0] mux_12647(input [0:0] sel);
    case (sel) 0: mux_12647 = 8'h0; 1: mux_12647 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12648;
  wire [7:0] v_12649;
  wire [7:0] v_12650;
  function [7:0] mux_12650(input [0:0] sel);
    case (sel) 0: mux_12650 = 8'h0; 1: mux_12650 = vout_peek_2167;
    endcase
  endfunction
  wire [7:0] v_12651;
  function [7:0] mux_12651(input [0:0] sel);
    case (sel) 0: mux_12651 = 8'h0; 1: mux_12651 = vout_peek_2159;
    endcase
  endfunction
  wire [7:0] v_12652;
  function [7:0] mux_12652(input [0:0] sel);
    case (sel) 0: mux_12652 = 8'h0; 1: mux_12652 = v_12653;
    endcase
  endfunction
  reg [7:0] v_12653 = 8'h0;
  wire [7:0] v_12654;
  wire [7:0] v_12655;
  function [7:0] mux_12655(input [0:0] sel);
    case (sel) 0: mux_12655 = 8'h0; 1: mux_12655 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12656;
  wire [7:0] v_12657;
  wire [7:0] v_12658;
  function [7:0] mux_12658(input [0:0] sel);
    case (sel) 0: mux_12658 = 8'h0; 1: mux_12658 = v_12659;
    endcase
  endfunction
  reg [7:0] v_12659 = 8'h0;
  wire [7:0] v_12660;
  wire [7:0] v_12661;
  function [7:0] mux_12661(input [0:0] sel);
    case (sel) 0: mux_12661 = 8'h0; 1: mux_12661 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12662;
  wire [7:0] v_12663;
  wire [7:0] v_12664;
  function [7:0] mux_12664(input [0:0] sel);
    case (sel) 0: mux_12664 = 8'h0; 1: mux_12664 = vout_peek_2153;
    endcase
  endfunction
  wire [7:0] v_12665;
  function [7:0] mux_12665(input [0:0] sel);
    case (sel) 0: mux_12665 = 8'h0; 1: mux_12665 = vout_peek_2145;
    endcase
  endfunction
  wire [7:0] v_12666;
  function [7:0] mux_12666(input [0:0] sel);
    case (sel) 0: mux_12666 = 8'h0; 1: mux_12666 = v_12667;
    endcase
  endfunction
  reg [7:0] v_12667 = 8'h0;
  wire [7:0] v_12668;
  wire [7:0] v_12669;
  function [7:0] mux_12669(input [0:0] sel);
    case (sel) 0: mux_12669 = 8'h0; 1: mux_12669 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12670;
  wire [7:0] v_12671;
  wire [7:0] v_12672;
  function [7:0] mux_12672(input [0:0] sel);
    case (sel) 0: mux_12672 = 8'h0; 1: mux_12672 = vout_peek_2139;
    endcase
  endfunction
  wire [7:0] v_12673;
  function [7:0] mux_12673(input [0:0] sel);
    case (sel) 0: mux_12673 = 8'h0; 1: mux_12673 = vout_peek_2131;
    endcase
  endfunction
  wire [7:0] v_12674;
  function [7:0] mux_12674(input [0:0] sel);
    case (sel) 0: mux_12674 = 8'h0; 1: mux_12674 = v_12675;
    endcase
  endfunction
  reg [7:0] v_12675 = 8'h0;
  wire [7:0] v_12676;
  wire [7:0] v_12677;
  function [7:0] mux_12677(input [0:0] sel);
    case (sel) 0: mux_12677 = 8'h0; 1: mux_12677 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12678;
  wire [7:0] v_12679;
  wire [7:0] v_12680;
  function [7:0] mux_12680(input [0:0] sel);
    case (sel) 0: mux_12680 = 8'h0; 1: mux_12680 = v_12681;
    endcase
  endfunction
  reg [7:0] v_12681 = 8'h0;
  wire [7:0] v_12682;
  wire [7:0] v_12683;
  function [7:0] mux_12683(input [0:0] sel);
    case (sel) 0: mux_12683 = 8'h0; 1: mux_12683 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12684;
  wire [7:0] v_12685;
  wire [7:0] v_12686;
  function [7:0] mux_12686(input [0:0] sel);
    case (sel) 0: mux_12686 = 8'h0; 1: mux_12686 = v_12687;
    endcase
  endfunction
  reg [7:0] v_12687 = 8'h0;
  wire [7:0] v_12688;
  wire [7:0] v_12689;
  function [7:0] mux_12689(input [0:0] sel);
    case (sel) 0: mux_12689 = 8'h0; 1: mux_12689 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12690;
  wire [7:0] v_12691;
  wire [7:0] v_12692;
  function [7:0] mux_12692(input [0:0] sel);
    case (sel) 0: mux_12692 = 8'h0; 1: mux_12692 = v_12693;
    endcase
  endfunction
  reg [7:0] v_12693 = 8'h0;
  wire [7:0] v_12694;
  wire [7:0] v_12695;
  function [7:0] mux_12695(input [0:0] sel);
    case (sel) 0: mux_12695 = 8'h0; 1: mux_12695 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12696;
  wire [7:0] v_12697;
  wire [7:0] v_12698;
  function [7:0] mux_12698(input [0:0] sel);
    case (sel) 0: mux_12698 = 8'h0; 1: mux_12698 = vout_peek_2125;
    endcase
  endfunction
  wire [7:0] v_12699;
  function [7:0] mux_12699(input [0:0] sel);
    case (sel) 0: mux_12699 = 8'h0; 1: mux_12699 = vout_peek_2117;
    endcase
  endfunction
  wire [7:0] v_12700;
  function [7:0] mux_12700(input [0:0] sel);
    case (sel) 0: mux_12700 = 8'h0; 1: mux_12700 = v_12701;
    endcase
  endfunction
  reg [7:0] v_12701 = 8'h0;
  wire [7:0] v_12702;
  wire [7:0] v_12703;
  function [7:0] mux_12703(input [0:0] sel);
    case (sel) 0: mux_12703 = 8'h0; 1: mux_12703 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12704;
  wire [7:0] v_12705;
  wire [7:0] v_12706;
  function [7:0] mux_12706(input [0:0] sel);
    case (sel) 0: mux_12706 = 8'h0; 1: mux_12706 = vout_peek_2111;
    endcase
  endfunction
  wire [7:0] v_12707;
  function [7:0] mux_12707(input [0:0] sel);
    case (sel) 0: mux_12707 = 8'h0; 1: mux_12707 = vout_peek_2103;
    endcase
  endfunction
  wire [7:0] v_12708;
  function [7:0] mux_12708(input [0:0] sel);
    case (sel) 0: mux_12708 = 8'h0; 1: mux_12708 = v_12709;
    endcase
  endfunction
  reg [7:0] v_12709 = 8'h0;
  wire [7:0] v_12710;
  wire [7:0] v_12711;
  function [7:0] mux_12711(input [0:0] sel);
    case (sel) 0: mux_12711 = 8'h0; 1: mux_12711 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12712;
  wire [7:0] v_12713;
  wire [7:0] v_12714;
  function [7:0] mux_12714(input [0:0] sel);
    case (sel) 0: mux_12714 = 8'h0; 1: mux_12714 = v_12715;
    endcase
  endfunction
  reg [7:0] v_12715 = 8'h0;
  wire [7:0] v_12716;
  wire [7:0] v_12717;
  function [7:0] mux_12717(input [0:0] sel);
    case (sel) 0: mux_12717 = 8'h0; 1: mux_12717 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12718;
  wire [7:0] v_12719;
  wire [7:0] v_12720;
  function [7:0] mux_12720(input [0:0] sel);
    case (sel) 0: mux_12720 = 8'h0; 1: mux_12720 = vout_peek_2097;
    endcase
  endfunction
  wire [7:0] v_12721;
  function [7:0] mux_12721(input [0:0] sel);
    case (sel) 0: mux_12721 = 8'h0; 1: mux_12721 = vout_peek_2089;
    endcase
  endfunction
  wire [7:0] v_12722;
  function [7:0] mux_12722(input [0:0] sel);
    case (sel) 0: mux_12722 = 8'h0; 1: mux_12722 = v_12723;
    endcase
  endfunction
  reg [7:0] v_12723 = 8'h0;
  wire [7:0] v_12724;
  wire [7:0] v_12725;
  function [7:0] mux_12725(input [0:0] sel);
    case (sel) 0: mux_12725 = 8'h0; 1: mux_12725 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12726;
  wire [7:0] v_12727;
  wire [7:0] v_12728;
  function [7:0] mux_12728(input [0:0] sel);
    case (sel) 0: mux_12728 = 8'h0; 1: mux_12728 = vout_peek_2083;
    endcase
  endfunction
  wire [7:0] v_12729;
  function [7:0] mux_12729(input [0:0] sel);
    case (sel) 0: mux_12729 = 8'h0; 1: mux_12729 = vout_peek_2075;
    endcase
  endfunction
  wire [7:0] v_12730;
  function [7:0] mux_12730(input [0:0] sel);
    case (sel) 0: mux_12730 = 8'h0; 1: mux_12730 = v_12731;
    endcase
  endfunction
  reg [7:0] v_12731 = 8'h0;
  wire [7:0] v_12732;
  wire [7:0] v_12733;
  function [7:0] mux_12733(input [0:0] sel);
    case (sel) 0: mux_12733 = 8'h0; 1: mux_12733 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12734;
  wire [7:0] v_12735;
  wire [7:0] v_12736;
  function [7:0] mux_12736(input [0:0] sel);
    case (sel) 0: mux_12736 = 8'h0; 1: mux_12736 = v_12737;
    endcase
  endfunction
  reg [7:0] v_12737 = 8'h0;
  wire [7:0] v_12738;
  wire [7:0] v_12739;
  function [7:0] mux_12739(input [0:0] sel);
    case (sel) 0: mux_12739 = 8'h0; 1: mux_12739 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12740;
  wire [7:0] v_12741;
  wire [7:0] v_12742;
  function [7:0] mux_12742(input [0:0] sel);
    case (sel) 0: mux_12742 = 8'h0; 1: mux_12742 = v_12743;
    endcase
  endfunction
  reg [7:0] v_12743 = 8'h0;
  wire [7:0] v_12744;
  wire [7:0] v_12745;
  function [7:0] mux_12745(input [0:0] sel);
    case (sel) 0: mux_12745 = 8'h0; 1: mux_12745 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12746;
  wire [7:0] v_12747;
  wire [7:0] v_12748;
  function [7:0] mux_12748(input [0:0] sel);
    case (sel) 0: mux_12748 = 8'h0; 1: mux_12748 = vout_peek_2069;
    endcase
  endfunction
  wire [7:0] v_12749;
  function [7:0] mux_12749(input [0:0] sel);
    case (sel) 0: mux_12749 = 8'h0; 1: mux_12749 = vout_peek_2061;
    endcase
  endfunction
  wire [7:0] v_12750;
  function [7:0] mux_12750(input [0:0] sel);
    case (sel) 0: mux_12750 = 8'h0; 1: mux_12750 = v_12751;
    endcase
  endfunction
  reg [7:0] v_12751 = 8'h0;
  wire [7:0] v_12752;
  wire [7:0] v_12753;
  function [7:0] mux_12753(input [0:0] sel);
    case (sel) 0: mux_12753 = 8'h0; 1: mux_12753 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12754;
  wire [7:0] v_12755;
  wire [7:0] v_12756;
  function [7:0] mux_12756(input [0:0] sel);
    case (sel) 0: mux_12756 = 8'h0; 1: mux_12756 = vout_peek_2055;
    endcase
  endfunction
  wire [7:0] v_12757;
  function [7:0] mux_12757(input [0:0] sel);
    case (sel) 0: mux_12757 = 8'h0; 1: mux_12757 = vout_peek_2047;
    endcase
  endfunction
  wire [7:0] v_12758;
  function [7:0] mux_12758(input [0:0] sel);
    case (sel) 0: mux_12758 = 8'h0; 1: mux_12758 = v_12759;
    endcase
  endfunction
  reg [7:0] v_12759 = 8'h0;
  wire [7:0] v_12760;
  wire [7:0] v_12761;
  function [7:0] mux_12761(input [0:0] sel);
    case (sel) 0: mux_12761 = 8'h0; 1: mux_12761 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12762;
  wire [7:0] v_12763;
  wire [7:0] v_12764;
  function [7:0] mux_12764(input [0:0] sel);
    case (sel) 0: mux_12764 = 8'h0; 1: mux_12764 = v_12765;
    endcase
  endfunction
  reg [7:0] v_12765 = 8'h0;
  wire [7:0] v_12766;
  wire [7:0] v_12767;
  function [7:0] mux_12767(input [0:0] sel);
    case (sel) 0: mux_12767 = 8'h0; 1: mux_12767 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12768;
  wire [7:0] v_12769;
  wire [7:0] v_12770;
  function [7:0] mux_12770(input [0:0] sel);
    case (sel) 0: mux_12770 = 8'h0; 1: mux_12770 = vout_peek_2041;
    endcase
  endfunction
  wire [7:0] v_12771;
  function [7:0] mux_12771(input [0:0] sel);
    case (sel) 0: mux_12771 = 8'h0; 1: mux_12771 = vout_peek_2033;
    endcase
  endfunction
  wire [7:0] v_12772;
  function [7:0] mux_12772(input [0:0] sel);
    case (sel) 0: mux_12772 = 8'h0; 1: mux_12772 = v_12773;
    endcase
  endfunction
  reg [7:0] v_12773 = 8'h0;
  wire [7:0] v_12774;
  wire [7:0] v_12775;
  function [7:0] mux_12775(input [0:0] sel);
    case (sel) 0: mux_12775 = 8'h0; 1: mux_12775 = 8'bxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_12776;
  wire [7:0] v_12777;
  wire [7:0] v_12778;
  function [7:0] mux_12778(input [0:0] sel);
    case (sel) 0: mux_12778 = 8'h0; 1: mux_12778 = vout_peek_2027;
    endcase
  endfunction
  wire [7:0] v_12779;
  function [7:0] mux_12779(input [0:0] sel);
    case (sel) 0: mux_12779 = 8'h0; 1: mux_12779 = vout_peek_2019;
    endcase
  endfunction
  wire [0:0] v_12780;
  wire [7:0] v_12781;
  // Instances
  //////////////////////////////////////////////////////////////////////////////
  assign v_0 = v_1 | v_4;
  assign v_1 = mux_1(v_2);
  assign v_2 = vout_canPeek_3 & 1'h1;
  pebbles_core
    pebbles_core_3
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_0),
       .in0_consume_en(vin0_consume_en_3),
       .out_canPeek(vout_canPeek_3),
       .out_peek(vout_peek_3));
  assign v_4 = mux_4(v_5);
  assign v_5 = ~v_2;
  assign v_6 = v_7 | v_12;
  assign v_7 = mux_7(v_8);
  assign v_8 = v_9 & 1'h1;
  assign v_9 = v_10 & vout_canPeek_11;
  assign v_10 = ~vout_canPeek_3;
  pebbles_core
    pebbles_core_11
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_6),
       .in0_consume_en(vin0_consume_en_11),
       .out_canPeek(vout_canPeek_11),
       .out_peek(vout_peek_11));
  assign v_12 = mux_12(v_13);
  assign v_13 = ~v_8;
  assign v_14 = v_15 | v_18;
  assign v_15 = mux_15(v_16);
  assign v_16 = vout_canPeek_17 & 1'h1;
  pebbles_core
    pebbles_core_17
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_14),
       .in0_consume_en(vin0_consume_en_17),
       .out_canPeek(vout_canPeek_17),
       .out_peek(vout_peek_17));
  assign v_18 = mux_18(v_19);
  assign v_19 = ~v_16;
  assign v_20 = v_21 | v_26;
  assign v_21 = mux_21(v_22);
  assign v_22 = v_23 & 1'h1;
  assign v_23 = v_24 & vout_canPeek_25;
  assign v_24 = ~vout_canPeek_17;
  pebbles_core
    pebbles_core_25
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_20),
       .in0_consume_en(vin0_consume_en_25),
       .out_canPeek(vout_canPeek_25),
       .out_peek(vout_peek_25));
  assign v_26 = mux_26(v_27);
  assign v_27 = ~v_22;
  assign v_28 = v_29 | v_32;
  assign v_29 = mux_29(v_30);
  assign v_30 = vout_canPeek_31 & 1'h1;
  pebbles_core
    pebbles_core_31
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_28),
       .in0_consume_en(vin0_consume_en_31),
       .out_canPeek(vout_canPeek_31),
       .out_peek(vout_peek_31));
  assign v_32 = mux_32(v_33);
  assign v_33 = ~v_30;
  assign v_34 = v_35 | v_40;
  assign v_35 = mux_35(v_36);
  assign v_36 = v_37 & 1'h1;
  assign v_37 = v_38 & vout_canPeek_39;
  assign v_38 = ~vout_canPeek_31;
  pebbles_core
    pebbles_core_39
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_34),
       .in0_consume_en(vin0_consume_en_39),
       .out_canPeek(vout_canPeek_39),
       .out_peek(vout_peek_39));
  assign v_40 = mux_40(v_41);
  assign v_41 = ~v_36;
  assign v_42 = v_43 | v_46;
  assign v_43 = mux_43(v_44);
  assign v_44 = vout_canPeek_45 & 1'h1;
  pebbles_core
    pebbles_core_45
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_42),
       .in0_consume_en(vin0_consume_en_45),
       .out_canPeek(vout_canPeek_45),
       .out_peek(vout_peek_45));
  assign v_46 = mux_46(v_47);
  assign v_47 = ~v_44;
  assign v_48 = v_49 | v_54;
  assign v_49 = mux_49(v_50);
  assign v_50 = v_51 & 1'h1;
  assign v_51 = v_52 & vout_canPeek_53;
  assign v_52 = ~vout_canPeek_45;
  pebbles_core
    pebbles_core_53
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_48),
       .in0_consume_en(vin0_consume_en_53),
       .out_canPeek(vout_canPeek_53),
       .out_peek(vout_peek_53));
  assign v_54 = mux_54(v_55);
  assign v_55 = ~v_50;
  assign v_56 = v_57 | v_60;
  assign v_57 = mux_57(v_58);
  assign v_58 = vout_canPeek_59 & 1'h1;
  pebbles_core
    pebbles_core_59
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_56),
       .in0_consume_en(vin0_consume_en_59),
       .out_canPeek(vout_canPeek_59),
       .out_peek(vout_peek_59));
  assign v_60 = mux_60(v_61);
  assign v_61 = ~v_58;
  assign v_62 = v_63 | v_68;
  assign v_63 = mux_63(v_64);
  assign v_64 = v_65 & 1'h1;
  assign v_65 = v_66 & vout_canPeek_67;
  assign v_66 = ~vout_canPeek_59;
  pebbles_core
    pebbles_core_67
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_62),
       .in0_consume_en(vin0_consume_en_67),
       .out_canPeek(vout_canPeek_67),
       .out_peek(vout_peek_67));
  assign v_68 = mux_68(v_69);
  assign v_69 = ~v_64;
  assign v_70 = v_71 | v_74;
  assign v_71 = mux_71(v_72);
  assign v_72 = vout_canPeek_73 & 1'h1;
  pebbles_core
    pebbles_core_73
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_70),
       .in0_consume_en(vin0_consume_en_73),
       .out_canPeek(vout_canPeek_73),
       .out_peek(vout_peek_73));
  assign v_74 = mux_74(v_75);
  assign v_75 = ~v_72;
  assign v_76 = v_77 | v_82;
  assign v_77 = mux_77(v_78);
  assign v_78 = v_79 & 1'h1;
  assign v_79 = v_80 & vout_canPeek_81;
  assign v_80 = ~vout_canPeek_73;
  pebbles_core
    pebbles_core_81
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_76),
       .in0_consume_en(vin0_consume_en_81),
       .out_canPeek(vout_canPeek_81),
       .out_peek(vout_peek_81));
  assign v_82 = mux_82(v_83);
  assign v_83 = ~v_78;
  assign v_84 = v_85 | v_88;
  assign v_85 = mux_85(v_86);
  assign v_86 = vout_canPeek_87 & 1'h1;
  pebbles_core
    pebbles_core_87
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_84),
       .in0_consume_en(vin0_consume_en_87),
       .out_canPeek(vout_canPeek_87),
       .out_peek(vout_peek_87));
  assign v_88 = mux_88(v_89);
  assign v_89 = ~v_86;
  assign v_90 = v_91 | v_96;
  assign v_91 = mux_91(v_92);
  assign v_92 = v_93 & 1'h1;
  assign v_93 = v_94 & vout_canPeek_95;
  assign v_94 = ~vout_canPeek_87;
  pebbles_core
    pebbles_core_95
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_90),
       .in0_consume_en(vin0_consume_en_95),
       .out_canPeek(vout_canPeek_95),
       .out_peek(vout_peek_95));
  assign v_96 = mux_96(v_97);
  assign v_97 = ~v_92;
  assign v_98 = v_99 | v_102;
  assign v_99 = mux_99(v_100);
  assign v_100 = vout_canPeek_101 & 1'h1;
  pebbles_core
    pebbles_core_101
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_98),
       .in0_consume_en(vin0_consume_en_101),
       .out_canPeek(vout_canPeek_101),
       .out_peek(vout_peek_101));
  assign v_102 = mux_102(v_103);
  assign v_103 = ~v_100;
  assign v_104 = v_105 | v_110;
  assign v_105 = mux_105(v_106);
  assign v_106 = v_107 & 1'h1;
  assign v_107 = v_108 & vout_canPeek_109;
  assign v_108 = ~vout_canPeek_101;
  pebbles_core
    pebbles_core_109
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_104),
       .in0_consume_en(vin0_consume_en_109),
       .out_canPeek(vout_canPeek_109),
       .out_peek(vout_peek_109));
  assign v_110 = mux_110(v_111);
  assign v_111 = ~v_106;
  assign v_112 = v_113 | v_116;
  assign v_113 = mux_113(v_114);
  assign v_114 = vout_canPeek_115 & 1'h1;
  pebbles_core
    pebbles_core_115
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_112),
       .in0_consume_en(vin0_consume_en_115),
       .out_canPeek(vout_canPeek_115),
       .out_peek(vout_peek_115));
  assign v_116 = mux_116(v_117);
  assign v_117 = ~v_114;
  assign v_118 = v_119 | v_124;
  assign v_119 = mux_119(v_120);
  assign v_120 = v_121 & 1'h1;
  assign v_121 = v_122 & vout_canPeek_123;
  assign v_122 = ~vout_canPeek_115;
  pebbles_core
    pebbles_core_123
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_118),
       .in0_consume_en(vin0_consume_en_123),
       .out_canPeek(vout_canPeek_123),
       .out_peek(vout_peek_123));
  assign v_124 = mux_124(v_125);
  assign v_125 = ~v_120;
  assign v_126 = v_127 | v_130;
  assign v_127 = mux_127(v_128);
  assign v_128 = vout_canPeek_129 & 1'h1;
  pebbles_core
    pebbles_core_129
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_126),
       .in0_consume_en(vin0_consume_en_129),
       .out_canPeek(vout_canPeek_129),
       .out_peek(vout_peek_129));
  assign v_130 = mux_130(v_131);
  assign v_131 = ~v_128;
  assign v_132 = v_133 | v_138;
  assign v_133 = mux_133(v_134);
  assign v_134 = v_135 & 1'h1;
  assign v_135 = v_136 & vout_canPeek_137;
  assign v_136 = ~vout_canPeek_129;
  pebbles_core
    pebbles_core_137
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_132),
       .in0_consume_en(vin0_consume_en_137),
       .out_canPeek(vout_canPeek_137),
       .out_peek(vout_peek_137));
  assign v_138 = mux_138(v_139);
  assign v_139 = ~v_134;
  assign v_140 = v_141 | v_144;
  assign v_141 = mux_141(v_142);
  assign v_142 = vout_canPeek_143 & 1'h1;
  pebbles_core
    pebbles_core_143
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_140),
       .in0_consume_en(vin0_consume_en_143),
       .out_canPeek(vout_canPeek_143),
       .out_peek(vout_peek_143));
  assign v_144 = mux_144(v_145);
  assign v_145 = ~v_142;
  assign v_146 = v_147 | v_152;
  assign v_147 = mux_147(v_148);
  assign v_148 = v_149 & 1'h1;
  assign v_149 = v_150 & vout_canPeek_151;
  assign v_150 = ~vout_canPeek_143;
  pebbles_core
    pebbles_core_151
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_146),
       .in0_consume_en(vin0_consume_en_151),
       .out_canPeek(vout_canPeek_151),
       .out_peek(vout_peek_151));
  assign v_152 = mux_152(v_153);
  assign v_153 = ~v_148;
  assign v_154 = v_155 | v_158;
  assign v_155 = mux_155(v_156);
  assign v_156 = vout_canPeek_157 & 1'h1;
  pebbles_core
    pebbles_core_157
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_154),
       .in0_consume_en(vin0_consume_en_157),
       .out_canPeek(vout_canPeek_157),
       .out_peek(vout_peek_157));
  assign v_158 = mux_158(v_159);
  assign v_159 = ~v_156;
  assign v_160 = v_161 | v_166;
  assign v_161 = mux_161(v_162);
  assign v_162 = v_163 & 1'h1;
  assign v_163 = v_164 & vout_canPeek_165;
  assign v_164 = ~vout_canPeek_157;
  pebbles_core
    pebbles_core_165
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_160),
       .in0_consume_en(vin0_consume_en_165),
       .out_canPeek(vout_canPeek_165),
       .out_peek(vout_peek_165));
  assign v_166 = mux_166(v_167);
  assign v_167 = ~v_162;
  assign v_168 = v_169 | v_172;
  assign v_169 = mux_169(v_170);
  assign v_170 = vout_canPeek_171 & 1'h1;
  pebbles_core
    pebbles_core_171
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_168),
       .in0_consume_en(vin0_consume_en_171),
       .out_canPeek(vout_canPeek_171),
       .out_peek(vout_peek_171));
  assign v_172 = mux_172(v_173);
  assign v_173 = ~v_170;
  assign v_174 = v_175 | v_180;
  assign v_175 = mux_175(v_176);
  assign v_176 = v_177 & 1'h1;
  assign v_177 = v_178 & vout_canPeek_179;
  assign v_178 = ~vout_canPeek_171;
  pebbles_core
    pebbles_core_179
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_174),
       .in0_consume_en(vin0_consume_en_179),
       .out_canPeek(vout_canPeek_179),
       .out_peek(vout_peek_179));
  assign v_180 = mux_180(v_181);
  assign v_181 = ~v_176;
  assign v_182 = v_183 | v_186;
  assign v_183 = mux_183(v_184);
  assign v_184 = vout_canPeek_185 & 1'h1;
  pebbles_core
    pebbles_core_185
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_182),
       .in0_consume_en(vin0_consume_en_185),
       .out_canPeek(vout_canPeek_185),
       .out_peek(vout_peek_185));
  assign v_186 = mux_186(v_187);
  assign v_187 = ~v_184;
  assign v_188 = v_189 | v_194;
  assign v_189 = mux_189(v_190);
  assign v_190 = v_191 & 1'h1;
  assign v_191 = v_192 & vout_canPeek_193;
  assign v_192 = ~vout_canPeek_185;
  pebbles_core
    pebbles_core_193
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_188),
       .in0_consume_en(vin0_consume_en_193),
       .out_canPeek(vout_canPeek_193),
       .out_peek(vout_peek_193));
  assign v_194 = mux_194(v_195);
  assign v_195 = ~v_190;
  assign v_196 = v_197 | v_200;
  assign v_197 = mux_197(v_198);
  assign v_198 = vout_canPeek_199 & 1'h1;
  pebbles_core
    pebbles_core_199
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_196),
       .in0_consume_en(vin0_consume_en_199),
       .out_canPeek(vout_canPeek_199),
       .out_peek(vout_peek_199));
  assign v_200 = mux_200(v_201);
  assign v_201 = ~v_198;
  assign v_202 = v_203 | v_208;
  assign v_203 = mux_203(v_204);
  assign v_204 = v_205 & 1'h1;
  assign v_205 = v_206 & vout_canPeek_207;
  assign v_206 = ~vout_canPeek_199;
  pebbles_core
    pebbles_core_207
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_202),
       .in0_consume_en(vin0_consume_en_207),
       .out_canPeek(vout_canPeek_207),
       .out_peek(vout_peek_207));
  assign v_208 = mux_208(v_209);
  assign v_209 = ~v_204;
  assign v_210 = v_211 | v_214;
  assign v_211 = mux_211(v_212);
  assign v_212 = vout_canPeek_213 & 1'h1;
  pebbles_core
    pebbles_core_213
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_210),
       .in0_consume_en(vin0_consume_en_213),
       .out_canPeek(vout_canPeek_213),
       .out_peek(vout_peek_213));
  assign v_214 = mux_214(v_215);
  assign v_215 = ~v_212;
  assign v_216 = v_217 | v_222;
  assign v_217 = mux_217(v_218);
  assign v_218 = v_219 & 1'h1;
  assign v_219 = v_220 & vout_canPeek_221;
  assign v_220 = ~vout_canPeek_213;
  pebbles_core
    pebbles_core_221
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_216),
       .in0_consume_en(vin0_consume_en_221),
       .out_canPeek(vout_canPeek_221),
       .out_peek(vout_peek_221));
  assign v_222 = mux_222(v_223);
  assign v_223 = ~v_218;
  assign v_224 = v_225 | v_228;
  assign v_225 = mux_225(v_226);
  assign v_226 = vout_canPeek_227 & 1'h1;
  pebbles_core
    pebbles_core_227
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_224),
       .in0_consume_en(vin0_consume_en_227),
       .out_canPeek(vout_canPeek_227),
       .out_peek(vout_peek_227));
  assign v_228 = mux_228(v_229);
  assign v_229 = ~v_226;
  assign v_230 = v_231 | v_236;
  assign v_231 = mux_231(v_232);
  assign v_232 = v_233 & 1'h1;
  assign v_233 = v_234 & vout_canPeek_235;
  assign v_234 = ~vout_canPeek_227;
  pebbles_core
    pebbles_core_235
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_230),
       .in0_consume_en(vin0_consume_en_235),
       .out_canPeek(vout_canPeek_235),
       .out_peek(vout_peek_235));
  assign v_236 = mux_236(v_237);
  assign v_237 = ~v_232;
  assign v_238 = v_239 | v_242;
  assign v_239 = mux_239(v_240);
  assign v_240 = vout_canPeek_241 & 1'h1;
  pebbles_core
    pebbles_core_241
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_238),
       .in0_consume_en(vin0_consume_en_241),
       .out_canPeek(vout_canPeek_241),
       .out_peek(vout_peek_241));
  assign v_242 = mux_242(v_243);
  assign v_243 = ~v_240;
  assign v_244 = v_245 | v_250;
  assign v_245 = mux_245(v_246);
  assign v_246 = v_247 & 1'h1;
  assign v_247 = v_248 & vout_canPeek_249;
  assign v_248 = ~vout_canPeek_241;
  pebbles_core
    pebbles_core_249
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_244),
       .in0_consume_en(vin0_consume_en_249),
       .out_canPeek(vout_canPeek_249),
       .out_peek(vout_peek_249));
  assign v_250 = mux_250(v_251);
  assign v_251 = ~v_246;
  assign v_252 = v_253 | v_256;
  assign v_253 = mux_253(v_254);
  assign v_254 = vout_canPeek_255 & 1'h1;
  pebbles_core
    pebbles_core_255
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_252),
       .in0_consume_en(vin0_consume_en_255),
       .out_canPeek(vout_canPeek_255),
       .out_peek(vout_peek_255));
  assign v_256 = mux_256(v_257);
  assign v_257 = ~v_254;
  assign v_258 = v_259 | v_264;
  assign v_259 = mux_259(v_260);
  assign v_260 = v_261 & 1'h1;
  assign v_261 = v_262 & vout_canPeek_263;
  assign v_262 = ~vout_canPeek_255;
  pebbles_core
    pebbles_core_263
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_258),
       .in0_consume_en(vin0_consume_en_263),
       .out_canPeek(vout_canPeek_263),
       .out_peek(vout_peek_263));
  assign v_264 = mux_264(v_265);
  assign v_265 = ~v_260;
  assign v_266 = v_267 | v_270;
  assign v_267 = mux_267(v_268);
  assign v_268 = vout_canPeek_269 & 1'h1;
  pebbles_core
    pebbles_core_269
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_266),
       .in0_consume_en(vin0_consume_en_269),
       .out_canPeek(vout_canPeek_269),
       .out_peek(vout_peek_269));
  assign v_270 = mux_270(v_271);
  assign v_271 = ~v_268;
  assign v_272 = v_273 | v_278;
  assign v_273 = mux_273(v_274);
  assign v_274 = v_275 & 1'h1;
  assign v_275 = v_276 & vout_canPeek_277;
  assign v_276 = ~vout_canPeek_269;
  pebbles_core
    pebbles_core_277
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_272),
       .in0_consume_en(vin0_consume_en_277),
       .out_canPeek(vout_canPeek_277),
       .out_peek(vout_peek_277));
  assign v_278 = mux_278(v_279);
  assign v_279 = ~v_274;
  assign v_280 = v_281 | v_284;
  assign v_281 = mux_281(v_282);
  assign v_282 = vout_canPeek_283 & 1'h1;
  pebbles_core
    pebbles_core_283
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_280),
       .in0_consume_en(vin0_consume_en_283),
       .out_canPeek(vout_canPeek_283),
       .out_peek(vout_peek_283));
  assign v_284 = mux_284(v_285);
  assign v_285 = ~v_282;
  assign v_286 = v_287 | v_292;
  assign v_287 = mux_287(v_288);
  assign v_288 = v_289 & 1'h1;
  assign v_289 = v_290 & vout_canPeek_291;
  assign v_290 = ~vout_canPeek_283;
  pebbles_core
    pebbles_core_291
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_286),
       .in0_consume_en(vin0_consume_en_291),
       .out_canPeek(vout_canPeek_291),
       .out_peek(vout_peek_291));
  assign v_292 = mux_292(v_293);
  assign v_293 = ~v_288;
  assign v_294 = v_295 | v_298;
  assign v_295 = mux_295(v_296);
  assign v_296 = vout_canPeek_297 & 1'h1;
  pebbles_core
    pebbles_core_297
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_294),
       .in0_consume_en(vin0_consume_en_297),
       .out_canPeek(vout_canPeek_297),
       .out_peek(vout_peek_297));
  assign v_298 = mux_298(v_299);
  assign v_299 = ~v_296;
  assign v_300 = v_301 | v_306;
  assign v_301 = mux_301(v_302);
  assign v_302 = v_303 & 1'h1;
  assign v_303 = v_304 & vout_canPeek_305;
  assign v_304 = ~vout_canPeek_297;
  pebbles_core
    pebbles_core_305
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_300),
       .in0_consume_en(vin0_consume_en_305),
       .out_canPeek(vout_canPeek_305),
       .out_peek(vout_peek_305));
  assign v_306 = mux_306(v_307);
  assign v_307 = ~v_302;
  assign v_308 = v_309 | v_312;
  assign v_309 = mux_309(v_310);
  assign v_310 = vout_canPeek_311 & 1'h1;
  pebbles_core
    pebbles_core_311
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_308),
       .in0_consume_en(vin0_consume_en_311),
       .out_canPeek(vout_canPeek_311),
       .out_peek(vout_peek_311));
  assign v_312 = mux_312(v_313);
  assign v_313 = ~v_310;
  assign v_314 = v_315 | v_320;
  assign v_315 = mux_315(v_316);
  assign v_316 = v_317 & 1'h1;
  assign v_317 = v_318 & vout_canPeek_319;
  assign v_318 = ~vout_canPeek_311;
  pebbles_core
    pebbles_core_319
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_314),
       .in0_consume_en(vin0_consume_en_319),
       .out_canPeek(vout_canPeek_319),
       .out_peek(vout_peek_319));
  assign v_320 = mux_320(v_321);
  assign v_321 = ~v_316;
  assign v_322 = v_323 | v_326;
  assign v_323 = mux_323(v_324);
  assign v_324 = vout_canPeek_325 & 1'h1;
  pebbles_core
    pebbles_core_325
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_322),
       .in0_consume_en(vin0_consume_en_325),
       .out_canPeek(vout_canPeek_325),
       .out_peek(vout_peek_325));
  assign v_326 = mux_326(v_327);
  assign v_327 = ~v_324;
  assign v_328 = v_329 | v_334;
  assign v_329 = mux_329(v_330);
  assign v_330 = v_331 & 1'h1;
  assign v_331 = v_332 & vout_canPeek_333;
  assign v_332 = ~vout_canPeek_325;
  pebbles_core
    pebbles_core_333
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_328),
       .in0_consume_en(vin0_consume_en_333),
       .out_canPeek(vout_canPeek_333),
       .out_peek(vout_peek_333));
  assign v_334 = mux_334(v_335);
  assign v_335 = ~v_330;
  assign v_336 = v_337 | v_340;
  assign v_337 = mux_337(v_338);
  assign v_338 = vout_canPeek_339 & 1'h1;
  pebbles_core
    pebbles_core_339
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_336),
       .in0_consume_en(vin0_consume_en_339),
       .out_canPeek(vout_canPeek_339),
       .out_peek(vout_peek_339));
  assign v_340 = mux_340(v_341);
  assign v_341 = ~v_338;
  assign v_342 = v_343 | v_348;
  assign v_343 = mux_343(v_344);
  assign v_344 = v_345 & 1'h1;
  assign v_345 = v_346 & vout_canPeek_347;
  assign v_346 = ~vout_canPeek_339;
  pebbles_core
    pebbles_core_347
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_342),
       .in0_consume_en(vin0_consume_en_347),
       .out_canPeek(vout_canPeek_347),
       .out_peek(vout_peek_347));
  assign v_348 = mux_348(v_349);
  assign v_349 = ~v_344;
  assign v_350 = v_351 | v_354;
  assign v_351 = mux_351(v_352);
  assign v_352 = vout_canPeek_353 & 1'h1;
  pebbles_core
    pebbles_core_353
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_350),
       .in0_consume_en(vin0_consume_en_353),
       .out_canPeek(vout_canPeek_353),
       .out_peek(vout_peek_353));
  assign v_354 = mux_354(v_355);
  assign v_355 = ~v_352;
  assign v_356 = v_357 | v_362;
  assign v_357 = mux_357(v_358);
  assign v_358 = v_359 & 1'h1;
  assign v_359 = v_360 & vout_canPeek_361;
  assign v_360 = ~vout_canPeek_353;
  pebbles_core
    pebbles_core_361
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_356),
       .in0_consume_en(vin0_consume_en_361),
       .out_canPeek(vout_canPeek_361),
       .out_peek(vout_peek_361));
  assign v_362 = mux_362(v_363);
  assign v_363 = ~v_358;
  assign v_364 = v_365 | v_368;
  assign v_365 = mux_365(v_366);
  assign v_366 = vout_canPeek_367 & 1'h1;
  pebbles_core
    pebbles_core_367
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_364),
       .in0_consume_en(vin0_consume_en_367),
       .out_canPeek(vout_canPeek_367),
       .out_peek(vout_peek_367));
  assign v_368 = mux_368(v_369);
  assign v_369 = ~v_366;
  assign v_370 = v_371 | v_376;
  assign v_371 = mux_371(v_372);
  assign v_372 = v_373 & 1'h1;
  assign v_373 = v_374 & vout_canPeek_375;
  assign v_374 = ~vout_canPeek_367;
  pebbles_core
    pebbles_core_375
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_370),
       .in0_consume_en(vin0_consume_en_375),
       .out_canPeek(vout_canPeek_375),
       .out_peek(vout_peek_375));
  assign v_376 = mux_376(v_377);
  assign v_377 = ~v_372;
  assign v_378 = v_379 | v_382;
  assign v_379 = mux_379(v_380);
  assign v_380 = vout_canPeek_381 & 1'h1;
  pebbles_core
    pebbles_core_381
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_378),
       .in0_consume_en(vin0_consume_en_381),
       .out_canPeek(vout_canPeek_381),
       .out_peek(vout_peek_381));
  assign v_382 = mux_382(v_383);
  assign v_383 = ~v_380;
  assign v_384 = v_385 | v_390;
  assign v_385 = mux_385(v_386);
  assign v_386 = v_387 & 1'h1;
  assign v_387 = v_388 & vout_canPeek_389;
  assign v_388 = ~vout_canPeek_381;
  pebbles_core
    pebbles_core_389
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_384),
       .in0_consume_en(vin0_consume_en_389),
       .out_canPeek(vout_canPeek_389),
       .out_peek(vout_peek_389));
  assign v_390 = mux_390(v_391);
  assign v_391 = ~v_386;
  assign v_392 = v_393 | v_396;
  assign v_393 = mux_393(v_394);
  assign v_394 = vout_canPeek_395 & 1'h1;
  pebbles_core
    pebbles_core_395
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_392),
       .in0_consume_en(vin0_consume_en_395),
       .out_canPeek(vout_canPeek_395),
       .out_peek(vout_peek_395));
  assign v_396 = mux_396(v_397);
  assign v_397 = ~v_394;
  assign v_398 = v_399 | v_404;
  assign v_399 = mux_399(v_400);
  assign v_400 = v_401 & 1'h1;
  assign v_401 = v_402 & vout_canPeek_403;
  assign v_402 = ~vout_canPeek_395;
  pebbles_core
    pebbles_core_403
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_398),
       .in0_consume_en(vin0_consume_en_403),
       .out_canPeek(vout_canPeek_403),
       .out_peek(vout_peek_403));
  assign v_404 = mux_404(v_405);
  assign v_405 = ~v_400;
  assign v_406 = v_407 | v_410;
  assign v_407 = mux_407(v_408);
  assign v_408 = vout_canPeek_409 & 1'h1;
  pebbles_core
    pebbles_core_409
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_406),
       .in0_consume_en(vin0_consume_en_409),
       .out_canPeek(vout_canPeek_409),
       .out_peek(vout_peek_409));
  assign v_410 = mux_410(v_411);
  assign v_411 = ~v_408;
  assign v_412 = v_413 | v_418;
  assign v_413 = mux_413(v_414);
  assign v_414 = v_415 & 1'h1;
  assign v_415 = v_416 & vout_canPeek_417;
  assign v_416 = ~vout_canPeek_409;
  pebbles_core
    pebbles_core_417
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_412),
       .in0_consume_en(vin0_consume_en_417),
       .out_canPeek(vout_canPeek_417),
       .out_peek(vout_peek_417));
  assign v_418 = mux_418(v_419);
  assign v_419 = ~v_414;
  assign v_420 = v_421 | v_424;
  assign v_421 = mux_421(v_422);
  assign v_422 = vout_canPeek_423 & 1'h1;
  pebbles_core
    pebbles_core_423
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_420),
       .in0_consume_en(vin0_consume_en_423),
       .out_canPeek(vout_canPeek_423),
       .out_peek(vout_peek_423));
  assign v_424 = mux_424(v_425);
  assign v_425 = ~v_422;
  assign v_426 = v_427 | v_432;
  assign v_427 = mux_427(v_428);
  assign v_428 = v_429 & 1'h1;
  assign v_429 = v_430 & vout_canPeek_431;
  assign v_430 = ~vout_canPeek_423;
  pebbles_core
    pebbles_core_431
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_426),
       .in0_consume_en(vin0_consume_en_431),
       .out_canPeek(vout_canPeek_431),
       .out_peek(vout_peek_431));
  assign v_432 = mux_432(v_433);
  assign v_433 = ~v_428;
  assign v_434 = v_435 | v_438;
  assign v_435 = mux_435(v_436);
  assign v_436 = vout_canPeek_437 & 1'h1;
  pebbles_core
    pebbles_core_437
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_434),
       .in0_consume_en(vin0_consume_en_437),
       .out_canPeek(vout_canPeek_437),
       .out_peek(vout_peek_437));
  assign v_438 = mux_438(v_439);
  assign v_439 = ~v_436;
  assign v_440 = v_441 | v_446;
  assign v_441 = mux_441(v_442);
  assign v_442 = v_443 & 1'h1;
  assign v_443 = v_444 & vout_canPeek_445;
  assign v_444 = ~vout_canPeek_437;
  pebbles_core
    pebbles_core_445
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_440),
       .in0_consume_en(vin0_consume_en_445),
       .out_canPeek(vout_canPeek_445),
       .out_peek(vout_peek_445));
  assign v_446 = mux_446(v_447);
  assign v_447 = ~v_442;
  assign v_448 = v_449 | v_452;
  assign v_449 = mux_449(v_450);
  assign v_450 = vout_canPeek_451 & 1'h1;
  pebbles_core
    pebbles_core_451
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_448),
       .in0_consume_en(vin0_consume_en_451),
       .out_canPeek(vout_canPeek_451),
       .out_peek(vout_peek_451));
  assign v_452 = mux_452(v_453);
  assign v_453 = ~v_450;
  assign v_454 = v_455 | v_460;
  assign v_455 = mux_455(v_456);
  assign v_456 = v_457 & 1'h1;
  assign v_457 = v_458 & vout_canPeek_459;
  assign v_458 = ~vout_canPeek_451;
  pebbles_core
    pebbles_core_459
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_454),
       .in0_consume_en(vin0_consume_en_459),
       .out_canPeek(vout_canPeek_459),
       .out_peek(vout_peek_459));
  assign v_460 = mux_460(v_461);
  assign v_461 = ~v_456;
  assign v_462 = v_463 | v_466;
  assign v_463 = mux_463(v_464);
  assign v_464 = vout_canPeek_465 & 1'h1;
  pebbles_core
    pebbles_core_465
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_462),
       .in0_consume_en(vin0_consume_en_465),
       .out_canPeek(vout_canPeek_465),
       .out_peek(vout_peek_465));
  assign v_466 = mux_466(v_467);
  assign v_467 = ~v_464;
  assign v_468 = v_469 | v_474;
  assign v_469 = mux_469(v_470);
  assign v_470 = v_471 & 1'h1;
  assign v_471 = v_472 & vout_canPeek_473;
  assign v_472 = ~vout_canPeek_465;
  pebbles_core
    pebbles_core_473
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_468),
       .in0_consume_en(vin0_consume_en_473),
       .out_canPeek(vout_canPeek_473),
       .out_peek(vout_peek_473));
  assign v_474 = mux_474(v_475);
  assign v_475 = ~v_470;
  assign v_476 = v_477 | v_480;
  assign v_477 = mux_477(v_478);
  assign v_478 = vout_canPeek_479 & 1'h1;
  pebbles_core
    pebbles_core_479
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_476),
       .in0_consume_en(vin0_consume_en_479),
       .out_canPeek(vout_canPeek_479),
       .out_peek(vout_peek_479));
  assign v_480 = mux_480(v_481);
  assign v_481 = ~v_478;
  assign v_482 = v_483 | v_488;
  assign v_483 = mux_483(v_484);
  assign v_484 = v_485 & 1'h1;
  assign v_485 = v_486 & vout_canPeek_487;
  assign v_486 = ~vout_canPeek_479;
  pebbles_core
    pebbles_core_487
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_482),
       .in0_consume_en(vin0_consume_en_487),
       .out_canPeek(vout_canPeek_487),
       .out_peek(vout_peek_487));
  assign v_488 = mux_488(v_489);
  assign v_489 = ~v_484;
  assign v_490 = v_491 | v_494;
  assign v_491 = mux_491(v_492);
  assign v_492 = vout_canPeek_493 & 1'h1;
  pebbles_core
    pebbles_core_493
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_490),
       .in0_consume_en(vin0_consume_en_493),
       .out_canPeek(vout_canPeek_493),
       .out_peek(vout_peek_493));
  assign v_494 = mux_494(v_495);
  assign v_495 = ~v_492;
  assign v_496 = v_497 | v_502;
  assign v_497 = mux_497(v_498);
  assign v_498 = v_499 & 1'h1;
  assign v_499 = v_500 & vout_canPeek_501;
  assign v_500 = ~vout_canPeek_493;
  pebbles_core
    pebbles_core_501
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_496),
       .in0_consume_en(vin0_consume_en_501),
       .out_canPeek(vout_canPeek_501),
       .out_peek(vout_peek_501));
  assign v_502 = mux_502(v_503);
  assign v_503 = ~v_498;
  assign v_504 = v_505 | v_508;
  assign v_505 = mux_505(v_506);
  assign v_506 = vout_canPeek_507 & 1'h1;
  pebbles_core
    pebbles_core_507
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_504),
       .in0_consume_en(vin0_consume_en_507),
       .out_canPeek(vout_canPeek_507),
       .out_peek(vout_peek_507));
  assign v_508 = mux_508(v_509);
  assign v_509 = ~v_506;
  assign v_510 = v_511 | v_516;
  assign v_511 = mux_511(v_512);
  assign v_512 = v_513 & 1'h1;
  assign v_513 = v_514 & vout_canPeek_515;
  assign v_514 = ~vout_canPeek_507;
  pebbles_core
    pebbles_core_515
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_510),
       .in0_consume_en(vin0_consume_en_515),
       .out_canPeek(vout_canPeek_515),
       .out_peek(vout_peek_515));
  assign v_516 = mux_516(v_517);
  assign v_517 = ~v_512;
  assign v_518 = v_519 | v_522;
  assign v_519 = mux_519(v_520);
  assign v_520 = vout_canPeek_521 & 1'h1;
  pebbles_core
    pebbles_core_521
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_518),
       .in0_consume_en(vin0_consume_en_521),
       .out_canPeek(vout_canPeek_521),
       .out_peek(vout_peek_521));
  assign v_522 = mux_522(v_523);
  assign v_523 = ~v_520;
  assign v_524 = v_525 | v_530;
  assign v_525 = mux_525(v_526);
  assign v_526 = v_527 & 1'h1;
  assign v_527 = v_528 & vout_canPeek_529;
  assign v_528 = ~vout_canPeek_521;
  pebbles_core
    pebbles_core_529
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_524),
       .in0_consume_en(vin0_consume_en_529),
       .out_canPeek(vout_canPeek_529),
       .out_peek(vout_peek_529));
  assign v_530 = mux_530(v_531);
  assign v_531 = ~v_526;
  assign v_532 = v_533 | v_536;
  assign v_533 = mux_533(v_534);
  assign v_534 = vout_canPeek_535 & 1'h1;
  pebbles_core
    pebbles_core_535
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_532),
       .in0_consume_en(vin0_consume_en_535),
       .out_canPeek(vout_canPeek_535),
       .out_peek(vout_peek_535));
  assign v_536 = mux_536(v_537);
  assign v_537 = ~v_534;
  assign v_538 = v_539 | v_544;
  assign v_539 = mux_539(v_540);
  assign v_540 = v_541 & 1'h1;
  assign v_541 = v_542 & vout_canPeek_543;
  assign v_542 = ~vout_canPeek_535;
  pebbles_core
    pebbles_core_543
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_538),
       .in0_consume_en(vin0_consume_en_543),
       .out_canPeek(vout_canPeek_543),
       .out_peek(vout_peek_543));
  assign v_544 = mux_544(v_545);
  assign v_545 = ~v_540;
  assign v_546 = v_547 | v_550;
  assign v_547 = mux_547(v_548);
  assign v_548 = vout_canPeek_549 & 1'h1;
  pebbles_core
    pebbles_core_549
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_546),
       .in0_consume_en(vin0_consume_en_549),
       .out_canPeek(vout_canPeek_549),
       .out_peek(vout_peek_549));
  assign v_550 = mux_550(v_551);
  assign v_551 = ~v_548;
  assign v_552 = v_553 | v_558;
  assign v_553 = mux_553(v_554);
  assign v_554 = v_555 & 1'h1;
  assign v_555 = v_556 & vout_canPeek_557;
  assign v_556 = ~vout_canPeek_549;
  pebbles_core
    pebbles_core_557
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_552),
       .in0_consume_en(vin0_consume_en_557),
       .out_canPeek(vout_canPeek_557),
       .out_peek(vout_peek_557));
  assign v_558 = mux_558(v_559);
  assign v_559 = ~v_554;
  assign v_560 = v_561 | v_564;
  assign v_561 = mux_561(v_562);
  assign v_562 = vout_canPeek_563 & 1'h1;
  pebbles_core
    pebbles_core_563
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_560),
       .in0_consume_en(vin0_consume_en_563),
       .out_canPeek(vout_canPeek_563),
       .out_peek(vout_peek_563));
  assign v_564 = mux_564(v_565);
  assign v_565 = ~v_562;
  assign v_566 = v_567 | v_572;
  assign v_567 = mux_567(v_568);
  assign v_568 = v_569 & 1'h1;
  assign v_569 = v_570 & vout_canPeek_571;
  assign v_570 = ~vout_canPeek_563;
  pebbles_core
    pebbles_core_571
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_566),
       .in0_consume_en(vin0_consume_en_571),
       .out_canPeek(vout_canPeek_571),
       .out_peek(vout_peek_571));
  assign v_572 = mux_572(v_573);
  assign v_573 = ~v_568;
  assign v_574 = v_575 | v_578;
  assign v_575 = mux_575(v_576);
  assign v_576 = vout_canPeek_577 & 1'h1;
  pebbles_core
    pebbles_core_577
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_574),
       .in0_consume_en(vin0_consume_en_577),
       .out_canPeek(vout_canPeek_577),
       .out_peek(vout_peek_577));
  assign v_578 = mux_578(v_579);
  assign v_579 = ~v_576;
  assign v_580 = v_581 | v_586;
  assign v_581 = mux_581(v_582);
  assign v_582 = v_583 & 1'h1;
  assign v_583 = v_584 & vout_canPeek_585;
  assign v_584 = ~vout_canPeek_577;
  pebbles_core
    pebbles_core_585
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_580),
       .in0_consume_en(vin0_consume_en_585),
       .out_canPeek(vout_canPeek_585),
       .out_peek(vout_peek_585));
  assign v_586 = mux_586(v_587);
  assign v_587 = ~v_582;
  assign v_588 = v_589 | v_592;
  assign v_589 = mux_589(v_590);
  assign v_590 = vout_canPeek_591 & 1'h1;
  pebbles_core
    pebbles_core_591
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_588),
       .in0_consume_en(vin0_consume_en_591),
       .out_canPeek(vout_canPeek_591),
       .out_peek(vout_peek_591));
  assign v_592 = mux_592(v_593);
  assign v_593 = ~v_590;
  assign v_594 = v_595 | v_600;
  assign v_595 = mux_595(v_596);
  assign v_596 = v_597 & 1'h1;
  assign v_597 = v_598 & vout_canPeek_599;
  assign v_598 = ~vout_canPeek_591;
  pebbles_core
    pebbles_core_599
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_594),
       .in0_consume_en(vin0_consume_en_599),
       .out_canPeek(vout_canPeek_599),
       .out_peek(vout_peek_599));
  assign v_600 = mux_600(v_601);
  assign v_601 = ~v_596;
  assign v_602 = v_603 | v_606;
  assign v_603 = mux_603(v_604);
  assign v_604 = vout_canPeek_605 & 1'h1;
  pebbles_core
    pebbles_core_605
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_602),
       .in0_consume_en(vin0_consume_en_605),
       .out_canPeek(vout_canPeek_605),
       .out_peek(vout_peek_605));
  assign v_606 = mux_606(v_607);
  assign v_607 = ~v_604;
  assign v_608 = v_609 | v_614;
  assign v_609 = mux_609(v_610);
  assign v_610 = v_611 & 1'h1;
  assign v_611 = v_612 & vout_canPeek_613;
  assign v_612 = ~vout_canPeek_605;
  pebbles_core
    pebbles_core_613
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_608),
       .in0_consume_en(vin0_consume_en_613),
       .out_canPeek(vout_canPeek_613),
       .out_peek(vout_peek_613));
  assign v_614 = mux_614(v_615);
  assign v_615 = ~v_610;
  assign v_616 = v_617 | v_620;
  assign v_617 = mux_617(v_618);
  assign v_618 = vout_canPeek_619 & 1'h1;
  pebbles_core
    pebbles_core_619
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_616),
       .in0_consume_en(vin0_consume_en_619),
       .out_canPeek(vout_canPeek_619),
       .out_peek(vout_peek_619));
  assign v_620 = mux_620(v_621);
  assign v_621 = ~v_618;
  assign v_622 = v_623 | v_628;
  assign v_623 = mux_623(v_624);
  assign v_624 = v_625 & 1'h1;
  assign v_625 = v_626 & vout_canPeek_627;
  assign v_626 = ~vout_canPeek_619;
  pebbles_core
    pebbles_core_627
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_622),
       .in0_consume_en(vin0_consume_en_627),
       .out_canPeek(vout_canPeek_627),
       .out_peek(vout_peek_627));
  assign v_628 = mux_628(v_629);
  assign v_629 = ~v_624;
  assign v_630 = v_631 | v_634;
  assign v_631 = mux_631(v_632);
  assign v_632 = vout_canPeek_633 & 1'h1;
  pebbles_core
    pebbles_core_633
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_630),
       .in0_consume_en(vin0_consume_en_633),
       .out_canPeek(vout_canPeek_633),
       .out_peek(vout_peek_633));
  assign v_634 = mux_634(v_635);
  assign v_635 = ~v_632;
  assign v_636 = v_637 | v_642;
  assign v_637 = mux_637(v_638);
  assign v_638 = v_639 & 1'h1;
  assign v_639 = v_640 & vout_canPeek_641;
  assign v_640 = ~vout_canPeek_633;
  pebbles_core
    pebbles_core_641
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_636),
       .in0_consume_en(vin0_consume_en_641),
       .out_canPeek(vout_canPeek_641),
       .out_peek(vout_peek_641));
  assign v_642 = mux_642(v_643);
  assign v_643 = ~v_638;
  assign v_644 = v_645 | v_648;
  assign v_645 = mux_645(v_646);
  assign v_646 = vout_canPeek_647 & 1'h1;
  pebbles_core
    pebbles_core_647
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_644),
       .in0_consume_en(vin0_consume_en_647),
       .out_canPeek(vout_canPeek_647),
       .out_peek(vout_peek_647));
  assign v_648 = mux_648(v_649);
  assign v_649 = ~v_646;
  assign v_650 = v_651 | v_656;
  assign v_651 = mux_651(v_652);
  assign v_652 = v_653 & 1'h1;
  assign v_653 = v_654 & vout_canPeek_655;
  assign v_654 = ~vout_canPeek_647;
  pebbles_core
    pebbles_core_655
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_650),
       .in0_consume_en(vin0_consume_en_655),
       .out_canPeek(vout_canPeek_655),
       .out_peek(vout_peek_655));
  assign v_656 = mux_656(v_657);
  assign v_657 = ~v_652;
  assign v_658 = v_659 | v_662;
  assign v_659 = mux_659(v_660);
  assign v_660 = vout_canPeek_661 & 1'h1;
  pebbles_core
    pebbles_core_661
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_658),
       .in0_consume_en(vin0_consume_en_661),
       .out_canPeek(vout_canPeek_661),
       .out_peek(vout_peek_661));
  assign v_662 = mux_662(v_663);
  assign v_663 = ~v_660;
  assign v_664 = v_665 | v_670;
  assign v_665 = mux_665(v_666);
  assign v_666 = v_667 & 1'h1;
  assign v_667 = v_668 & vout_canPeek_669;
  assign v_668 = ~vout_canPeek_661;
  pebbles_core
    pebbles_core_669
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_664),
       .in0_consume_en(vin0_consume_en_669),
       .out_canPeek(vout_canPeek_669),
       .out_peek(vout_peek_669));
  assign v_670 = mux_670(v_671);
  assign v_671 = ~v_666;
  assign v_672 = v_673 | v_676;
  assign v_673 = mux_673(v_674);
  assign v_674 = vout_canPeek_675 & 1'h1;
  pebbles_core
    pebbles_core_675
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_672),
       .in0_consume_en(vin0_consume_en_675),
       .out_canPeek(vout_canPeek_675),
       .out_peek(vout_peek_675));
  assign v_676 = mux_676(v_677);
  assign v_677 = ~v_674;
  assign v_678 = v_679 | v_684;
  assign v_679 = mux_679(v_680);
  assign v_680 = v_681 & 1'h1;
  assign v_681 = v_682 & vout_canPeek_683;
  assign v_682 = ~vout_canPeek_675;
  pebbles_core
    pebbles_core_683
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_678),
       .in0_consume_en(vin0_consume_en_683),
       .out_canPeek(vout_canPeek_683),
       .out_peek(vout_peek_683));
  assign v_684 = mux_684(v_685);
  assign v_685 = ~v_680;
  assign v_686 = v_687 | v_690;
  assign v_687 = mux_687(v_688);
  assign v_688 = vout_canPeek_689 & 1'h1;
  pebbles_core
    pebbles_core_689
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_686),
       .in0_consume_en(vin0_consume_en_689),
       .out_canPeek(vout_canPeek_689),
       .out_peek(vout_peek_689));
  assign v_690 = mux_690(v_691);
  assign v_691 = ~v_688;
  assign v_692 = v_693 | v_698;
  assign v_693 = mux_693(v_694);
  assign v_694 = v_695 & 1'h1;
  assign v_695 = v_696 & vout_canPeek_697;
  assign v_696 = ~vout_canPeek_689;
  pebbles_core
    pebbles_core_697
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_692),
       .in0_consume_en(vin0_consume_en_697),
       .out_canPeek(vout_canPeek_697),
       .out_peek(vout_peek_697));
  assign v_698 = mux_698(v_699);
  assign v_699 = ~v_694;
  assign v_700 = v_701 | v_704;
  assign v_701 = mux_701(v_702);
  assign v_702 = vout_canPeek_703 & 1'h1;
  pebbles_core
    pebbles_core_703
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_700),
       .in0_consume_en(vin0_consume_en_703),
       .out_canPeek(vout_canPeek_703),
       .out_peek(vout_peek_703));
  assign v_704 = mux_704(v_705);
  assign v_705 = ~v_702;
  assign v_706 = v_707 | v_712;
  assign v_707 = mux_707(v_708);
  assign v_708 = v_709 & 1'h1;
  assign v_709 = v_710 & vout_canPeek_711;
  assign v_710 = ~vout_canPeek_703;
  pebbles_core
    pebbles_core_711
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_706),
       .in0_consume_en(vin0_consume_en_711),
       .out_canPeek(vout_canPeek_711),
       .out_peek(vout_peek_711));
  assign v_712 = mux_712(v_713);
  assign v_713 = ~v_708;
  assign v_714 = v_715 | v_718;
  assign v_715 = mux_715(v_716);
  assign v_716 = vout_canPeek_717 & 1'h1;
  pebbles_core
    pebbles_core_717
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_714),
       .in0_consume_en(vin0_consume_en_717),
       .out_canPeek(vout_canPeek_717),
       .out_peek(vout_peek_717));
  assign v_718 = mux_718(v_719);
  assign v_719 = ~v_716;
  assign v_720 = v_721 | v_726;
  assign v_721 = mux_721(v_722);
  assign v_722 = v_723 & 1'h1;
  assign v_723 = v_724 & vout_canPeek_725;
  assign v_724 = ~vout_canPeek_717;
  pebbles_core
    pebbles_core_725
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_720),
       .in0_consume_en(vin0_consume_en_725),
       .out_canPeek(vout_canPeek_725),
       .out_peek(vout_peek_725));
  assign v_726 = mux_726(v_727);
  assign v_727 = ~v_722;
  assign v_728 = v_729 | v_732;
  assign v_729 = mux_729(v_730);
  assign v_730 = vout_canPeek_731 & 1'h1;
  pebbles_core
    pebbles_core_731
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_728),
       .in0_consume_en(vin0_consume_en_731),
       .out_canPeek(vout_canPeek_731),
       .out_peek(vout_peek_731));
  assign v_732 = mux_732(v_733);
  assign v_733 = ~v_730;
  assign v_734 = v_735 | v_740;
  assign v_735 = mux_735(v_736);
  assign v_736 = v_737 & 1'h1;
  assign v_737 = v_738 & vout_canPeek_739;
  assign v_738 = ~vout_canPeek_731;
  pebbles_core
    pebbles_core_739
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_734),
       .in0_consume_en(vin0_consume_en_739),
       .out_canPeek(vout_canPeek_739),
       .out_peek(vout_peek_739));
  assign v_740 = mux_740(v_741);
  assign v_741 = ~v_736;
  assign v_742 = v_743 | v_746;
  assign v_743 = mux_743(v_744);
  assign v_744 = vout_canPeek_745 & 1'h1;
  pebbles_core
    pebbles_core_745
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_742),
       .in0_consume_en(vin0_consume_en_745),
       .out_canPeek(vout_canPeek_745),
       .out_peek(vout_peek_745));
  assign v_746 = mux_746(v_747);
  assign v_747 = ~v_744;
  assign v_748 = v_749 | v_754;
  assign v_749 = mux_749(v_750);
  assign v_750 = v_751 & 1'h1;
  assign v_751 = v_752 & vout_canPeek_753;
  assign v_752 = ~vout_canPeek_745;
  pebbles_core
    pebbles_core_753
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_748),
       .in0_consume_en(vin0_consume_en_753),
       .out_canPeek(vout_canPeek_753),
       .out_peek(vout_peek_753));
  assign v_754 = mux_754(v_755);
  assign v_755 = ~v_750;
  assign v_756 = v_757 | v_760;
  assign v_757 = mux_757(v_758);
  assign v_758 = vout_canPeek_759 & 1'h1;
  pebbles_core
    pebbles_core_759
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_756),
       .in0_consume_en(vin0_consume_en_759),
       .out_canPeek(vout_canPeek_759),
       .out_peek(vout_peek_759));
  assign v_760 = mux_760(v_761);
  assign v_761 = ~v_758;
  assign v_762 = v_763 | v_768;
  assign v_763 = mux_763(v_764);
  assign v_764 = v_765 & 1'h1;
  assign v_765 = v_766 & vout_canPeek_767;
  assign v_766 = ~vout_canPeek_759;
  pebbles_core
    pebbles_core_767
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_762),
       .in0_consume_en(vin0_consume_en_767),
       .out_canPeek(vout_canPeek_767),
       .out_peek(vout_peek_767));
  assign v_768 = mux_768(v_769);
  assign v_769 = ~v_764;
  assign v_770 = v_771 | v_774;
  assign v_771 = mux_771(v_772);
  assign v_772 = vout_canPeek_773 & 1'h1;
  pebbles_core
    pebbles_core_773
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_770),
       .in0_consume_en(vin0_consume_en_773),
       .out_canPeek(vout_canPeek_773),
       .out_peek(vout_peek_773));
  assign v_774 = mux_774(v_775);
  assign v_775 = ~v_772;
  assign v_776 = v_777 | v_782;
  assign v_777 = mux_777(v_778);
  assign v_778 = v_779 & 1'h1;
  assign v_779 = v_780 & vout_canPeek_781;
  assign v_780 = ~vout_canPeek_773;
  pebbles_core
    pebbles_core_781
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_776),
       .in0_consume_en(vin0_consume_en_781),
       .out_canPeek(vout_canPeek_781),
       .out_peek(vout_peek_781));
  assign v_782 = mux_782(v_783);
  assign v_783 = ~v_778;
  assign v_784 = v_785 | v_788;
  assign v_785 = mux_785(v_786);
  assign v_786 = vout_canPeek_787 & 1'h1;
  pebbles_core
    pebbles_core_787
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_784),
       .in0_consume_en(vin0_consume_en_787),
       .out_canPeek(vout_canPeek_787),
       .out_peek(vout_peek_787));
  assign v_788 = mux_788(v_789);
  assign v_789 = ~v_786;
  assign v_790 = v_791 | v_796;
  assign v_791 = mux_791(v_792);
  assign v_792 = v_793 & 1'h1;
  assign v_793 = v_794 & vout_canPeek_795;
  assign v_794 = ~vout_canPeek_787;
  pebbles_core
    pebbles_core_795
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_790),
       .in0_consume_en(vin0_consume_en_795),
       .out_canPeek(vout_canPeek_795),
       .out_peek(vout_peek_795));
  assign v_796 = mux_796(v_797);
  assign v_797 = ~v_792;
  assign v_798 = v_799 | v_802;
  assign v_799 = mux_799(v_800);
  assign v_800 = vout_canPeek_801 & 1'h1;
  pebbles_core
    pebbles_core_801
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_798),
       .in0_consume_en(vin0_consume_en_801),
       .out_canPeek(vout_canPeek_801),
       .out_peek(vout_peek_801));
  assign v_802 = mux_802(v_803);
  assign v_803 = ~v_800;
  assign v_804 = v_805 | v_810;
  assign v_805 = mux_805(v_806);
  assign v_806 = v_807 & 1'h1;
  assign v_807 = v_808 & vout_canPeek_809;
  assign v_808 = ~vout_canPeek_801;
  pebbles_core
    pebbles_core_809
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_804),
       .in0_consume_en(vin0_consume_en_809),
       .out_canPeek(vout_canPeek_809),
       .out_peek(vout_peek_809));
  assign v_810 = mux_810(v_811);
  assign v_811 = ~v_806;
  assign v_812 = v_813 | v_816;
  assign v_813 = mux_813(v_814);
  assign v_814 = vout_canPeek_815 & 1'h1;
  pebbles_core
    pebbles_core_815
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_812),
       .in0_consume_en(vin0_consume_en_815),
       .out_canPeek(vout_canPeek_815),
       .out_peek(vout_peek_815));
  assign v_816 = mux_816(v_817);
  assign v_817 = ~v_814;
  assign v_818 = v_819 | v_824;
  assign v_819 = mux_819(v_820);
  assign v_820 = v_821 & 1'h1;
  assign v_821 = v_822 & vout_canPeek_823;
  assign v_822 = ~vout_canPeek_815;
  pebbles_core
    pebbles_core_823
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_818),
       .in0_consume_en(vin0_consume_en_823),
       .out_canPeek(vout_canPeek_823),
       .out_peek(vout_peek_823));
  assign v_824 = mux_824(v_825);
  assign v_825 = ~v_820;
  assign v_826 = v_827 | v_830;
  assign v_827 = mux_827(v_828);
  assign v_828 = vout_canPeek_829 & 1'h1;
  pebbles_core
    pebbles_core_829
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_826),
       .in0_consume_en(vin0_consume_en_829),
       .out_canPeek(vout_canPeek_829),
       .out_peek(vout_peek_829));
  assign v_830 = mux_830(v_831);
  assign v_831 = ~v_828;
  assign v_832 = v_833 | v_838;
  assign v_833 = mux_833(v_834);
  assign v_834 = v_835 & 1'h1;
  assign v_835 = v_836 & vout_canPeek_837;
  assign v_836 = ~vout_canPeek_829;
  pebbles_core
    pebbles_core_837
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_832),
       .in0_consume_en(vin0_consume_en_837),
       .out_canPeek(vout_canPeek_837),
       .out_peek(vout_peek_837));
  assign v_838 = mux_838(v_839);
  assign v_839 = ~v_834;
  assign v_840 = v_841 | v_844;
  assign v_841 = mux_841(v_842);
  assign v_842 = vout_canPeek_843 & 1'h1;
  pebbles_core
    pebbles_core_843
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_840),
       .in0_consume_en(vin0_consume_en_843),
       .out_canPeek(vout_canPeek_843),
       .out_peek(vout_peek_843));
  assign v_844 = mux_844(v_845);
  assign v_845 = ~v_842;
  assign v_846 = v_847 | v_852;
  assign v_847 = mux_847(v_848);
  assign v_848 = v_849 & 1'h1;
  assign v_849 = v_850 & vout_canPeek_851;
  assign v_850 = ~vout_canPeek_843;
  pebbles_core
    pebbles_core_851
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_846),
       .in0_consume_en(vin0_consume_en_851),
       .out_canPeek(vout_canPeek_851),
       .out_peek(vout_peek_851));
  assign v_852 = mux_852(v_853);
  assign v_853 = ~v_848;
  assign v_854 = v_855 | v_858;
  assign v_855 = mux_855(v_856);
  assign v_856 = vout_canPeek_857 & 1'h1;
  pebbles_core
    pebbles_core_857
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_854),
       .in0_consume_en(vin0_consume_en_857),
       .out_canPeek(vout_canPeek_857),
       .out_peek(vout_peek_857));
  assign v_858 = mux_858(v_859);
  assign v_859 = ~v_856;
  assign v_860 = v_861 | v_866;
  assign v_861 = mux_861(v_862);
  assign v_862 = v_863 & 1'h1;
  assign v_863 = v_864 & vout_canPeek_865;
  assign v_864 = ~vout_canPeek_857;
  pebbles_core
    pebbles_core_865
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_860),
       .in0_consume_en(vin0_consume_en_865),
       .out_canPeek(vout_canPeek_865),
       .out_peek(vout_peek_865));
  assign v_866 = mux_866(v_867);
  assign v_867 = ~v_862;
  assign v_868 = v_869 | v_872;
  assign v_869 = mux_869(v_870);
  assign v_870 = vout_canPeek_871 & 1'h1;
  pebbles_core
    pebbles_core_871
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_868),
       .in0_consume_en(vin0_consume_en_871),
       .out_canPeek(vout_canPeek_871),
       .out_peek(vout_peek_871));
  assign v_872 = mux_872(v_873);
  assign v_873 = ~v_870;
  assign v_874 = v_875 | v_880;
  assign v_875 = mux_875(v_876);
  assign v_876 = v_877 & 1'h1;
  assign v_877 = v_878 & vout_canPeek_879;
  assign v_878 = ~vout_canPeek_871;
  pebbles_core
    pebbles_core_879
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_874),
       .in0_consume_en(vin0_consume_en_879),
       .out_canPeek(vout_canPeek_879),
       .out_peek(vout_peek_879));
  assign v_880 = mux_880(v_881);
  assign v_881 = ~v_876;
  assign v_882 = v_883 | v_886;
  assign v_883 = mux_883(v_884);
  assign v_884 = vout_canPeek_885 & 1'h1;
  pebbles_core
    pebbles_core_885
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_882),
       .in0_consume_en(vin0_consume_en_885),
       .out_canPeek(vout_canPeek_885),
       .out_peek(vout_peek_885));
  assign v_886 = mux_886(v_887);
  assign v_887 = ~v_884;
  assign v_888 = v_889 | v_894;
  assign v_889 = mux_889(v_890);
  assign v_890 = v_891 & 1'h1;
  assign v_891 = v_892 & vout_canPeek_893;
  assign v_892 = ~vout_canPeek_885;
  pebbles_core
    pebbles_core_893
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_888),
       .in0_consume_en(vin0_consume_en_893),
       .out_canPeek(vout_canPeek_893),
       .out_peek(vout_peek_893));
  assign v_894 = mux_894(v_895);
  assign v_895 = ~v_890;
  assign v_896 = v_897 | v_900;
  assign v_897 = mux_897(v_898);
  assign v_898 = vout_canPeek_899 & 1'h1;
  pebbles_core
    pebbles_core_899
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_896),
       .in0_consume_en(vin0_consume_en_899),
       .out_canPeek(vout_canPeek_899),
       .out_peek(vout_peek_899));
  assign v_900 = mux_900(v_901);
  assign v_901 = ~v_898;
  assign v_902 = v_903 | v_908;
  assign v_903 = mux_903(v_904);
  assign v_904 = v_905 & 1'h1;
  assign v_905 = v_906 & vout_canPeek_907;
  assign v_906 = ~vout_canPeek_899;
  pebbles_core
    pebbles_core_907
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_902),
       .in0_consume_en(vin0_consume_en_907),
       .out_canPeek(vout_canPeek_907),
       .out_peek(vout_peek_907));
  assign v_908 = mux_908(v_909);
  assign v_909 = ~v_904;
  assign v_910 = v_911 | v_914;
  assign v_911 = mux_911(v_912);
  assign v_912 = vout_canPeek_913 & 1'h1;
  pebbles_core
    pebbles_core_913
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_910),
       .in0_consume_en(vin0_consume_en_913),
       .out_canPeek(vout_canPeek_913),
       .out_peek(vout_peek_913));
  assign v_914 = mux_914(v_915);
  assign v_915 = ~v_912;
  assign v_916 = v_917 | v_922;
  assign v_917 = mux_917(v_918);
  assign v_918 = v_919 & 1'h1;
  assign v_919 = v_920 & vout_canPeek_921;
  assign v_920 = ~vout_canPeek_913;
  pebbles_core
    pebbles_core_921
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_916),
       .in0_consume_en(vin0_consume_en_921),
       .out_canPeek(vout_canPeek_921),
       .out_peek(vout_peek_921));
  assign v_922 = mux_922(v_923);
  assign v_923 = ~v_918;
  assign v_924 = v_925 | v_928;
  assign v_925 = mux_925(v_926);
  assign v_926 = vout_canPeek_927 & 1'h1;
  pebbles_core
    pebbles_core_927
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_924),
       .in0_consume_en(vin0_consume_en_927),
       .out_canPeek(vout_canPeek_927),
       .out_peek(vout_peek_927));
  assign v_928 = mux_928(v_929);
  assign v_929 = ~v_926;
  assign v_930 = v_931 | v_936;
  assign v_931 = mux_931(v_932);
  assign v_932 = v_933 & 1'h1;
  assign v_933 = v_934 & vout_canPeek_935;
  assign v_934 = ~vout_canPeek_927;
  pebbles_core
    pebbles_core_935
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_930),
       .in0_consume_en(vin0_consume_en_935),
       .out_canPeek(vout_canPeek_935),
       .out_peek(vout_peek_935));
  assign v_936 = mux_936(v_937);
  assign v_937 = ~v_932;
  assign v_938 = v_939 | v_942;
  assign v_939 = mux_939(v_940);
  assign v_940 = vout_canPeek_941 & 1'h1;
  pebbles_core
    pebbles_core_941
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_938),
       .in0_consume_en(vin0_consume_en_941),
       .out_canPeek(vout_canPeek_941),
       .out_peek(vout_peek_941));
  assign v_942 = mux_942(v_943);
  assign v_943 = ~v_940;
  assign v_944 = v_945 | v_950;
  assign v_945 = mux_945(v_946);
  assign v_946 = v_947 & 1'h1;
  assign v_947 = v_948 & vout_canPeek_949;
  assign v_948 = ~vout_canPeek_941;
  pebbles_core
    pebbles_core_949
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_944),
       .in0_consume_en(vin0_consume_en_949),
       .out_canPeek(vout_canPeek_949),
       .out_peek(vout_peek_949));
  assign v_950 = mux_950(v_951);
  assign v_951 = ~v_946;
  assign v_952 = v_953 | v_956;
  assign v_953 = mux_953(v_954);
  assign v_954 = vout_canPeek_955 & 1'h1;
  pebbles_core
    pebbles_core_955
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_952),
       .in0_consume_en(vin0_consume_en_955),
       .out_canPeek(vout_canPeek_955),
       .out_peek(vout_peek_955));
  assign v_956 = mux_956(v_957);
  assign v_957 = ~v_954;
  assign v_958 = v_959 | v_964;
  assign v_959 = mux_959(v_960);
  assign v_960 = v_961 & 1'h1;
  assign v_961 = v_962 & vout_canPeek_963;
  assign v_962 = ~vout_canPeek_955;
  pebbles_core
    pebbles_core_963
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_958),
       .in0_consume_en(vin0_consume_en_963),
       .out_canPeek(vout_canPeek_963),
       .out_peek(vout_peek_963));
  assign v_964 = mux_964(v_965);
  assign v_965 = ~v_960;
  assign v_966 = v_967 | v_970;
  assign v_967 = mux_967(v_968);
  assign v_968 = vout_canPeek_969 & 1'h1;
  pebbles_core
    pebbles_core_969
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_966),
       .in0_consume_en(vin0_consume_en_969),
       .out_canPeek(vout_canPeek_969),
       .out_peek(vout_peek_969));
  assign v_970 = mux_970(v_971);
  assign v_971 = ~v_968;
  assign v_972 = v_973 | v_978;
  assign v_973 = mux_973(v_974);
  assign v_974 = v_975 & 1'h1;
  assign v_975 = v_976 & vout_canPeek_977;
  assign v_976 = ~vout_canPeek_969;
  pebbles_core
    pebbles_core_977
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_972),
       .in0_consume_en(vin0_consume_en_977),
       .out_canPeek(vout_canPeek_977),
       .out_peek(vout_peek_977));
  assign v_978 = mux_978(v_979);
  assign v_979 = ~v_974;
  assign v_980 = v_981 | v_984;
  assign v_981 = mux_981(v_982);
  assign v_982 = vout_canPeek_983 & 1'h1;
  pebbles_core
    pebbles_core_983
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_980),
       .in0_consume_en(vin0_consume_en_983),
       .out_canPeek(vout_canPeek_983),
       .out_peek(vout_peek_983));
  assign v_984 = mux_984(v_985);
  assign v_985 = ~v_982;
  assign v_986 = v_987 | v_992;
  assign v_987 = mux_987(v_988);
  assign v_988 = v_989 & 1'h1;
  assign v_989 = v_990 & vout_canPeek_991;
  assign v_990 = ~vout_canPeek_983;
  pebbles_core
    pebbles_core_991
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_986),
       .in0_consume_en(vin0_consume_en_991),
       .out_canPeek(vout_canPeek_991),
       .out_peek(vout_peek_991));
  assign v_992 = mux_992(v_993);
  assign v_993 = ~v_988;
  assign v_994 = v_995 | v_998;
  assign v_995 = mux_995(v_996);
  assign v_996 = vout_canPeek_997 & 1'h1;
  pebbles_core
    pebbles_core_997
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_994),
       .in0_consume_en(vin0_consume_en_997),
       .out_canPeek(vout_canPeek_997),
       .out_peek(vout_peek_997));
  assign v_998 = mux_998(v_999);
  assign v_999 = ~v_996;
  assign v_1000 = v_1001 | v_1006;
  assign v_1001 = mux_1001(v_1002);
  assign v_1002 = v_1003 & 1'h1;
  assign v_1003 = v_1004 & vout_canPeek_1005;
  assign v_1004 = ~vout_canPeek_997;
  pebbles_core
    pebbles_core_1005
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1000),
       .in0_consume_en(vin0_consume_en_1005),
       .out_canPeek(vout_canPeek_1005),
       .out_peek(vout_peek_1005));
  assign v_1006 = mux_1006(v_1007);
  assign v_1007 = ~v_1002;
  assign v_1008 = v_1009 | v_1012;
  assign v_1009 = mux_1009(v_1010);
  assign v_1010 = vout_canPeek_1011 & 1'h1;
  pebbles_core
    pebbles_core_1011
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1008),
       .in0_consume_en(vin0_consume_en_1011),
       .out_canPeek(vout_canPeek_1011),
       .out_peek(vout_peek_1011));
  assign v_1012 = mux_1012(v_1013);
  assign v_1013 = ~v_1010;
  assign v_1014 = v_1015 | v_1020;
  assign v_1015 = mux_1015(v_1016);
  assign v_1016 = v_1017 & 1'h1;
  assign v_1017 = v_1018 & vout_canPeek_1019;
  assign v_1018 = ~vout_canPeek_1011;
  pebbles_core
    pebbles_core_1019
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1014),
       .in0_consume_en(vin0_consume_en_1019),
       .out_canPeek(vout_canPeek_1019),
       .out_peek(vout_peek_1019));
  assign v_1020 = mux_1020(v_1021);
  assign v_1021 = ~v_1016;
  assign v_1022 = v_1023 | v_1026;
  assign v_1023 = mux_1023(v_1024);
  assign v_1024 = vout_canPeek_1025 & 1'h1;
  pebbles_core
    pebbles_core_1025
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1022),
       .in0_consume_en(vin0_consume_en_1025),
       .out_canPeek(vout_canPeek_1025),
       .out_peek(vout_peek_1025));
  assign v_1026 = mux_1026(v_1027);
  assign v_1027 = ~v_1024;
  assign v_1028 = v_1029 | v_1034;
  assign v_1029 = mux_1029(v_1030);
  assign v_1030 = v_1031 & 1'h1;
  assign v_1031 = v_1032 & vout_canPeek_1033;
  assign v_1032 = ~vout_canPeek_1025;
  pebbles_core
    pebbles_core_1033
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1028),
       .in0_consume_en(vin0_consume_en_1033),
       .out_canPeek(vout_canPeek_1033),
       .out_peek(vout_peek_1033));
  assign v_1034 = mux_1034(v_1035);
  assign v_1035 = ~v_1030;
  assign v_1036 = v_1037 | v_1040;
  assign v_1037 = mux_1037(v_1038);
  assign v_1038 = vout_canPeek_1039 & 1'h1;
  pebbles_core
    pebbles_core_1039
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1036),
       .in0_consume_en(vin0_consume_en_1039),
       .out_canPeek(vout_canPeek_1039),
       .out_peek(vout_peek_1039));
  assign v_1040 = mux_1040(v_1041);
  assign v_1041 = ~v_1038;
  assign v_1042 = v_1043 | v_1048;
  assign v_1043 = mux_1043(v_1044);
  assign v_1044 = v_1045 & 1'h1;
  assign v_1045 = v_1046 & vout_canPeek_1047;
  assign v_1046 = ~vout_canPeek_1039;
  pebbles_core
    pebbles_core_1047
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1042),
       .in0_consume_en(vin0_consume_en_1047),
       .out_canPeek(vout_canPeek_1047),
       .out_peek(vout_peek_1047));
  assign v_1048 = mux_1048(v_1049);
  assign v_1049 = ~v_1044;
  assign v_1050 = v_1051 | v_1054;
  assign v_1051 = mux_1051(v_1052);
  assign v_1052 = vout_canPeek_1053 & 1'h1;
  pebbles_core
    pebbles_core_1053
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1050),
       .in0_consume_en(vin0_consume_en_1053),
       .out_canPeek(vout_canPeek_1053),
       .out_peek(vout_peek_1053));
  assign v_1054 = mux_1054(v_1055);
  assign v_1055 = ~v_1052;
  assign v_1056 = v_1057 | v_1062;
  assign v_1057 = mux_1057(v_1058);
  assign v_1058 = v_1059 & 1'h1;
  assign v_1059 = v_1060 & vout_canPeek_1061;
  assign v_1060 = ~vout_canPeek_1053;
  pebbles_core
    pebbles_core_1061
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1056),
       .in0_consume_en(vin0_consume_en_1061),
       .out_canPeek(vout_canPeek_1061),
       .out_peek(vout_peek_1061));
  assign v_1062 = mux_1062(v_1063);
  assign v_1063 = ~v_1058;
  assign v_1064 = v_1065 | v_1068;
  assign v_1065 = mux_1065(v_1066);
  assign v_1066 = vout_canPeek_1067 & 1'h1;
  pebbles_core
    pebbles_core_1067
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1064),
       .in0_consume_en(vin0_consume_en_1067),
       .out_canPeek(vout_canPeek_1067),
       .out_peek(vout_peek_1067));
  assign v_1068 = mux_1068(v_1069);
  assign v_1069 = ~v_1066;
  assign v_1070 = v_1071 | v_1076;
  assign v_1071 = mux_1071(v_1072);
  assign v_1072 = v_1073 & 1'h1;
  assign v_1073 = v_1074 & vout_canPeek_1075;
  assign v_1074 = ~vout_canPeek_1067;
  pebbles_core
    pebbles_core_1075
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1070),
       .in0_consume_en(vin0_consume_en_1075),
       .out_canPeek(vout_canPeek_1075),
       .out_peek(vout_peek_1075));
  assign v_1076 = mux_1076(v_1077);
  assign v_1077 = ~v_1072;
  assign v_1078 = v_1079 | v_1082;
  assign v_1079 = mux_1079(v_1080);
  assign v_1080 = vout_canPeek_1081 & 1'h1;
  pebbles_core
    pebbles_core_1081
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1078),
       .in0_consume_en(vin0_consume_en_1081),
       .out_canPeek(vout_canPeek_1081),
       .out_peek(vout_peek_1081));
  assign v_1082 = mux_1082(v_1083);
  assign v_1083 = ~v_1080;
  assign v_1084 = v_1085 | v_1090;
  assign v_1085 = mux_1085(v_1086);
  assign v_1086 = v_1087 & 1'h1;
  assign v_1087 = v_1088 & vout_canPeek_1089;
  assign v_1088 = ~vout_canPeek_1081;
  pebbles_core
    pebbles_core_1089
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1084),
       .in0_consume_en(vin0_consume_en_1089),
       .out_canPeek(vout_canPeek_1089),
       .out_peek(vout_peek_1089));
  assign v_1090 = mux_1090(v_1091);
  assign v_1091 = ~v_1086;
  assign v_1092 = v_1093 | v_1096;
  assign v_1093 = mux_1093(v_1094);
  assign v_1094 = vout_canPeek_1095 & 1'h1;
  pebbles_core
    pebbles_core_1095
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1092),
       .in0_consume_en(vin0_consume_en_1095),
       .out_canPeek(vout_canPeek_1095),
       .out_peek(vout_peek_1095));
  assign v_1096 = mux_1096(v_1097);
  assign v_1097 = ~v_1094;
  assign v_1098 = v_1099 | v_1104;
  assign v_1099 = mux_1099(v_1100);
  assign v_1100 = v_1101 & 1'h1;
  assign v_1101 = v_1102 & vout_canPeek_1103;
  assign v_1102 = ~vout_canPeek_1095;
  pebbles_core
    pebbles_core_1103
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1098),
       .in0_consume_en(vin0_consume_en_1103),
       .out_canPeek(vout_canPeek_1103),
       .out_peek(vout_peek_1103));
  assign v_1104 = mux_1104(v_1105);
  assign v_1105 = ~v_1100;
  assign v_1106 = v_1107 | v_1110;
  assign v_1107 = mux_1107(v_1108);
  assign v_1108 = vout_canPeek_1109 & 1'h1;
  pebbles_core
    pebbles_core_1109
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1106),
       .in0_consume_en(vin0_consume_en_1109),
       .out_canPeek(vout_canPeek_1109),
       .out_peek(vout_peek_1109));
  assign v_1110 = mux_1110(v_1111);
  assign v_1111 = ~v_1108;
  assign v_1112 = v_1113 | v_1118;
  assign v_1113 = mux_1113(v_1114);
  assign v_1114 = v_1115 & 1'h1;
  assign v_1115 = v_1116 & vout_canPeek_1117;
  assign v_1116 = ~vout_canPeek_1109;
  pebbles_core
    pebbles_core_1117
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1112),
       .in0_consume_en(vin0_consume_en_1117),
       .out_canPeek(vout_canPeek_1117),
       .out_peek(vout_peek_1117));
  assign v_1118 = mux_1118(v_1119);
  assign v_1119 = ~v_1114;
  assign v_1120 = v_1121 | v_1124;
  assign v_1121 = mux_1121(v_1122);
  assign v_1122 = vout_canPeek_1123 & 1'h1;
  pebbles_core
    pebbles_core_1123
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1120),
       .in0_consume_en(vin0_consume_en_1123),
       .out_canPeek(vout_canPeek_1123),
       .out_peek(vout_peek_1123));
  assign v_1124 = mux_1124(v_1125);
  assign v_1125 = ~v_1122;
  assign v_1126 = v_1127 | v_1132;
  assign v_1127 = mux_1127(v_1128);
  assign v_1128 = v_1129 & 1'h1;
  assign v_1129 = v_1130 & vout_canPeek_1131;
  assign v_1130 = ~vout_canPeek_1123;
  pebbles_core
    pebbles_core_1131
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1126),
       .in0_consume_en(vin0_consume_en_1131),
       .out_canPeek(vout_canPeek_1131),
       .out_peek(vout_peek_1131));
  assign v_1132 = mux_1132(v_1133);
  assign v_1133 = ~v_1128;
  assign v_1134 = v_1135 | v_1138;
  assign v_1135 = mux_1135(v_1136);
  assign v_1136 = vout_canPeek_1137 & 1'h1;
  pebbles_core
    pebbles_core_1137
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1134),
       .in0_consume_en(vin0_consume_en_1137),
       .out_canPeek(vout_canPeek_1137),
       .out_peek(vout_peek_1137));
  assign v_1138 = mux_1138(v_1139);
  assign v_1139 = ~v_1136;
  assign v_1140 = v_1141 | v_1146;
  assign v_1141 = mux_1141(v_1142);
  assign v_1142 = v_1143 & 1'h1;
  assign v_1143 = v_1144 & vout_canPeek_1145;
  assign v_1144 = ~vout_canPeek_1137;
  pebbles_core
    pebbles_core_1145
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1140),
       .in0_consume_en(vin0_consume_en_1145),
       .out_canPeek(vout_canPeek_1145),
       .out_peek(vout_peek_1145));
  assign v_1146 = mux_1146(v_1147);
  assign v_1147 = ~v_1142;
  assign v_1148 = v_1149 | v_1152;
  assign v_1149 = mux_1149(v_1150);
  assign v_1150 = vout_canPeek_1151 & 1'h1;
  pebbles_core
    pebbles_core_1151
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1148),
       .in0_consume_en(vin0_consume_en_1151),
       .out_canPeek(vout_canPeek_1151),
       .out_peek(vout_peek_1151));
  assign v_1152 = mux_1152(v_1153);
  assign v_1153 = ~v_1150;
  assign v_1154 = v_1155 | v_1160;
  assign v_1155 = mux_1155(v_1156);
  assign v_1156 = v_1157 & 1'h1;
  assign v_1157 = v_1158 & vout_canPeek_1159;
  assign v_1158 = ~vout_canPeek_1151;
  pebbles_core
    pebbles_core_1159
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1154),
       .in0_consume_en(vin0_consume_en_1159),
       .out_canPeek(vout_canPeek_1159),
       .out_peek(vout_peek_1159));
  assign v_1160 = mux_1160(v_1161);
  assign v_1161 = ~v_1156;
  assign v_1162 = v_1163 | v_1166;
  assign v_1163 = mux_1163(v_1164);
  assign v_1164 = vout_canPeek_1165 & 1'h1;
  pebbles_core
    pebbles_core_1165
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1162),
       .in0_consume_en(vin0_consume_en_1165),
       .out_canPeek(vout_canPeek_1165),
       .out_peek(vout_peek_1165));
  assign v_1166 = mux_1166(v_1167);
  assign v_1167 = ~v_1164;
  assign v_1168 = v_1169 | v_1174;
  assign v_1169 = mux_1169(v_1170);
  assign v_1170 = v_1171 & 1'h1;
  assign v_1171 = v_1172 & vout_canPeek_1173;
  assign v_1172 = ~vout_canPeek_1165;
  pebbles_core
    pebbles_core_1173
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1168),
       .in0_consume_en(vin0_consume_en_1173),
       .out_canPeek(vout_canPeek_1173),
       .out_peek(vout_peek_1173));
  assign v_1174 = mux_1174(v_1175);
  assign v_1175 = ~v_1170;
  assign v_1176 = v_1177 | v_1180;
  assign v_1177 = mux_1177(v_1178);
  assign v_1178 = vout_canPeek_1179 & 1'h1;
  pebbles_core
    pebbles_core_1179
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1176),
       .in0_consume_en(vin0_consume_en_1179),
       .out_canPeek(vout_canPeek_1179),
       .out_peek(vout_peek_1179));
  assign v_1180 = mux_1180(v_1181);
  assign v_1181 = ~v_1178;
  assign v_1182 = v_1183 | v_1188;
  assign v_1183 = mux_1183(v_1184);
  assign v_1184 = v_1185 & 1'h1;
  assign v_1185 = v_1186 & vout_canPeek_1187;
  assign v_1186 = ~vout_canPeek_1179;
  pebbles_core
    pebbles_core_1187
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1182),
       .in0_consume_en(vin0_consume_en_1187),
       .out_canPeek(vout_canPeek_1187),
       .out_peek(vout_peek_1187));
  assign v_1188 = mux_1188(v_1189);
  assign v_1189 = ~v_1184;
  assign v_1190 = v_1191 | v_1194;
  assign v_1191 = mux_1191(v_1192);
  assign v_1192 = vout_canPeek_1193 & 1'h1;
  pebbles_core
    pebbles_core_1193
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1190),
       .in0_consume_en(vin0_consume_en_1193),
       .out_canPeek(vout_canPeek_1193),
       .out_peek(vout_peek_1193));
  assign v_1194 = mux_1194(v_1195);
  assign v_1195 = ~v_1192;
  assign v_1196 = v_1197 | v_1202;
  assign v_1197 = mux_1197(v_1198);
  assign v_1198 = v_1199 & 1'h1;
  assign v_1199 = v_1200 & vout_canPeek_1201;
  assign v_1200 = ~vout_canPeek_1193;
  pebbles_core
    pebbles_core_1201
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1196),
       .in0_consume_en(vin0_consume_en_1201),
       .out_canPeek(vout_canPeek_1201),
       .out_peek(vout_peek_1201));
  assign v_1202 = mux_1202(v_1203);
  assign v_1203 = ~v_1198;
  assign v_1204 = v_1205 | v_1208;
  assign v_1205 = mux_1205(v_1206);
  assign v_1206 = vout_canPeek_1207 & 1'h1;
  pebbles_core
    pebbles_core_1207
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1204),
       .in0_consume_en(vin0_consume_en_1207),
       .out_canPeek(vout_canPeek_1207),
       .out_peek(vout_peek_1207));
  assign v_1208 = mux_1208(v_1209);
  assign v_1209 = ~v_1206;
  assign v_1210 = v_1211 | v_1216;
  assign v_1211 = mux_1211(v_1212);
  assign v_1212 = v_1213 & 1'h1;
  assign v_1213 = v_1214 & vout_canPeek_1215;
  assign v_1214 = ~vout_canPeek_1207;
  pebbles_core
    pebbles_core_1215
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1210),
       .in0_consume_en(vin0_consume_en_1215),
       .out_canPeek(vout_canPeek_1215),
       .out_peek(vout_peek_1215));
  assign v_1216 = mux_1216(v_1217);
  assign v_1217 = ~v_1212;
  assign v_1218 = v_1219 | v_1222;
  assign v_1219 = mux_1219(v_1220);
  assign v_1220 = vout_canPeek_1221 & 1'h1;
  pebbles_core
    pebbles_core_1221
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1218),
       .in0_consume_en(vin0_consume_en_1221),
       .out_canPeek(vout_canPeek_1221),
       .out_peek(vout_peek_1221));
  assign v_1222 = mux_1222(v_1223);
  assign v_1223 = ~v_1220;
  assign v_1224 = v_1225 | v_1230;
  assign v_1225 = mux_1225(v_1226);
  assign v_1226 = v_1227 & 1'h1;
  assign v_1227 = v_1228 & vout_canPeek_1229;
  assign v_1228 = ~vout_canPeek_1221;
  pebbles_core
    pebbles_core_1229
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1224),
       .in0_consume_en(vin0_consume_en_1229),
       .out_canPeek(vout_canPeek_1229),
       .out_peek(vout_peek_1229));
  assign v_1230 = mux_1230(v_1231);
  assign v_1231 = ~v_1226;
  assign v_1232 = v_1233 | v_1236;
  assign v_1233 = mux_1233(v_1234);
  assign v_1234 = vout_canPeek_1235 & 1'h1;
  pebbles_core
    pebbles_core_1235
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1232),
       .in0_consume_en(vin0_consume_en_1235),
       .out_canPeek(vout_canPeek_1235),
       .out_peek(vout_peek_1235));
  assign v_1236 = mux_1236(v_1237);
  assign v_1237 = ~v_1234;
  assign v_1238 = v_1239 | v_1244;
  assign v_1239 = mux_1239(v_1240);
  assign v_1240 = v_1241 & 1'h1;
  assign v_1241 = v_1242 & vout_canPeek_1243;
  assign v_1242 = ~vout_canPeek_1235;
  pebbles_core
    pebbles_core_1243
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1238),
       .in0_consume_en(vin0_consume_en_1243),
       .out_canPeek(vout_canPeek_1243),
       .out_peek(vout_peek_1243));
  assign v_1244 = mux_1244(v_1245);
  assign v_1245 = ~v_1240;
  assign v_1246 = v_1247 | v_1250;
  assign v_1247 = mux_1247(v_1248);
  assign v_1248 = vout_canPeek_1249 & 1'h1;
  pebbles_core
    pebbles_core_1249
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1246),
       .in0_consume_en(vin0_consume_en_1249),
       .out_canPeek(vout_canPeek_1249),
       .out_peek(vout_peek_1249));
  assign v_1250 = mux_1250(v_1251);
  assign v_1251 = ~v_1248;
  assign v_1252 = v_1253 | v_1258;
  assign v_1253 = mux_1253(v_1254);
  assign v_1254 = v_1255 & 1'h1;
  assign v_1255 = v_1256 & vout_canPeek_1257;
  assign v_1256 = ~vout_canPeek_1249;
  pebbles_core
    pebbles_core_1257
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1252),
       .in0_consume_en(vin0_consume_en_1257),
       .out_canPeek(vout_canPeek_1257),
       .out_peek(vout_peek_1257));
  assign v_1258 = mux_1258(v_1259);
  assign v_1259 = ~v_1254;
  assign v_1260 = v_1261 | v_1264;
  assign v_1261 = mux_1261(v_1262);
  assign v_1262 = vout_canPeek_1263 & 1'h1;
  pebbles_core
    pebbles_core_1263
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1260),
       .in0_consume_en(vin0_consume_en_1263),
       .out_canPeek(vout_canPeek_1263),
       .out_peek(vout_peek_1263));
  assign v_1264 = mux_1264(v_1265);
  assign v_1265 = ~v_1262;
  assign v_1266 = v_1267 | v_1272;
  assign v_1267 = mux_1267(v_1268);
  assign v_1268 = v_1269 & 1'h1;
  assign v_1269 = v_1270 & vout_canPeek_1271;
  assign v_1270 = ~vout_canPeek_1263;
  pebbles_core
    pebbles_core_1271
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1266),
       .in0_consume_en(vin0_consume_en_1271),
       .out_canPeek(vout_canPeek_1271),
       .out_peek(vout_peek_1271));
  assign v_1272 = mux_1272(v_1273);
  assign v_1273 = ~v_1268;
  assign v_1274 = v_1275 | v_1278;
  assign v_1275 = mux_1275(v_1276);
  assign v_1276 = vout_canPeek_1277 & 1'h1;
  pebbles_core
    pebbles_core_1277
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1274),
       .in0_consume_en(vin0_consume_en_1277),
       .out_canPeek(vout_canPeek_1277),
       .out_peek(vout_peek_1277));
  assign v_1278 = mux_1278(v_1279);
  assign v_1279 = ~v_1276;
  assign v_1280 = v_1281 | v_1286;
  assign v_1281 = mux_1281(v_1282);
  assign v_1282 = v_1283 & 1'h1;
  assign v_1283 = v_1284 & vout_canPeek_1285;
  assign v_1284 = ~vout_canPeek_1277;
  pebbles_core
    pebbles_core_1285
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1280),
       .in0_consume_en(vin0_consume_en_1285),
       .out_canPeek(vout_canPeek_1285),
       .out_peek(vout_peek_1285));
  assign v_1286 = mux_1286(v_1287);
  assign v_1287 = ~v_1282;
  assign v_1288 = v_1289 | v_1292;
  assign v_1289 = mux_1289(v_1290);
  assign v_1290 = vout_canPeek_1291 & 1'h1;
  pebbles_core
    pebbles_core_1291
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1288),
       .in0_consume_en(vin0_consume_en_1291),
       .out_canPeek(vout_canPeek_1291),
       .out_peek(vout_peek_1291));
  assign v_1292 = mux_1292(v_1293);
  assign v_1293 = ~v_1290;
  assign v_1294 = v_1295 | v_1300;
  assign v_1295 = mux_1295(v_1296);
  assign v_1296 = v_1297 & 1'h1;
  assign v_1297 = v_1298 & vout_canPeek_1299;
  assign v_1298 = ~vout_canPeek_1291;
  pebbles_core
    pebbles_core_1299
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1294),
       .in0_consume_en(vin0_consume_en_1299),
       .out_canPeek(vout_canPeek_1299),
       .out_peek(vout_peek_1299));
  assign v_1300 = mux_1300(v_1301);
  assign v_1301 = ~v_1296;
  assign v_1302 = v_1303 | v_1306;
  assign v_1303 = mux_1303(v_1304);
  assign v_1304 = vout_canPeek_1305 & 1'h1;
  pebbles_core
    pebbles_core_1305
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1302),
       .in0_consume_en(vin0_consume_en_1305),
       .out_canPeek(vout_canPeek_1305),
       .out_peek(vout_peek_1305));
  assign v_1306 = mux_1306(v_1307);
  assign v_1307 = ~v_1304;
  assign v_1308 = v_1309 | v_1314;
  assign v_1309 = mux_1309(v_1310);
  assign v_1310 = v_1311 & 1'h1;
  assign v_1311 = v_1312 & vout_canPeek_1313;
  assign v_1312 = ~vout_canPeek_1305;
  pebbles_core
    pebbles_core_1313
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1308),
       .in0_consume_en(vin0_consume_en_1313),
       .out_canPeek(vout_canPeek_1313),
       .out_peek(vout_peek_1313));
  assign v_1314 = mux_1314(v_1315);
  assign v_1315 = ~v_1310;
  assign v_1316 = v_1317 | v_1320;
  assign v_1317 = mux_1317(v_1318);
  assign v_1318 = vout_canPeek_1319 & 1'h1;
  pebbles_core
    pebbles_core_1319
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1316),
       .in0_consume_en(vin0_consume_en_1319),
       .out_canPeek(vout_canPeek_1319),
       .out_peek(vout_peek_1319));
  assign v_1320 = mux_1320(v_1321);
  assign v_1321 = ~v_1318;
  assign v_1322 = v_1323 | v_1328;
  assign v_1323 = mux_1323(v_1324);
  assign v_1324 = v_1325 & 1'h1;
  assign v_1325 = v_1326 & vout_canPeek_1327;
  assign v_1326 = ~vout_canPeek_1319;
  pebbles_core
    pebbles_core_1327
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1322),
       .in0_consume_en(vin0_consume_en_1327),
       .out_canPeek(vout_canPeek_1327),
       .out_peek(vout_peek_1327));
  assign v_1328 = mux_1328(v_1329);
  assign v_1329 = ~v_1324;
  assign v_1330 = v_1331 | v_1334;
  assign v_1331 = mux_1331(v_1332);
  assign v_1332 = vout_canPeek_1333 & 1'h1;
  pebbles_core
    pebbles_core_1333
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1330),
       .in0_consume_en(vin0_consume_en_1333),
       .out_canPeek(vout_canPeek_1333),
       .out_peek(vout_peek_1333));
  assign v_1334 = mux_1334(v_1335);
  assign v_1335 = ~v_1332;
  assign v_1336 = v_1337 | v_1342;
  assign v_1337 = mux_1337(v_1338);
  assign v_1338 = v_1339 & 1'h1;
  assign v_1339 = v_1340 & vout_canPeek_1341;
  assign v_1340 = ~vout_canPeek_1333;
  pebbles_core
    pebbles_core_1341
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1336),
       .in0_consume_en(vin0_consume_en_1341),
       .out_canPeek(vout_canPeek_1341),
       .out_peek(vout_peek_1341));
  assign v_1342 = mux_1342(v_1343);
  assign v_1343 = ~v_1338;
  assign v_1344 = v_1345 | v_1348;
  assign v_1345 = mux_1345(v_1346);
  assign v_1346 = vout_canPeek_1347 & 1'h1;
  pebbles_core
    pebbles_core_1347
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1344),
       .in0_consume_en(vin0_consume_en_1347),
       .out_canPeek(vout_canPeek_1347),
       .out_peek(vout_peek_1347));
  assign v_1348 = mux_1348(v_1349);
  assign v_1349 = ~v_1346;
  assign v_1350 = v_1351 | v_1356;
  assign v_1351 = mux_1351(v_1352);
  assign v_1352 = v_1353 & 1'h1;
  assign v_1353 = v_1354 & vout_canPeek_1355;
  assign v_1354 = ~vout_canPeek_1347;
  pebbles_core
    pebbles_core_1355
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1350),
       .in0_consume_en(vin0_consume_en_1355),
       .out_canPeek(vout_canPeek_1355),
       .out_peek(vout_peek_1355));
  assign v_1356 = mux_1356(v_1357);
  assign v_1357 = ~v_1352;
  assign v_1358 = v_1359 | v_1362;
  assign v_1359 = mux_1359(v_1360);
  assign v_1360 = vout_canPeek_1361 & 1'h1;
  pebbles_core
    pebbles_core_1361
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1358),
       .in0_consume_en(vin0_consume_en_1361),
       .out_canPeek(vout_canPeek_1361),
       .out_peek(vout_peek_1361));
  assign v_1362 = mux_1362(v_1363);
  assign v_1363 = ~v_1360;
  assign v_1364 = v_1365 | v_1370;
  assign v_1365 = mux_1365(v_1366);
  assign v_1366 = v_1367 & 1'h1;
  assign v_1367 = v_1368 & vout_canPeek_1369;
  assign v_1368 = ~vout_canPeek_1361;
  pebbles_core
    pebbles_core_1369
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1364),
       .in0_consume_en(vin0_consume_en_1369),
       .out_canPeek(vout_canPeek_1369),
       .out_peek(vout_peek_1369));
  assign v_1370 = mux_1370(v_1371);
  assign v_1371 = ~v_1366;
  assign v_1372 = v_1373 | v_1376;
  assign v_1373 = mux_1373(v_1374);
  assign v_1374 = vout_canPeek_1375 & 1'h1;
  pebbles_core
    pebbles_core_1375
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1372),
       .in0_consume_en(vin0_consume_en_1375),
       .out_canPeek(vout_canPeek_1375),
       .out_peek(vout_peek_1375));
  assign v_1376 = mux_1376(v_1377);
  assign v_1377 = ~v_1374;
  assign v_1378 = v_1379 | v_1384;
  assign v_1379 = mux_1379(v_1380);
  assign v_1380 = v_1381 & 1'h1;
  assign v_1381 = v_1382 & vout_canPeek_1383;
  assign v_1382 = ~vout_canPeek_1375;
  pebbles_core
    pebbles_core_1383
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1378),
       .in0_consume_en(vin0_consume_en_1383),
       .out_canPeek(vout_canPeek_1383),
       .out_peek(vout_peek_1383));
  assign v_1384 = mux_1384(v_1385);
  assign v_1385 = ~v_1380;
  assign v_1386 = v_1387 | v_1390;
  assign v_1387 = mux_1387(v_1388);
  assign v_1388 = vout_canPeek_1389 & 1'h1;
  pebbles_core
    pebbles_core_1389
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1386),
       .in0_consume_en(vin0_consume_en_1389),
       .out_canPeek(vout_canPeek_1389),
       .out_peek(vout_peek_1389));
  assign v_1390 = mux_1390(v_1391);
  assign v_1391 = ~v_1388;
  assign v_1392 = v_1393 | v_1398;
  assign v_1393 = mux_1393(v_1394);
  assign v_1394 = v_1395 & 1'h1;
  assign v_1395 = v_1396 & vout_canPeek_1397;
  assign v_1396 = ~vout_canPeek_1389;
  pebbles_core
    pebbles_core_1397
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1392),
       .in0_consume_en(vin0_consume_en_1397),
       .out_canPeek(vout_canPeek_1397),
       .out_peek(vout_peek_1397));
  assign v_1398 = mux_1398(v_1399);
  assign v_1399 = ~v_1394;
  assign v_1400 = v_1401 | v_1404;
  assign v_1401 = mux_1401(v_1402);
  assign v_1402 = vout_canPeek_1403 & 1'h1;
  pebbles_core
    pebbles_core_1403
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1400),
       .in0_consume_en(vin0_consume_en_1403),
       .out_canPeek(vout_canPeek_1403),
       .out_peek(vout_peek_1403));
  assign v_1404 = mux_1404(v_1405);
  assign v_1405 = ~v_1402;
  assign v_1406 = v_1407 | v_1412;
  assign v_1407 = mux_1407(v_1408);
  assign v_1408 = v_1409 & 1'h1;
  assign v_1409 = v_1410 & vout_canPeek_1411;
  assign v_1410 = ~vout_canPeek_1403;
  pebbles_core
    pebbles_core_1411
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1406),
       .in0_consume_en(vin0_consume_en_1411),
       .out_canPeek(vout_canPeek_1411),
       .out_peek(vout_peek_1411));
  assign v_1412 = mux_1412(v_1413);
  assign v_1413 = ~v_1408;
  assign v_1414 = v_1415 | v_1418;
  assign v_1415 = mux_1415(v_1416);
  assign v_1416 = vout_canPeek_1417 & 1'h1;
  pebbles_core
    pebbles_core_1417
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1414),
       .in0_consume_en(vin0_consume_en_1417),
       .out_canPeek(vout_canPeek_1417),
       .out_peek(vout_peek_1417));
  assign v_1418 = mux_1418(v_1419);
  assign v_1419 = ~v_1416;
  assign v_1420 = v_1421 | v_1426;
  assign v_1421 = mux_1421(v_1422);
  assign v_1422 = v_1423 & 1'h1;
  assign v_1423 = v_1424 & vout_canPeek_1425;
  assign v_1424 = ~vout_canPeek_1417;
  pebbles_core
    pebbles_core_1425
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1420),
       .in0_consume_en(vin0_consume_en_1425),
       .out_canPeek(vout_canPeek_1425),
       .out_peek(vout_peek_1425));
  assign v_1426 = mux_1426(v_1427);
  assign v_1427 = ~v_1422;
  assign v_1428 = v_1429 | v_1432;
  assign v_1429 = mux_1429(v_1430);
  assign v_1430 = vout_canPeek_1431 & 1'h1;
  pebbles_core
    pebbles_core_1431
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1428),
       .in0_consume_en(vin0_consume_en_1431),
       .out_canPeek(vout_canPeek_1431),
       .out_peek(vout_peek_1431));
  assign v_1432 = mux_1432(v_1433);
  assign v_1433 = ~v_1430;
  assign v_1434 = v_1435 | v_1440;
  assign v_1435 = mux_1435(v_1436);
  assign v_1436 = v_1437 & 1'h1;
  assign v_1437 = v_1438 & vout_canPeek_1439;
  assign v_1438 = ~vout_canPeek_1431;
  pebbles_core
    pebbles_core_1439
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1434),
       .in0_consume_en(vin0_consume_en_1439),
       .out_canPeek(vout_canPeek_1439),
       .out_peek(vout_peek_1439));
  assign v_1440 = mux_1440(v_1441);
  assign v_1441 = ~v_1436;
  assign v_1442 = v_1443 | v_1446;
  assign v_1443 = mux_1443(v_1444);
  assign v_1444 = vout_canPeek_1445 & 1'h1;
  pebbles_core
    pebbles_core_1445
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1442),
       .in0_consume_en(vin0_consume_en_1445),
       .out_canPeek(vout_canPeek_1445),
       .out_peek(vout_peek_1445));
  assign v_1446 = mux_1446(v_1447);
  assign v_1447 = ~v_1444;
  assign v_1448 = v_1449 | v_1454;
  assign v_1449 = mux_1449(v_1450);
  assign v_1450 = v_1451 & 1'h1;
  assign v_1451 = v_1452 & vout_canPeek_1453;
  assign v_1452 = ~vout_canPeek_1445;
  pebbles_core
    pebbles_core_1453
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1448),
       .in0_consume_en(vin0_consume_en_1453),
       .out_canPeek(vout_canPeek_1453),
       .out_peek(vout_peek_1453));
  assign v_1454 = mux_1454(v_1455);
  assign v_1455 = ~v_1450;
  assign v_1456 = v_1457 | v_1460;
  assign v_1457 = mux_1457(v_1458);
  assign v_1458 = vout_canPeek_1459 & 1'h1;
  pebbles_core
    pebbles_core_1459
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1456),
       .in0_consume_en(vin0_consume_en_1459),
       .out_canPeek(vout_canPeek_1459),
       .out_peek(vout_peek_1459));
  assign v_1460 = mux_1460(v_1461);
  assign v_1461 = ~v_1458;
  assign v_1462 = v_1463 | v_1468;
  assign v_1463 = mux_1463(v_1464);
  assign v_1464 = v_1465 & 1'h1;
  assign v_1465 = v_1466 & vout_canPeek_1467;
  assign v_1466 = ~vout_canPeek_1459;
  pebbles_core
    pebbles_core_1467
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1462),
       .in0_consume_en(vin0_consume_en_1467),
       .out_canPeek(vout_canPeek_1467),
       .out_peek(vout_peek_1467));
  assign v_1468 = mux_1468(v_1469);
  assign v_1469 = ~v_1464;
  assign v_1470 = v_1471 | v_1474;
  assign v_1471 = mux_1471(v_1472);
  assign v_1472 = vout_canPeek_1473 & 1'h1;
  pebbles_core
    pebbles_core_1473
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1470),
       .in0_consume_en(vin0_consume_en_1473),
       .out_canPeek(vout_canPeek_1473),
       .out_peek(vout_peek_1473));
  assign v_1474 = mux_1474(v_1475);
  assign v_1475 = ~v_1472;
  assign v_1476 = v_1477 | v_1482;
  assign v_1477 = mux_1477(v_1478);
  assign v_1478 = v_1479 & 1'h1;
  assign v_1479 = v_1480 & vout_canPeek_1481;
  assign v_1480 = ~vout_canPeek_1473;
  pebbles_core
    pebbles_core_1481
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1476),
       .in0_consume_en(vin0_consume_en_1481),
       .out_canPeek(vout_canPeek_1481),
       .out_peek(vout_peek_1481));
  assign v_1482 = mux_1482(v_1483);
  assign v_1483 = ~v_1478;
  assign v_1484 = v_1485 | v_1488;
  assign v_1485 = mux_1485(v_1486);
  assign v_1486 = vout_canPeek_1487 & 1'h1;
  pebbles_core
    pebbles_core_1487
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1484),
       .in0_consume_en(vin0_consume_en_1487),
       .out_canPeek(vout_canPeek_1487),
       .out_peek(vout_peek_1487));
  assign v_1488 = mux_1488(v_1489);
  assign v_1489 = ~v_1486;
  assign v_1490 = v_1491 | v_1496;
  assign v_1491 = mux_1491(v_1492);
  assign v_1492 = v_1493 & 1'h1;
  assign v_1493 = v_1494 & vout_canPeek_1495;
  assign v_1494 = ~vout_canPeek_1487;
  pebbles_core
    pebbles_core_1495
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1490),
       .in0_consume_en(vin0_consume_en_1495),
       .out_canPeek(vout_canPeek_1495),
       .out_peek(vout_peek_1495));
  assign v_1496 = mux_1496(v_1497);
  assign v_1497 = ~v_1492;
  assign v_1498 = v_1499 | v_1502;
  assign v_1499 = mux_1499(v_1500);
  assign v_1500 = vout_canPeek_1501 & 1'h1;
  pebbles_core
    pebbles_core_1501
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1498),
       .in0_consume_en(vin0_consume_en_1501),
       .out_canPeek(vout_canPeek_1501),
       .out_peek(vout_peek_1501));
  assign v_1502 = mux_1502(v_1503);
  assign v_1503 = ~v_1500;
  assign v_1504 = v_1505 | v_1510;
  assign v_1505 = mux_1505(v_1506);
  assign v_1506 = v_1507 & 1'h1;
  assign v_1507 = v_1508 & vout_canPeek_1509;
  assign v_1508 = ~vout_canPeek_1501;
  pebbles_core
    pebbles_core_1509
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1504),
       .in0_consume_en(vin0_consume_en_1509),
       .out_canPeek(vout_canPeek_1509),
       .out_peek(vout_peek_1509));
  assign v_1510 = mux_1510(v_1511);
  assign v_1511 = ~v_1506;
  assign v_1512 = v_1513 | v_1516;
  assign v_1513 = mux_1513(v_1514);
  assign v_1514 = vout_canPeek_1515 & 1'h1;
  pebbles_core
    pebbles_core_1515
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1512),
       .in0_consume_en(vin0_consume_en_1515),
       .out_canPeek(vout_canPeek_1515),
       .out_peek(vout_peek_1515));
  assign v_1516 = mux_1516(v_1517);
  assign v_1517 = ~v_1514;
  assign v_1518 = v_1519 | v_1524;
  assign v_1519 = mux_1519(v_1520);
  assign v_1520 = v_1521 & 1'h1;
  assign v_1521 = v_1522 & vout_canPeek_1523;
  assign v_1522 = ~vout_canPeek_1515;
  pebbles_core
    pebbles_core_1523
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1518),
       .in0_consume_en(vin0_consume_en_1523),
       .out_canPeek(vout_canPeek_1523),
       .out_peek(vout_peek_1523));
  assign v_1524 = mux_1524(v_1525);
  assign v_1525 = ~v_1520;
  assign v_1526 = v_1527 | v_1530;
  assign v_1527 = mux_1527(v_1528);
  assign v_1528 = vout_canPeek_1529 & 1'h1;
  pebbles_core
    pebbles_core_1529
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1526),
       .in0_consume_en(vin0_consume_en_1529),
       .out_canPeek(vout_canPeek_1529),
       .out_peek(vout_peek_1529));
  assign v_1530 = mux_1530(v_1531);
  assign v_1531 = ~v_1528;
  assign v_1532 = v_1533 | v_1538;
  assign v_1533 = mux_1533(v_1534);
  assign v_1534 = v_1535 & 1'h1;
  assign v_1535 = v_1536 & vout_canPeek_1537;
  assign v_1536 = ~vout_canPeek_1529;
  pebbles_core
    pebbles_core_1537
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1532),
       .in0_consume_en(vin0_consume_en_1537),
       .out_canPeek(vout_canPeek_1537),
       .out_peek(vout_peek_1537));
  assign v_1538 = mux_1538(v_1539);
  assign v_1539 = ~v_1534;
  assign v_1540 = v_1541 | v_1544;
  assign v_1541 = mux_1541(v_1542);
  assign v_1542 = vout_canPeek_1543 & 1'h1;
  pebbles_core
    pebbles_core_1543
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1540),
       .in0_consume_en(vin0_consume_en_1543),
       .out_canPeek(vout_canPeek_1543),
       .out_peek(vout_peek_1543));
  assign v_1544 = mux_1544(v_1545);
  assign v_1545 = ~v_1542;
  assign v_1546 = v_1547 | v_1552;
  assign v_1547 = mux_1547(v_1548);
  assign v_1548 = v_1549 & 1'h1;
  assign v_1549 = v_1550 & vout_canPeek_1551;
  assign v_1550 = ~vout_canPeek_1543;
  pebbles_core
    pebbles_core_1551
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1546),
       .in0_consume_en(vin0_consume_en_1551),
       .out_canPeek(vout_canPeek_1551),
       .out_peek(vout_peek_1551));
  assign v_1552 = mux_1552(v_1553);
  assign v_1553 = ~v_1548;
  assign v_1554 = v_1555 | v_1558;
  assign v_1555 = mux_1555(v_1556);
  assign v_1556 = vout_canPeek_1557 & 1'h1;
  pebbles_core
    pebbles_core_1557
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1554),
       .in0_consume_en(vin0_consume_en_1557),
       .out_canPeek(vout_canPeek_1557),
       .out_peek(vout_peek_1557));
  assign v_1558 = mux_1558(v_1559);
  assign v_1559 = ~v_1556;
  assign v_1560 = v_1561 | v_1566;
  assign v_1561 = mux_1561(v_1562);
  assign v_1562 = v_1563 & 1'h1;
  assign v_1563 = v_1564 & vout_canPeek_1565;
  assign v_1564 = ~vout_canPeek_1557;
  pebbles_core
    pebbles_core_1565
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1560),
       .in0_consume_en(vin0_consume_en_1565),
       .out_canPeek(vout_canPeek_1565),
       .out_peek(vout_peek_1565));
  assign v_1566 = mux_1566(v_1567);
  assign v_1567 = ~v_1562;
  assign v_1568 = v_1569 | v_1572;
  assign v_1569 = mux_1569(v_1570);
  assign v_1570 = vout_canPeek_1571 & 1'h1;
  pebbles_core
    pebbles_core_1571
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1568),
       .in0_consume_en(vin0_consume_en_1571),
       .out_canPeek(vout_canPeek_1571),
       .out_peek(vout_peek_1571));
  assign v_1572 = mux_1572(v_1573);
  assign v_1573 = ~v_1570;
  assign v_1574 = v_1575 | v_1580;
  assign v_1575 = mux_1575(v_1576);
  assign v_1576 = v_1577 & 1'h1;
  assign v_1577 = v_1578 & vout_canPeek_1579;
  assign v_1578 = ~vout_canPeek_1571;
  pebbles_core
    pebbles_core_1579
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1574),
       .in0_consume_en(vin0_consume_en_1579),
       .out_canPeek(vout_canPeek_1579),
       .out_peek(vout_peek_1579));
  assign v_1580 = mux_1580(v_1581);
  assign v_1581 = ~v_1576;
  assign v_1582 = v_1583 | v_1586;
  assign v_1583 = mux_1583(v_1584);
  assign v_1584 = vout_canPeek_1585 & 1'h1;
  pebbles_core
    pebbles_core_1585
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1582),
       .in0_consume_en(vin0_consume_en_1585),
       .out_canPeek(vout_canPeek_1585),
       .out_peek(vout_peek_1585));
  assign v_1586 = mux_1586(v_1587);
  assign v_1587 = ~v_1584;
  assign v_1588 = v_1589 | v_1594;
  assign v_1589 = mux_1589(v_1590);
  assign v_1590 = v_1591 & 1'h1;
  assign v_1591 = v_1592 & vout_canPeek_1593;
  assign v_1592 = ~vout_canPeek_1585;
  pebbles_core
    pebbles_core_1593
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1588),
       .in0_consume_en(vin0_consume_en_1593),
       .out_canPeek(vout_canPeek_1593),
       .out_peek(vout_peek_1593));
  assign v_1594 = mux_1594(v_1595);
  assign v_1595 = ~v_1590;
  assign v_1596 = v_1597 | v_1600;
  assign v_1597 = mux_1597(v_1598);
  assign v_1598 = vout_canPeek_1599 & 1'h1;
  pebbles_core
    pebbles_core_1599
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1596),
       .in0_consume_en(vin0_consume_en_1599),
       .out_canPeek(vout_canPeek_1599),
       .out_peek(vout_peek_1599));
  assign v_1600 = mux_1600(v_1601);
  assign v_1601 = ~v_1598;
  assign v_1602 = v_1603 | v_1608;
  assign v_1603 = mux_1603(v_1604);
  assign v_1604 = v_1605 & 1'h1;
  assign v_1605 = v_1606 & vout_canPeek_1607;
  assign v_1606 = ~vout_canPeek_1599;
  pebbles_core
    pebbles_core_1607
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1602),
       .in0_consume_en(vin0_consume_en_1607),
       .out_canPeek(vout_canPeek_1607),
       .out_peek(vout_peek_1607));
  assign v_1608 = mux_1608(v_1609);
  assign v_1609 = ~v_1604;
  assign v_1610 = v_1611 | v_1614;
  assign v_1611 = mux_1611(v_1612);
  assign v_1612 = vout_canPeek_1613 & 1'h1;
  pebbles_core
    pebbles_core_1613
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1610),
       .in0_consume_en(vin0_consume_en_1613),
       .out_canPeek(vout_canPeek_1613),
       .out_peek(vout_peek_1613));
  assign v_1614 = mux_1614(v_1615);
  assign v_1615 = ~v_1612;
  assign v_1616 = v_1617 | v_1622;
  assign v_1617 = mux_1617(v_1618);
  assign v_1618 = v_1619 & 1'h1;
  assign v_1619 = v_1620 & vout_canPeek_1621;
  assign v_1620 = ~vout_canPeek_1613;
  pebbles_core
    pebbles_core_1621
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1616),
       .in0_consume_en(vin0_consume_en_1621),
       .out_canPeek(vout_canPeek_1621),
       .out_peek(vout_peek_1621));
  assign v_1622 = mux_1622(v_1623);
  assign v_1623 = ~v_1618;
  assign v_1624 = v_1625 | v_1628;
  assign v_1625 = mux_1625(v_1626);
  assign v_1626 = vout_canPeek_1627 & 1'h1;
  pebbles_core
    pebbles_core_1627
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1624),
       .in0_consume_en(vin0_consume_en_1627),
       .out_canPeek(vout_canPeek_1627),
       .out_peek(vout_peek_1627));
  assign v_1628 = mux_1628(v_1629);
  assign v_1629 = ~v_1626;
  assign v_1630 = v_1631 | v_1636;
  assign v_1631 = mux_1631(v_1632);
  assign v_1632 = v_1633 & 1'h1;
  assign v_1633 = v_1634 & vout_canPeek_1635;
  assign v_1634 = ~vout_canPeek_1627;
  pebbles_core
    pebbles_core_1635
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1630),
       .in0_consume_en(vin0_consume_en_1635),
       .out_canPeek(vout_canPeek_1635),
       .out_peek(vout_peek_1635));
  assign v_1636 = mux_1636(v_1637);
  assign v_1637 = ~v_1632;
  assign v_1638 = v_1639 | v_1642;
  assign v_1639 = mux_1639(v_1640);
  assign v_1640 = vout_canPeek_1641 & 1'h1;
  pebbles_core
    pebbles_core_1641
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1638),
       .in0_consume_en(vin0_consume_en_1641),
       .out_canPeek(vout_canPeek_1641),
       .out_peek(vout_peek_1641));
  assign v_1642 = mux_1642(v_1643);
  assign v_1643 = ~v_1640;
  assign v_1644 = v_1645 | v_1650;
  assign v_1645 = mux_1645(v_1646);
  assign v_1646 = v_1647 & 1'h1;
  assign v_1647 = v_1648 & vout_canPeek_1649;
  assign v_1648 = ~vout_canPeek_1641;
  pebbles_core
    pebbles_core_1649
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1644),
       .in0_consume_en(vin0_consume_en_1649),
       .out_canPeek(vout_canPeek_1649),
       .out_peek(vout_peek_1649));
  assign v_1650 = mux_1650(v_1651);
  assign v_1651 = ~v_1646;
  assign v_1652 = v_1653 | v_1656;
  assign v_1653 = mux_1653(v_1654);
  assign v_1654 = vout_canPeek_1655 & 1'h1;
  pebbles_core
    pebbles_core_1655
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1652),
       .in0_consume_en(vin0_consume_en_1655),
       .out_canPeek(vout_canPeek_1655),
       .out_peek(vout_peek_1655));
  assign v_1656 = mux_1656(v_1657);
  assign v_1657 = ~v_1654;
  assign v_1658 = v_1659 | v_1664;
  assign v_1659 = mux_1659(v_1660);
  assign v_1660 = v_1661 & 1'h1;
  assign v_1661 = v_1662 & vout_canPeek_1663;
  assign v_1662 = ~vout_canPeek_1655;
  pebbles_core
    pebbles_core_1663
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1658),
       .in0_consume_en(vin0_consume_en_1663),
       .out_canPeek(vout_canPeek_1663),
       .out_peek(vout_peek_1663));
  assign v_1664 = mux_1664(v_1665);
  assign v_1665 = ~v_1660;
  assign v_1666 = v_1667 | v_1670;
  assign v_1667 = mux_1667(v_1668);
  assign v_1668 = vout_canPeek_1669 & 1'h1;
  pebbles_core
    pebbles_core_1669
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1666),
       .in0_consume_en(vin0_consume_en_1669),
       .out_canPeek(vout_canPeek_1669),
       .out_peek(vout_peek_1669));
  assign v_1670 = mux_1670(v_1671);
  assign v_1671 = ~v_1668;
  assign v_1672 = v_1673 | v_1678;
  assign v_1673 = mux_1673(v_1674);
  assign v_1674 = v_1675 & 1'h1;
  assign v_1675 = v_1676 & vout_canPeek_1677;
  assign v_1676 = ~vout_canPeek_1669;
  pebbles_core
    pebbles_core_1677
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1672),
       .in0_consume_en(vin0_consume_en_1677),
       .out_canPeek(vout_canPeek_1677),
       .out_peek(vout_peek_1677));
  assign v_1678 = mux_1678(v_1679);
  assign v_1679 = ~v_1674;
  assign v_1680 = v_1681 | v_1684;
  assign v_1681 = mux_1681(v_1682);
  assign v_1682 = vout_canPeek_1683 & 1'h1;
  pebbles_core
    pebbles_core_1683
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1680),
       .in0_consume_en(vin0_consume_en_1683),
       .out_canPeek(vout_canPeek_1683),
       .out_peek(vout_peek_1683));
  assign v_1684 = mux_1684(v_1685);
  assign v_1685 = ~v_1682;
  assign v_1686 = v_1687 | v_1692;
  assign v_1687 = mux_1687(v_1688);
  assign v_1688 = v_1689 & 1'h1;
  assign v_1689 = v_1690 & vout_canPeek_1691;
  assign v_1690 = ~vout_canPeek_1683;
  pebbles_core
    pebbles_core_1691
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1686),
       .in0_consume_en(vin0_consume_en_1691),
       .out_canPeek(vout_canPeek_1691),
       .out_peek(vout_peek_1691));
  assign v_1692 = mux_1692(v_1693);
  assign v_1693 = ~v_1688;
  assign v_1694 = v_1695 | v_1698;
  assign v_1695 = mux_1695(v_1696);
  assign v_1696 = vout_canPeek_1697 & 1'h1;
  pebbles_core
    pebbles_core_1697
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1694),
       .in0_consume_en(vin0_consume_en_1697),
       .out_canPeek(vout_canPeek_1697),
       .out_peek(vout_peek_1697));
  assign v_1698 = mux_1698(v_1699);
  assign v_1699 = ~v_1696;
  assign v_1700 = v_1701 | v_1706;
  assign v_1701 = mux_1701(v_1702);
  assign v_1702 = v_1703 & 1'h1;
  assign v_1703 = v_1704 & vout_canPeek_1705;
  assign v_1704 = ~vout_canPeek_1697;
  pebbles_core
    pebbles_core_1705
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1700),
       .in0_consume_en(vin0_consume_en_1705),
       .out_canPeek(vout_canPeek_1705),
       .out_peek(vout_peek_1705));
  assign v_1706 = mux_1706(v_1707);
  assign v_1707 = ~v_1702;
  assign v_1708 = v_1709 | v_1712;
  assign v_1709 = mux_1709(v_1710);
  assign v_1710 = vout_canPeek_1711 & 1'h1;
  pebbles_core
    pebbles_core_1711
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1708),
       .in0_consume_en(vin0_consume_en_1711),
       .out_canPeek(vout_canPeek_1711),
       .out_peek(vout_peek_1711));
  assign v_1712 = mux_1712(v_1713);
  assign v_1713 = ~v_1710;
  assign v_1714 = v_1715 | v_1720;
  assign v_1715 = mux_1715(v_1716);
  assign v_1716 = v_1717 & 1'h1;
  assign v_1717 = v_1718 & vout_canPeek_1719;
  assign v_1718 = ~vout_canPeek_1711;
  pebbles_core
    pebbles_core_1719
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1714),
       .in0_consume_en(vin0_consume_en_1719),
       .out_canPeek(vout_canPeek_1719),
       .out_peek(vout_peek_1719));
  assign v_1720 = mux_1720(v_1721);
  assign v_1721 = ~v_1716;
  assign v_1722 = v_1723 | v_1726;
  assign v_1723 = mux_1723(v_1724);
  assign v_1724 = vout_canPeek_1725 & 1'h1;
  pebbles_core
    pebbles_core_1725
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1722),
       .in0_consume_en(vin0_consume_en_1725),
       .out_canPeek(vout_canPeek_1725),
       .out_peek(vout_peek_1725));
  assign v_1726 = mux_1726(v_1727);
  assign v_1727 = ~v_1724;
  assign v_1728 = v_1729 | v_1734;
  assign v_1729 = mux_1729(v_1730);
  assign v_1730 = v_1731 & 1'h1;
  assign v_1731 = v_1732 & vout_canPeek_1733;
  assign v_1732 = ~vout_canPeek_1725;
  pebbles_core
    pebbles_core_1733
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1728),
       .in0_consume_en(vin0_consume_en_1733),
       .out_canPeek(vout_canPeek_1733),
       .out_peek(vout_peek_1733));
  assign v_1734 = mux_1734(v_1735);
  assign v_1735 = ~v_1730;
  assign v_1736 = v_1737 | v_1740;
  assign v_1737 = mux_1737(v_1738);
  assign v_1738 = vout_canPeek_1739 & 1'h1;
  pebbles_core
    pebbles_core_1739
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1736),
       .in0_consume_en(vin0_consume_en_1739),
       .out_canPeek(vout_canPeek_1739),
       .out_peek(vout_peek_1739));
  assign v_1740 = mux_1740(v_1741);
  assign v_1741 = ~v_1738;
  assign v_1742 = v_1743 | v_1748;
  assign v_1743 = mux_1743(v_1744);
  assign v_1744 = v_1745 & 1'h1;
  assign v_1745 = v_1746 & vout_canPeek_1747;
  assign v_1746 = ~vout_canPeek_1739;
  pebbles_core
    pebbles_core_1747
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1742),
       .in0_consume_en(vin0_consume_en_1747),
       .out_canPeek(vout_canPeek_1747),
       .out_peek(vout_peek_1747));
  assign v_1748 = mux_1748(v_1749);
  assign v_1749 = ~v_1744;
  assign v_1750 = v_1751 | v_1754;
  assign v_1751 = mux_1751(v_1752);
  assign v_1752 = vout_canPeek_1753 & 1'h1;
  pebbles_core
    pebbles_core_1753
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1750),
       .in0_consume_en(vin0_consume_en_1753),
       .out_canPeek(vout_canPeek_1753),
       .out_peek(vout_peek_1753));
  assign v_1754 = mux_1754(v_1755);
  assign v_1755 = ~v_1752;
  assign v_1756 = v_1757 | v_1762;
  assign v_1757 = mux_1757(v_1758);
  assign v_1758 = v_1759 & 1'h1;
  assign v_1759 = v_1760 & vout_canPeek_1761;
  assign v_1760 = ~vout_canPeek_1753;
  pebbles_core
    pebbles_core_1761
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1756),
       .in0_consume_en(vin0_consume_en_1761),
       .out_canPeek(vout_canPeek_1761),
       .out_peek(vout_peek_1761));
  assign v_1762 = mux_1762(v_1763);
  assign v_1763 = ~v_1758;
  assign v_1764 = v_1765 | v_1768;
  assign v_1765 = mux_1765(v_1766);
  assign v_1766 = vout_canPeek_1767 & 1'h1;
  pebbles_core
    pebbles_core_1767
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1764),
       .in0_consume_en(vin0_consume_en_1767),
       .out_canPeek(vout_canPeek_1767),
       .out_peek(vout_peek_1767));
  assign v_1768 = mux_1768(v_1769);
  assign v_1769 = ~v_1766;
  assign v_1770 = v_1771 | v_1776;
  assign v_1771 = mux_1771(v_1772);
  assign v_1772 = v_1773 & 1'h1;
  assign v_1773 = v_1774 & vout_canPeek_1775;
  assign v_1774 = ~vout_canPeek_1767;
  pebbles_core
    pebbles_core_1775
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1770),
       .in0_consume_en(vin0_consume_en_1775),
       .out_canPeek(vout_canPeek_1775),
       .out_peek(vout_peek_1775));
  assign v_1776 = mux_1776(v_1777);
  assign v_1777 = ~v_1772;
  assign v_1778 = v_1779 | v_1782;
  assign v_1779 = mux_1779(v_1780);
  assign v_1780 = vout_canPeek_1781 & 1'h1;
  pebbles_core
    pebbles_core_1781
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1778),
       .in0_consume_en(vin0_consume_en_1781),
       .out_canPeek(vout_canPeek_1781),
       .out_peek(vout_peek_1781));
  assign v_1782 = mux_1782(v_1783);
  assign v_1783 = ~v_1780;
  assign v_1784 = v_1785 | v_1790;
  assign v_1785 = mux_1785(v_1786);
  assign v_1786 = v_1787 & 1'h1;
  assign v_1787 = v_1788 & vout_canPeek_1789;
  assign v_1788 = ~vout_canPeek_1781;
  pebbles_core
    pebbles_core_1789
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1784),
       .in0_consume_en(vin0_consume_en_1789),
       .out_canPeek(vout_canPeek_1789),
       .out_peek(vout_peek_1789));
  assign v_1790 = mux_1790(v_1791);
  assign v_1791 = ~v_1786;
  assign v_1792 = v_1793 | v_1796;
  assign v_1793 = mux_1793(v_1794);
  assign v_1794 = vout_canPeek_1795 & 1'h1;
  pebbles_core
    pebbles_core_1795
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1792),
       .in0_consume_en(vin0_consume_en_1795),
       .out_canPeek(vout_canPeek_1795),
       .out_peek(vout_peek_1795));
  assign v_1796 = mux_1796(v_1797);
  assign v_1797 = ~v_1794;
  assign v_1798 = v_1799 | v_1804;
  assign v_1799 = mux_1799(v_1800);
  assign v_1800 = v_1801 & 1'h1;
  assign v_1801 = v_1802 & vout_canPeek_1803;
  assign v_1802 = ~vout_canPeek_1795;
  pebbles_core
    pebbles_core_1803
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1798),
       .in0_consume_en(vin0_consume_en_1803),
       .out_canPeek(vout_canPeek_1803),
       .out_peek(vout_peek_1803));
  assign v_1804 = mux_1804(v_1805);
  assign v_1805 = ~v_1800;
  assign v_1806 = v_1807 | v_1810;
  assign v_1807 = mux_1807(v_1808);
  assign v_1808 = vout_canPeek_1809 & 1'h1;
  pebbles_core
    pebbles_core_1809
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1806),
       .in0_consume_en(vin0_consume_en_1809),
       .out_canPeek(vout_canPeek_1809),
       .out_peek(vout_peek_1809));
  assign v_1810 = mux_1810(v_1811);
  assign v_1811 = ~v_1808;
  assign v_1812 = v_1813 | v_1818;
  assign v_1813 = mux_1813(v_1814);
  assign v_1814 = v_1815 & 1'h1;
  assign v_1815 = v_1816 & vout_canPeek_1817;
  assign v_1816 = ~vout_canPeek_1809;
  pebbles_core
    pebbles_core_1817
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1812),
       .in0_consume_en(vin0_consume_en_1817),
       .out_canPeek(vout_canPeek_1817),
       .out_peek(vout_peek_1817));
  assign v_1818 = mux_1818(v_1819);
  assign v_1819 = ~v_1814;
  assign v_1820 = v_1821 | v_1824;
  assign v_1821 = mux_1821(v_1822);
  assign v_1822 = vout_canPeek_1823 & 1'h1;
  pebbles_core
    pebbles_core_1823
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1820),
       .in0_consume_en(vin0_consume_en_1823),
       .out_canPeek(vout_canPeek_1823),
       .out_peek(vout_peek_1823));
  assign v_1824 = mux_1824(v_1825);
  assign v_1825 = ~v_1822;
  assign v_1826 = v_1827 | v_1832;
  assign v_1827 = mux_1827(v_1828);
  assign v_1828 = v_1829 & 1'h1;
  assign v_1829 = v_1830 & vout_canPeek_1831;
  assign v_1830 = ~vout_canPeek_1823;
  pebbles_core
    pebbles_core_1831
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1826),
       .in0_consume_en(vin0_consume_en_1831),
       .out_canPeek(vout_canPeek_1831),
       .out_peek(vout_peek_1831));
  assign v_1832 = mux_1832(v_1833);
  assign v_1833 = ~v_1828;
  assign v_1834 = v_1835 | v_1838;
  assign v_1835 = mux_1835(v_1836);
  assign v_1836 = vout_canPeek_1837 & 1'h1;
  pebbles_core
    pebbles_core_1837
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1834),
       .in0_consume_en(vin0_consume_en_1837),
       .out_canPeek(vout_canPeek_1837),
       .out_peek(vout_peek_1837));
  assign v_1838 = mux_1838(v_1839);
  assign v_1839 = ~v_1836;
  assign v_1840 = v_1841 | v_1846;
  assign v_1841 = mux_1841(v_1842);
  assign v_1842 = v_1843 & 1'h1;
  assign v_1843 = v_1844 & vout_canPeek_1845;
  assign v_1844 = ~vout_canPeek_1837;
  pebbles_core
    pebbles_core_1845
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1840),
       .in0_consume_en(vin0_consume_en_1845),
       .out_canPeek(vout_canPeek_1845),
       .out_peek(vout_peek_1845));
  assign v_1846 = mux_1846(v_1847);
  assign v_1847 = ~v_1842;
  assign v_1848 = v_1849 | v_1852;
  assign v_1849 = mux_1849(v_1850);
  assign v_1850 = vout_canPeek_1851 & 1'h1;
  pebbles_core
    pebbles_core_1851
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1848),
       .in0_consume_en(vin0_consume_en_1851),
       .out_canPeek(vout_canPeek_1851),
       .out_peek(vout_peek_1851));
  assign v_1852 = mux_1852(v_1853);
  assign v_1853 = ~v_1850;
  assign v_1854 = v_1855 | v_1860;
  assign v_1855 = mux_1855(v_1856);
  assign v_1856 = v_1857 & 1'h1;
  assign v_1857 = v_1858 & vout_canPeek_1859;
  assign v_1858 = ~vout_canPeek_1851;
  pebbles_core
    pebbles_core_1859
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1854),
       .in0_consume_en(vin0_consume_en_1859),
       .out_canPeek(vout_canPeek_1859),
       .out_peek(vout_peek_1859));
  assign v_1860 = mux_1860(v_1861);
  assign v_1861 = ~v_1856;
  assign v_1862 = v_1863 | v_1866;
  assign v_1863 = mux_1863(v_1864);
  assign v_1864 = vout_canPeek_1865 & 1'h1;
  pebbles_core
    pebbles_core_1865
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1862),
       .in0_consume_en(vin0_consume_en_1865),
       .out_canPeek(vout_canPeek_1865),
       .out_peek(vout_peek_1865));
  assign v_1866 = mux_1866(v_1867);
  assign v_1867 = ~v_1864;
  assign v_1868 = v_1869 | v_1874;
  assign v_1869 = mux_1869(v_1870);
  assign v_1870 = v_1871 & 1'h1;
  assign v_1871 = v_1872 & vout_canPeek_1873;
  assign v_1872 = ~vout_canPeek_1865;
  pebbles_core
    pebbles_core_1873
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1868),
       .in0_consume_en(vin0_consume_en_1873),
       .out_canPeek(vout_canPeek_1873),
       .out_peek(vout_peek_1873));
  assign v_1874 = mux_1874(v_1875);
  assign v_1875 = ~v_1870;
  assign v_1876 = v_1877 | v_1880;
  assign v_1877 = mux_1877(v_1878);
  assign v_1878 = vout_canPeek_1879 & 1'h1;
  pebbles_core
    pebbles_core_1879
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1876),
       .in0_consume_en(vin0_consume_en_1879),
       .out_canPeek(vout_canPeek_1879),
       .out_peek(vout_peek_1879));
  assign v_1880 = mux_1880(v_1881);
  assign v_1881 = ~v_1878;
  assign v_1882 = v_1883 | v_1888;
  assign v_1883 = mux_1883(v_1884);
  assign v_1884 = v_1885 & 1'h1;
  assign v_1885 = v_1886 & vout_canPeek_1887;
  assign v_1886 = ~vout_canPeek_1879;
  pebbles_core
    pebbles_core_1887
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1882),
       .in0_consume_en(vin0_consume_en_1887),
       .out_canPeek(vout_canPeek_1887),
       .out_peek(vout_peek_1887));
  assign v_1888 = mux_1888(v_1889);
  assign v_1889 = ~v_1884;
  assign v_1890 = v_1891 | v_1894;
  assign v_1891 = mux_1891(v_1892);
  assign v_1892 = vout_canPeek_1893 & 1'h1;
  pebbles_core
    pebbles_core_1893
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1890),
       .in0_consume_en(vin0_consume_en_1893),
       .out_canPeek(vout_canPeek_1893),
       .out_peek(vout_peek_1893));
  assign v_1894 = mux_1894(v_1895);
  assign v_1895 = ~v_1892;
  assign v_1896 = v_1897 | v_1902;
  assign v_1897 = mux_1897(v_1898);
  assign v_1898 = v_1899 & 1'h1;
  assign v_1899 = v_1900 & vout_canPeek_1901;
  assign v_1900 = ~vout_canPeek_1893;
  pebbles_core
    pebbles_core_1901
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1896),
       .in0_consume_en(vin0_consume_en_1901),
       .out_canPeek(vout_canPeek_1901),
       .out_peek(vout_peek_1901));
  assign v_1902 = mux_1902(v_1903);
  assign v_1903 = ~v_1898;
  assign v_1904 = v_1905 | v_1908;
  assign v_1905 = mux_1905(v_1906);
  assign v_1906 = vout_canPeek_1907 & 1'h1;
  pebbles_core
    pebbles_core_1907
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1904),
       .in0_consume_en(vin0_consume_en_1907),
       .out_canPeek(vout_canPeek_1907),
       .out_peek(vout_peek_1907));
  assign v_1908 = mux_1908(v_1909);
  assign v_1909 = ~v_1906;
  assign v_1910 = v_1911 | v_1916;
  assign v_1911 = mux_1911(v_1912);
  assign v_1912 = v_1913 & 1'h1;
  assign v_1913 = v_1914 & vout_canPeek_1915;
  assign v_1914 = ~vout_canPeek_1907;
  pebbles_core
    pebbles_core_1915
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1910),
       .in0_consume_en(vin0_consume_en_1915),
       .out_canPeek(vout_canPeek_1915),
       .out_peek(vout_peek_1915));
  assign v_1916 = mux_1916(v_1917);
  assign v_1917 = ~v_1912;
  assign v_1918 = v_1919 | v_1922;
  assign v_1919 = mux_1919(v_1920);
  assign v_1920 = vout_canPeek_1921 & 1'h1;
  pebbles_core
    pebbles_core_1921
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1918),
       .in0_consume_en(vin0_consume_en_1921),
       .out_canPeek(vout_canPeek_1921),
       .out_peek(vout_peek_1921));
  assign v_1922 = mux_1922(v_1923);
  assign v_1923 = ~v_1920;
  assign v_1924 = v_1925 | v_1930;
  assign v_1925 = mux_1925(v_1926);
  assign v_1926 = v_1927 & 1'h1;
  assign v_1927 = v_1928 & vout_canPeek_1929;
  assign v_1928 = ~vout_canPeek_1921;
  pebbles_core
    pebbles_core_1929
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1924),
       .in0_consume_en(vin0_consume_en_1929),
       .out_canPeek(vout_canPeek_1929),
       .out_peek(vout_peek_1929));
  assign v_1930 = mux_1930(v_1931);
  assign v_1931 = ~v_1926;
  assign v_1932 = v_1933 | v_1936;
  assign v_1933 = mux_1933(v_1934);
  assign v_1934 = vout_canPeek_1935 & 1'h1;
  pebbles_core
    pebbles_core_1935
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1932),
       .in0_consume_en(vin0_consume_en_1935),
       .out_canPeek(vout_canPeek_1935),
       .out_peek(vout_peek_1935));
  assign v_1936 = mux_1936(v_1937);
  assign v_1937 = ~v_1934;
  assign v_1938 = v_1939 | v_1944;
  assign v_1939 = mux_1939(v_1940);
  assign v_1940 = v_1941 & 1'h1;
  assign v_1941 = v_1942 & vout_canPeek_1943;
  assign v_1942 = ~vout_canPeek_1935;
  pebbles_core
    pebbles_core_1943
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1938),
       .in0_consume_en(vin0_consume_en_1943),
       .out_canPeek(vout_canPeek_1943),
       .out_peek(vout_peek_1943));
  assign v_1944 = mux_1944(v_1945);
  assign v_1945 = ~v_1940;
  assign v_1946 = v_1947 | v_1950;
  assign v_1947 = mux_1947(v_1948);
  assign v_1948 = vout_canPeek_1949 & 1'h1;
  pebbles_core
    pebbles_core_1949
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1946),
       .in0_consume_en(vin0_consume_en_1949),
       .out_canPeek(vout_canPeek_1949),
       .out_peek(vout_peek_1949));
  assign v_1950 = mux_1950(v_1951);
  assign v_1951 = ~v_1948;
  assign v_1952 = v_1953 | v_1958;
  assign v_1953 = mux_1953(v_1954);
  assign v_1954 = v_1955 & 1'h1;
  assign v_1955 = v_1956 & vout_canPeek_1957;
  assign v_1956 = ~vout_canPeek_1949;
  pebbles_core
    pebbles_core_1957
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1952),
       .in0_consume_en(vin0_consume_en_1957),
       .out_canPeek(vout_canPeek_1957),
       .out_peek(vout_peek_1957));
  assign v_1958 = mux_1958(v_1959);
  assign v_1959 = ~v_1954;
  assign v_1960 = v_1961 | v_1964;
  assign v_1961 = mux_1961(v_1962);
  assign v_1962 = vout_canPeek_1963 & 1'h1;
  pebbles_core
    pebbles_core_1963
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1960),
       .in0_consume_en(vin0_consume_en_1963),
       .out_canPeek(vout_canPeek_1963),
       .out_peek(vout_peek_1963));
  assign v_1964 = mux_1964(v_1965);
  assign v_1965 = ~v_1962;
  assign v_1966 = v_1967 | v_1972;
  assign v_1967 = mux_1967(v_1968);
  assign v_1968 = v_1969 & 1'h1;
  assign v_1969 = v_1970 & vout_canPeek_1971;
  assign v_1970 = ~vout_canPeek_1963;
  pebbles_core
    pebbles_core_1971
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1966),
       .in0_consume_en(vin0_consume_en_1971),
       .out_canPeek(vout_canPeek_1971),
       .out_peek(vout_peek_1971));
  assign v_1972 = mux_1972(v_1973);
  assign v_1973 = ~v_1968;
  assign v_1974 = v_1975 | v_1978;
  assign v_1975 = mux_1975(v_1976);
  assign v_1976 = vout_canPeek_1977 & 1'h1;
  pebbles_core
    pebbles_core_1977
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1974),
       .in0_consume_en(vin0_consume_en_1977),
       .out_canPeek(vout_canPeek_1977),
       .out_peek(vout_peek_1977));
  assign v_1978 = mux_1978(v_1979);
  assign v_1979 = ~v_1976;
  assign v_1980 = v_1981 | v_1986;
  assign v_1981 = mux_1981(v_1982);
  assign v_1982 = v_1983 & 1'h1;
  assign v_1983 = v_1984 & vout_canPeek_1985;
  assign v_1984 = ~vout_canPeek_1977;
  pebbles_core
    pebbles_core_1985
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1980),
       .in0_consume_en(vin0_consume_en_1985),
       .out_canPeek(vout_canPeek_1985),
       .out_peek(vout_peek_1985));
  assign v_1986 = mux_1986(v_1987);
  assign v_1987 = ~v_1982;
  assign v_1988 = v_1989 | v_1992;
  assign v_1989 = mux_1989(v_1990);
  assign v_1990 = vout_canPeek_1991 & 1'h1;
  pebbles_core
    pebbles_core_1991
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1988),
       .in0_consume_en(vin0_consume_en_1991),
       .out_canPeek(vout_canPeek_1991),
       .out_peek(vout_peek_1991));
  assign v_1992 = mux_1992(v_1993);
  assign v_1993 = ~v_1990;
  assign v_1994 = v_1995 | v_2000;
  assign v_1995 = mux_1995(v_1996);
  assign v_1996 = v_1997 & 1'h1;
  assign v_1997 = v_1998 & vout_canPeek_1999;
  assign v_1998 = ~vout_canPeek_1991;
  pebbles_core
    pebbles_core_1999
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_1994),
       .in0_consume_en(vin0_consume_en_1999),
       .out_canPeek(vout_canPeek_1999),
       .out_peek(vout_peek_1999));
  assign v_2000 = mux_2000(v_2001);
  assign v_2001 = ~v_1996;
  assign v_2002 = v_2003 | v_2006;
  assign v_2003 = mux_2003(v_2004);
  assign v_2004 = vout_canPeek_2005 & 1'h1;
  pebbles_core
    pebbles_core_2005
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2002),
       .in0_consume_en(vin0_consume_en_2005),
       .out_canPeek(vout_canPeek_2005),
       .out_peek(vout_peek_2005));
  assign v_2006 = mux_2006(v_2007);
  assign v_2007 = ~v_2004;
  assign v_2008 = v_2009 | v_2014;
  assign v_2009 = mux_2009(v_2010);
  assign v_2010 = v_2011 & 1'h1;
  assign v_2011 = v_2012 & vout_canPeek_2013;
  assign v_2012 = ~vout_canPeek_2005;
  pebbles_core
    pebbles_core_2013
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2008),
       .in0_consume_en(vin0_consume_en_2013),
       .out_canPeek(vout_canPeek_2013),
       .out_peek(vout_peek_2013));
  assign v_2014 = mux_2014(v_2015);
  assign v_2015 = ~v_2010;
  assign v_2016 = v_2017 | v_2020;
  assign v_2017 = mux_2017(v_2018);
  assign v_2018 = vout_canPeek_2019 & 1'h1;
  pebbles_core
    pebbles_core_2019
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2016),
       .in0_consume_en(vin0_consume_en_2019),
       .out_canPeek(vout_canPeek_2019),
       .out_peek(vout_peek_2019));
  assign v_2020 = mux_2020(v_2021);
  assign v_2021 = ~v_2018;
  assign v_2022 = v_2023 | v_2028;
  assign v_2023 = mux_2023(v_2024);
  assign v_2024 = v_2025 & 1'h1;
  assign v_2025 = v_2026 & vout_canPeek_2027;
  assign v_2026 = ~vout_canPeek_2019;
  pebbles_core
    pebbles_core_2027
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2022),
       .in0_consume_en(vin0_consume_en_2027),
       .out_canPeek(vout_canPeek_2027),
       .out_peek(vout_peek_2027));
  assign v_2028 = mux_2028(v_2029);
  assign v_2029 = ~v_2024;
  assign v_2030 = v_2031 | v_2034;
  assign v_2031 = mux_2031(v_2032);
  assign v_2032 = vout_canPeek_2033 & 1'h1;
  pebbles_core
    pebbles_core_2033
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2030),
       .in0_consume_en(vin0_consume_en_2033),
       .out_canPeek(vout_canPeek_2033),
       .out_peek(vout_peek_2033));
  assign v_2034 = mux_2034(v_2035);
  assign v_2035 = ~v_2032;
  assign v_2036 = v_2037 | v_2042;
  assign v_2037 = mux_2037(v_2038);
  assign v_2038 = v_2039 & 1'h1;
  assign v_2039 = v_2040 & vout_canPeek_2041;
  assign v_2040 = ~vout_canPeek_2033;
  pebbles_core
    pebbles_core_2041
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2036),
       .in0_consume_en(vin0_consume_en_2041),
       .out_canPeek(vout_canPeek_2041),
       .out_peek(vout_peek_2041));
  assign v_2042 = mux_2042(v_2043);
  assign v_2043 = ~v_2038;
  assign v_2044 = v_2045 | v_2048;
  assign v_2045 = mux_2045(v_2046);
  assign v_2046 = vout_canPeek_2047 & 1'h1;
  pebbles_core
    pebbles_core_2047
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2044),
       .in0_consume_en(vin0_consume_en_2047),
       .out_canPeek(vout_canPeek_2047),
       .out_peek(vout_peek_2047));
  assign v_2048 = mux_2048(v_2049);
  assign v_2049 = ~v_2046;
  assign v_2050 = v_2051 | v_2056;
  assign v_2051 = mux_2051(v_2052);
  assign v_2052 = v_2053 & 1'h1;
  assign v_2053 = v_2054 & vout_canPeek_2055;
  assign v_2054 = ~vout_canPeek_2047;
  pebbles_core
    pebbles_core_2055
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2050),
       .in0_consume_en(vin0_consume_en_2055),
       .out_canPeek(vout_canPeek_2055),
       .out_peek(vout_peek_2055));
  assign v_2056 = mux_2056(v_2057);
  assign v_2057 = ~v_2052;
  assign v_2058 = v_2059 | v_2062;
  assign v_2059 = mux_2059(v_2060);
  assign v_2060 = vout_canPeek_2061 & 1'h1;
  pebbles_core
    pebbles_core_2061
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2058),
       .in0_consume_en(vin0_consume_en_2061),
       .out_canPeek(vout_canPeek_2061),
       .out_peek(vout_peek_2061));
  assign v_2062 = mux_2062(v_2063);
  assign v_2063 = ~v_2060;
  assign v_2064 = v_2065 | v_2070;
  assign v_2065 = mux_2065(v_2066);
  assign v_2066 = v_2067 & 1'h1;
  assign v_2067 = v_2068 & vout_canPeek_2069;
  assign v_2068 = ~vout_canPeek_2061;
  pebbles_core
    pebbles_core_2069
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2064),
       .in0_consume_en(vin0_consume_en_2069),
       .out_canPeek(vout_canPeek_2069),
       .out_peek(vout_peek_2069));
  assign v_2070 = mux_2070(v_2071);
  assign v_2071 = ~v_2066;
  assign v_2072 = v_2073 | v_2076;
  assign v_2073 = mux_2073(v_2074);
  assign v_2074 = vout_canPeek_2075 & 1'h1;
  pebbles_core
    pebbles_core_2075
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2072),
       .in0_consume_en(vin0_consume_en_2075),
       .out_canPeek(vout_canPeek_2075),
       .out_peek(vout_peek_2075));
  assign v_2076 = mux_2076(v_2077);
  assign v_2077 = ~v_2074;
  assign v_2078 = v_2079 | v_2084;
  assign v_2079 = mux_2079(v_2080);
  assign v_2080 = v_2081 & 1'h1;
  assign v_2081 = v_2082 & vout_canPeek_2083;
  assign v_2082 = ~vout_canPeek_2075;
  pebbles_core
    pebbles_core_2083
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2078),
       .in0_consume_en(vin0_consume_en_2083),
       .out_canPeek(vout_canPeek_2083),
       .out_peek(vout_peek_2083));
  assign v_2084 = mux_2084(v_2085);
  assign v_2085 = ~v_2080;
  assign v_2086 = v_2087 | v_2090;
  assign v_2087 = mux_2087(v_2088);
  assign v_2088 = vout_canPeek_2089 & 1'h1;
  pebbles_core
    pebbles_core_2089
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2086),
       .in0_consume_en(vin0_consume_en_2089),
       .out_canPeek(vout_canPeek_2089),
       .out_peek(vout_peek_2089));
  assign v_2090 = mux_2090(v_2091);
  assign v_2091 = ~v_2088;
  assign v_2092 = v_2093 | v_2098;
  assign v_2093 = mux_2093(v_2094);
  assign v_2094 = v_2095 & 1'h1;
  assign v_2095 = v_2096 & vout_canPeek_2097;
  assign v_2096 = ~vout_canPeek_2089;
  pebbles_core
    pebbles_core_2097
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2092),
       .in0_consume_en(vin0_consume_en_2097),
       .out_canPeek(vout_canPeek_2097),
       .out_peek(vout_peek_2097));
  assign v_2098 = mux_2098(v_2099);
  assign v_2099 = ~v_2094;
  assign v_2100 = v_2101 | v_2104;
  assign v_2101 = mux_2101(v_2102);
  assign v_2102 = vout_canPeek_2103 & 1'h1;
  pebbles_core
    pebbles_core_2103
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2100),
       .in0_consume_en(vin0_consume_en_2103),
       .out_canPeek(vout_canPeek_2103),
       .out_peek(vout_peek_2103));
  assign v_2104 = mux_2104(v_2105);
  assign v_2105 = ~v_2102;
  assign v_2106 = v_2107 | v_2112;
  assign v_2107 = mux_2107(v_2108);
  assign v_2108 = v_2109 & 1'h1;
  assign v_2109 = v_2110 & vout_canPeek_2111;
  assign v_2110 = ~vout_canPeek_2103;
  pebbles_core
    pebbles_core_2111
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2106),
       .in0_consume_en(vin0_consume_en_2111),
       .out_canPeek(vout_canPeek_2111),
       .out_peek(vout_peek_2111));
  assign v_2112 = mux_2112(v_2113);
  assign v_2113 = ~v_2108;
  assign v_2114 = v_2115 | v_2118;
  assign v_2115 = mux_2115(v_2116);
  assign v_2116 = vout_canPeek_2117 & 1'h1;
  pebbles_core
    pebbles_core_2117
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2114),
       .in0_consume_en(vin0_consume_en_2117),
       .out_canPeek(vout_canPeek_2117),
       .out_peek(vout_peek_2117));
  assign v_2118 = mux_2118(v_2119);
  assign v_2119 = ~v_2116;
  assign v_2120 = v_2121 | v_2126;
  assign v_2121 = mux_2121(v_2122);
  assign v_2122 = v_2123 & 1'h1;
  assign v_2123 = v_2124 & vout_canPeek_2125;
  assign v_2124 = ~vout_canPeek_2117;
  pebbles_core
    pebbles_core_2125
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2120),
       .in0_consume_en(vin0_consume_en_2125),
       .out_canPeek(vout_canPeek_2125),
       .out_peek(vout_peek_2125));
  assign v_2126 = mux_2126(v_2127);
  assign v_2127 = ~v_2122;
  assign v_2128 = v_2129 | v_2132;
  assign v_2129 = mux_2129(v_2130);
  assign v_2130 = vout_canPeek_2131 & 1'h1;
  pebbles_core
    pebbles_core_2131
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2128),
       .in0_consume_en(vin0_consume_en_2131),
       .out_canPeek(vout_canPeek_2131),
       .out_peek(vout_peek_2131));
  assign v_2132 = mux_2132(v_2133);
  assign v_2133 = ~v_2130;
  assign v_2134 = v_2135 | v_2140;
  assign v_2135 = mux_2135(v_2136);
  assign v_2136 = v_2137 & 1'h1;
  assign v_2137 = v_2138 & vout_canPeek_2139;
  assign v_2138 = ~vout_canPeek_2131;
  pebbles_core
    pebbles_core_2139
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2134),
       .in0_consume_en(vin0_consume_en_2139),
       .out_canPeek(vout_canPeek_2139),
       .out_peek(vout_peek_2139));
  assign v_2140 = mux_2140(v_2141);
  assign v_2141 = ~v_2136;
  assign v_2142 = v_2143 | v_2146;
  assign v_2143 = mux_2143(v_2144);
  assign v_2144 = vout_canPeek_2145 & 1'h1;
  pebbles_core
    pebbles_core_2145
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2142),
       .in0_consume_en(vin0_consume_en_2145),
       .out_canPeek(vout_canPeek_2145),
       .out_peek(vout_peek_2145));
  assign v_2146 = mux_2146(v_2147);
  assign v_2147 = ~v_2144;
  assign v_2148 = v_2149 | v_2154;
  assign v_2149 = mux_2149(v_2150);
  assign v_2150 = v_2151 & 1'h1;
  assign v_2151 = v_2152 & vout_canPeek_2153;
  assign v_2152 = ~vout_canPeek_2145;
  pebbles_core
    pebbles_core_2153
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2148),
       .in0_consume_en(vin0_consume_en_2153),
       .out_canPeek(vout_canPeek_2153),
       .out_peek(vout_peek_2153));
  assign v_2154 = mux_2154(v_2155);
  assign v_2155 = ~v_2150;
  assign v_2156 = v_2157 | v_2160;
  assign v_2157 = mux_2157(v_2158);
  assign v_2158 = vout_canPeek_2159 & 1'h1;
  pebbles_core
    pebbles_core_2159
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2156),
       .in0_consume_en(vin0_consume_en_2159),
       .out_canPeek(vout_canPeek_2159),
       .out_peek(vout_peek_2159));
  assign v_2160 = mux_2160(v_2161);
  assign v_2161 = ~v_2158;
  assign v_2162 = v_2163 | v_2168;
  assign v_2163 = mux_2163(v_2164);
  assign v_2164 = v_2165 & 1'h1;
  assign v_2165 = v_2166 & vout_canPeek_2167;
  assign v_2166 = ~vout_canPeek_2159;
  pebbles_core
    pebbles_core_2167
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2162),
       .in0_consume_en(vin0_consume_en_2167),
       .out_canPeek(vout_canPeek_2167),
       .out_peek(vout_peek_2167));
  assign v_2168 = mux_2168(v_2169);
  assign v_2169 = ~v_2164;
  assign v_2170 = v_2171 | v_2174;
  assign v_2171 = mux_2171(v_2172);
  assign v_2172 = vout_canPeek_2173 & 1'h1;
  pebbles_core
    pebbles_core_2173
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2170),
       .in0_consume_en(vin0_consume_en_2173),
       .out_canPeek(vout_canPeek_2173),
       .out_peek(vout_peek_2173));
  assign v_2174 = mux_2174(v_2175);
  assign v_2175 = ~v_2172;
  assign v_2176 = v_2177 | v_2182;
  assign v_2177 = mux_2177(v_2178);
  assign v_2178 = v_2179 & 1'h1;
  assign v_2179 = v_2180 & vout_canPeek_2181;
  assign v_2180 = ~vout_canPeek_2173;
  pebbles_core
    pebbles_core_2181
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2176),
       .in0_consume_en(vin0_consume_en_2181),
       .out_canPeek(vout_canPeek_2181),
       .out_peek(vout_peek_2181));
  assign v_2182 = mux_2182(v_2183);
  assign v_2183 = ~v_2178;
  assign v_2184 = v_2185 | v_2188;
  assign v_2185 = mux_2185(v_2186);
  assign v_2186 = vout_canPeek_2187 & 1'h1;
  pebbles_core
    pebbles_core_2187
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2184),
       .in0_consume_en(vin0_consume_en_2187),
       .out_canPeek(vout_canPeek_2187),
       .out_peek(vout_peek_2187));
  assign v_2188 = mux_2188(v_2189);
  assign v_2189 = ~v_2186;
  assign v_2190 = v_2191 | v_2196;
  assign v_2191 = mux_2191(v_2192);
  assign v_2192 = v_2193 & 1'h1;
  assign v_2193 = v_2194 & vout_canPeek_2195;
  assign v_2194 = ~vout_canPeek_2187;
  pebbles_core
    pebbles_core_2195
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2190),
       .in0_consume_en(vin0_consume_en_2195),
       .out_canPeek(vout_canPeek_2195),
       .out_peek(vout_peek_2195));
  assign v_2196 = mux_2196(v_2197);
  assign v_2197 = ~v_2192;
  assign v_2198 = v_2199 | v_2202;
  assign v_2199 = mux_2199(v_2200);
  assign v_2200 = vout_canPeek_2201 & 1'h1;
  pebbles_core
    pebbles_core_2201
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2198),
       .in0_consume_en(vin0_consume_en_2201),
       .out_canPeek(vout_canPeek_2201),
       .out_peek(vout_peek_2201));
  assign v_2202 = mux_2202(v_2203);
  assign v_2203 = ~v_2200;
  assign v_2204 = v_2205 | v_2210;
  assign v_2205 = mux_2205(v_2206);
  assign v_2206 = v_2207 & 1'h1;
  assign v_2207 = v_2208 & vout_canPeek_2209;
  assign v_2208 = ~vout_canPeek_2201;
  pebbles_core
    pebbles_core_2209
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2204),
       .in0_consume_en(vin0_consume_en_2209),
       .out_canPeek(vout_canPeek_2209),
       .out_peek(vout_peek_2209));
  assign v_2210 = mux_2210(v_2211);
  assign v_2211 = ~v_2206;
  assign v_2212 = v_2213 | v_2216;
  assign v_2213 = mux_2213(v_2214);
  assign v_2214 = vout_canPeek_2215 & 1'h1;
  pebbles_core
    pebbles_core_2215
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2212),
       .in0_consume_en(vin0_consume_en_2215),
       .out_canPeek(vout_canPeek_2215),
       .out_peek(vout_peek_2215));
  assign v_2216 = mux_2216(v_2217);
  assign v_2217 = ~v_2214;
  assign v_2218 = v_2219 | v_2224;
  assign v_2219 = mux_2219(v_2220);
  assign v_2220 = v_2221 & 1'h1;
  assign v_2221 = v_2222 & vout_canPeek_2223;
  assign v_2222 = ~vout_canPeek_2215;
  pebbles_core
    pebbles_core_2223
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2218),
       .in0_consume_en(vin0_consume_en_2223),
       .out_canPeek(vout_canPeek_2223),
       .out_peek(vout_peek_2223));
  assign v_2224 = mux_2224(v_2225);
  assign v_2225 = ~v_2220;
  assign v_2226 = v_2227 | v_2230;
  assign v_2227 = mux_2227(v_2228);
  assign v_2228 = vout_canPeek_2229 & 1'h1;
  pebbles_core
    pebbles_core_2229
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2226),
       .in0_consume_en(vin0_consume_en_2229),
       .out_canPeek(vout_canPeek_2229),
       .out_peek(vout_peek_2229));
  assign v_2230 = mux_2230(v_2231);
  assign v_2231 = ~v_2228;
  assign v_2232 = v_2233 | v_2238;
  assign v_2233 = mux_2233(v_2234);
  assign v_2234 = v_2235 & 1'h1;
  assign v_2235 = v_2236 & vout_canPeek_2237;
  assign v_2236 = ~vout_canPeek_2229;
  pebbles_core
    pebbles_core_2237
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2232),
       .in0_consume_en(vin0_consume_en_2237),
       .out_canPeek(vout_canPeek_2237),
       .out_peek(vout_peek_2237));
  assign v_2238 = mux_2238(v_2239);
  assign v_2239 = ~v_2234;
  assign v_2240 = v_2241 | v_2244;
  assign v_2241 = mux_2241(v_2242);
  assign v_2242 = vout_canPeek_2243 & 1'h1;
  pebbles_core
    pebbles_core_2243
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2240),
       .in0_consume_en(vin0_consume_en_2243),
       .out_canPeek(vout_canPeek_2243),
       .out_peek(vout_peek_2243));
  assign v_2244 = mux_2244(v_2245);
  assign v_2245 = ~v_2242;
  assign v_2246 = v_2247 | v_2252;
  assign v_2247 = mux_2247(v_2248);
  assign v_2248 = v_2249 & 1'h1;
  assign v_2249 = v_2250 & vout_canPeek_2251;
  assign v_2250 = ~vout_canPeek_2243;
  pebbles_core
    pebbles_core_2251
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2246),
       .in0_consume_en(vin0_consume_en_2251),
       .out_canPeek(vout_canPeek_2251),
       .out_peek(vout_peek_2251));
  assign v_2252 = mux_2252(v_2253);
  assign v_2253 = ~v_2248;
  assign v_2254 = v_2255 | v_2258;
  assign v_2255 = mux_2255(v_2256);
  assign v_2256 = vout_canPeek_2257 & 1'h1;
  pebbles_core
    pebbles_core_2257
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2254),
       .in0_consume_en(vin0_consume_en_2257),
       .out_canPeek(vout_canPeek_2257),
       .out_peek(vout_peek_2257));
  assign v_2258 = mux_2258(v_2259);
  assign v_2259 = ~v_2256;
  assign v_2260 = v_2261 | v_2266;
  assign v_2261 = mux_2261(v_2262);
  assign v_2262 = v_2263 & 1'h1;
  assign v_2263 = v_2264 & vout_canPeek_2265;
  assign v_2264 = ~vout_canPeek_2257;
  pebbles_core
    pebbles_core_2265
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2260),
       .in0_consume_en(vin0_consume_en_2265),
       .out_canPeek(vout_canPeek_2265),
       .out_peek(vout_peek_2265));
  assign v_2266 = mux_2266(v_2267);
  assign v_2267 = ~v_2262;
  assign v_2268 = v_2269 | v_2272;
  assign v_2269 = mux_2269(v_2270);
  assign v_2270 = vout_canPeek_2271 & 1'h1;
  pebbles_core
    pebbles_core_2271
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2268),
       .in0_consume_en(vin0_consume_en_2271),
       .out_canPeek(vout_canPeek_2271),
       .out_peek(vout_peek_2271));
  assign v_2272 = mux_2272(v_2273);
  assign v_2273 = ~v_2270;
  assign v_2274 = v_2275 | v_2280;
  assign v_2275 = mux_2275(v_2276);
  assign v_2276 = v_2277 & 1'h1;
  assign v_2277 = v_2278 & vout_canPeek_2279;
  assign v_2278 = ~vout_canPeek_2271;
  pebbles_core
    pebbles_core_2279
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2274),
       .in0_consume_en(vin0_consume_en_2279),
       .out_canPeek(vout_canPeek_2279),
       .out_peek(vout_peek_2279));
  assign v_2280 = mux_2280(v_2281);
  assign v_2281 = ~v_2276;
  assign v_2282 = v_2283 | v_2286;
  assign v_2283 = mux_2283(v_2284);
  assign v_2284 = vout_canPeek_2285 & 1'h1;
  pebbles_core
    pebbles_core_2285
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2282),
       .in0_consume_en(vin0_consume_en_2285),
       .out_canPeek(vout_canPeek_2285),
       .out_peek(vout_peek_2285));
  assign v_2286 = mux_2286(v_2287);
  assign v_2287 = ~v_2284;
  assign v_2288 = v_2289 | v_2294;
  assign v_2289 = mux_2289(v_2290);
  assign v_2290 = v_2291 & 1'h1;
  assign v_2291 = v_2292 & vout_canPeek_2293;
  assign v_2292 = ~vout_canPeek_2285;
  pebbles_core
    pebbles_core_2293
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2288),
       .in0_consume_en(vin0_consume_en_2293),
       .out_canPeek(vout_canPeek_2293),
       .out_peek(vout_peek_2293));
  assign v_2294 = mux_2294(v_2295);
  assign v_2295 = ~v_2290;
  assign v_2296 = v_2297 | v_2300;
  assign v_2297 = mux_2297(v_2298);
  assign v_2298 = vout_canPeek_2299 & 1'h1;
  pebbles_core
    pebbles_core_2299
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2296),
       .in0_consume_en(vin0_consume_en_2299),
       .out_canPeek(vout_canPeek_2299),
       .out_peek(vout_peek_2299));
  assign v_2300 = mux_2300(v_2301);
  assign v_2301 = ~v_2298;
  assign v_2302 = v_2303 | v_2308;
  assign v_2303 = mux_2303(v_2304);
  assign v_2304 = v_2305 & 1'h1;
  assign v_2305 = v_2306 & vout_canPeek_2307;
  assign v_2306 = ~vout_canPeek_2299;
  pebbles_core
    pebbles_core_2307
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2302),
       .in0_consume_en(vin0_consume_en_2307),
       .out_canPeek(vout_canPeek_2307),
       .out_peek(vout_peek_2307));
  assign v_2308 = mux_2308(v_2309);
  assign v_2309 = ~v_2304;
  assign v_2310 = v_2311 | v_2314;
  assign v_2311 = mux_2311(v_2312);
  assign v_2312 = vout_canPeek_2313 & 1'h1;
  pebbles_core
    pebbles_core_2313
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2310),
       .in0_consume_en(vin0_consume_en_2313),
       .out_canPeek(vout_canPeek_2313),
       .out_peek(vout_peek_2313));
  assign v_2314 = mux_2314(v_2315);
  assign v_2315 = ~v_2312;
  assign v_2316 = v_2317 | v_2322;
  assign v_2317 = mux_2317(v_2318);
  assign v_2318 = v_2319 & 1'h1;
  assign v_2319 = v_2320 & vout_canPeek_2321;
  assign v_2320 = ~vout_canPeek_2313;
  pebbles_core
    pebbles_core_2321
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2316),
       .in0_consume_en(vin0_consume_en_2321),
       .out_canPeek(vout_canPeek_2321),
       .out_peek(vout_peek_2321));
  assign v_2322 = mux_2322(v_2323);
  assign v_2323 = ~v_2318;
  assign v_2324 = v_2325 | v_2328;
  assign v_2325 = mux_2325(v_2326);
  assign v_2326 = vout_canPeek_2327 & 1'h1;
  pebbles_core
    pebbles_core_2327
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2324),
       .in0_consume_en(vin0_consume_en_2327),
       .out_canPeek(vout_canPeek_2327),
       .out_peek(vout_peek_2327));
  assign v_2328 = mux_2328(v_2329);
  assign v_2329 = ~v_2326;
  assign v_2330 = v_2331 | v_2336;
  assign v_2331 = mux_2331(v_2332);
  assign v_2332 = v_2333 & 1'h1;
  assign v_2333 = v_2334 & vout_canPeek_2335;
  assign v_2334 = ~vout_canPeek_2327;
  pebbles_core
    pebbles_core_2335
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2330),
       .in0_consume_en(vin0_consume_en_2335),
       .out_canPeek(vout_canPeek_2335),
       .out_peek(vout_peek_2335));
  assign v_2336 = mux_2336(v_2337);
  assign v_2337 = ~v_2332;
  assign v_2338 = v_2339 | v_2342;
  assign v_2339 = mux_2339(v_2340);
  assign v_2340 = vout_canPeek_2341 & 1'h1;
  pebbles_core
    pebbles_core_2341
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2338),
       .in0_consume_en(vin0_consume_en_2341),
       .out_canPeek(vout_canPeek_2341),
       .out_peek(vout_peek_2341));
  assign v_2342 = mux_2342(v_2343);
  assign v_2343 = ~v_2340;
  assign v_2344 = v_2345 | v_2350;
  assign v_2345 = mux_2345(v_2346);
  assign v_2346 = v_2347 & 1'h1;
  assign v_2347 = v_2348 & vout_canPeek_2349;
  assign v_2348 = ~vout_canPeek_2341;
  pebbles_core
    pebbles_core_2349
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2344),
       .in0_consume_en(vin0_consume_en_2349),
       .out_canPeek(vout_canPeek_2349),
       .out_peek(vout_peek_2349));
  assign v_2350 = mux_2350(v_2351);
  assign v_2351 = ~v_2346;
  assign v_2352 = v_2353 | v_2356;
  assign v_2353 = mux_2353(v_2354);
  assign v_2354 = vout_canPeek_2355 & 1'h1;
  pebbles_core
    pebbles_core_2355
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2352),
       .in0_consume_en(vin0_consume_en_2355),
       .out_canPeek(vout_canPeek_2355),
       .out_peek(vout_peek_2355));
  assign v_2356 = mux_2356(v_2357);
  assign v_2357 = ~v_2354;
  assign v_2358 = v_2359 | v_2364;
  assign v_2359 = mux_2359(v_2360);
  assign v_2360 = v_2361 & 1'h1;
  assign v_2361 = v_2362 & vout_canPeek_2363;
  assign v_2362 = ~vout_canPeek_2355;
  pebbles_core
    pebbles_core_2363
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2358),
       .in0_consume_en(vin0_consume_en_2363),
       .out_canPeek(vout_canPeek_2363),
       .out_peek(vout_peek_2363));
  assign v_2364 = mux_2364(v_2365);
  assign v_2365 = ~v_2360;
  assign v_2366 = v_2367 | v_2370;
  assign v_2367 = mux_2367(v_2368);
  assign v_2368 = vout_canPeek_2369 & 1'h1;
  pebbles_core
    pebbles_core_2369
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2366),
       .in0_consume_en(vin0_consume_en_2369),
       .out_canPeek(vout_canPeek_2369),
       .out_peek(vout_peek_2369));
  assign v_2370 = mux_2370(v_2371);
  assign v_2371 = ~v_2368;
  assign v_2372 = v_2373 | v_2378;
  assign v_2373 = mux_2373(v_2374);
  assign v_2374 = v_2375 & 1'h1;
  assign v_2375 = v_2376 & vout_canPeek_2377;
  assign v_2376 = ~vout_canPeek_2369;
  pebbles_core
    pebbles_core_2377
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2372),
       .in0_consume_en(vin0_consume_en_2377),
       .out_canPeek(vout_canPeek_2377),
       .out_peek(vout_peek_2377));
  assign v_2378 = mux_2378(v_2379);
  assign v_2379 = ~v_2374;
  assign v_2380 = v_2381 | v_2384;
  assign v_2381 = mux_2381(v_2382);
  assign v_2382 = vout_canPeek_2383 & 1'h1;
  pebbles_core
    pebbles_core_2383
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2380),
       .in0_consume_en(vin0_consume_en_2383),
       .out_canPeek(vout_canPeek_2383),
       .out_peek(vout_peek_2383));
  assign v_2384 = mux_2384(v_2385);
  assign v_2385 = ~v_2382;
  assign v_2386 = v_2387 | v_2392;
  assign v_2387 = mux_2387(v_2388);
  assign v_2388 = v_2389 & 1'h1;
  assign v_2389 = v_2390 & vout_canPeek_2391;
  assign v_2390 = ~vout_canPeek_2383;
  pebbles_core
    pebbles_core_2391
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2386),
       .in0_consume_en(vin0_consume_en_2391),
       .out_canPeek(vout_canPeek_2391),
       .out_peek(vout_peek_2391));
  assign v_2392 = mux_2392(v_2393);
  assign v_2393 = ~v_2388;
  assign v_2394 = v_2395 | v_2398;
  assign v_2395 = mux_2395(v_2396);
  assign v_2396 = vout_canPeek_2397 & 1'h1;
  pebbles_core
    pebbles_core_2397
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2394),
       .in0_consume_en(vin0_consume_en_2397),
       .out_canPeek(vout_canPeek_2397),
       .out_peek(vout_peek_2397));
  assign v_2398 = mux_2398(v_2399);
  assign v_2399 = ~v_2396;
  assign v_2400 = v_2401 | v_2406;
  assign v_2401 = mux_2401(v_2402);
  assign v_2402 = v_2403 & 1'h1;
  assign v_2403 = v_2404 & vout_canPeek_2405;
  assign v_2404 = ~vout_canPeek_2397;
  pebbles_core
    pebbles_core_2405
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2400),
       .in0_consume_en(vin0_consume_en_2405),
       .out_canPeek(vout_canPeek_2405),
       .out_peek(vout_peek_2405));
  assign v_2406 = mux_2406(v_2407);
  assign v_2407 = ~v_2402;
  assign v_2408 = v_2409 | v_2412;
  assign v_2409 = mux_2409(v_2410);
  assign v_2410 = vout_canPeek_2411 & 1'h1;
  pebbles_core
    pebbles_core_2411
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2408),
       .in0_consume_en(vin0_consume_en_2411),
       .out_canPeek(vout_canPeek_2411),
       .out_peek(vout_peek_2411));
  assign v_2412 = mux_2412(v_2413);
  assign v_2413 = ~v_2410;
  assign v_2414 = v_2415 | v_2420;
  assign v_2415 = mux_2415(v_2416);
  assign v_2416 = v_2417 & 1'h1;
  assign v_2417 = v_2418 & vout_canPeek_2419;
  assign v_2418 = ~vout_canPeek_2411;
  pebbles_core
    pebbles_core_2419
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2414),
       .in0_consume_en(vin0_consume_en_2419),
       .out_canPeek(vout_canPeek_2419),
       .out_peek(vout_peek_2419));
  assign v_2420 = mux_2420(v_2421);
  assign v_2421 = ~v_2416;
  assign v_2422 = v_2423 | v_2426;
  assign v_2423 = mux_2423(v_2424);
  assign v_2424 = vout_canPeek_2425 & 1'h1;
  pebbles_core
    pebbles_core_2425
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2422),
       .in0_consume_en(vin0_consume_en_2425),
       .out_canPeek(vout_canPeek_2425),
       .out_peek(vout_peek_2425));
  assign v_2426 = mux_2426(v_2427);
  assign v_2427 = ~v_2424;
  assign v_2428 = v_2429 | v_2434;
  assign v_2429 = mux_2429(v_2430);
  assign v_2430 = v_2431 & 1'h1;
  assign v_2431 = v_2432 & vout_canPeek_2433;
  assign v_2432 = ~vout_canPeek_2425;
  pebbles_core
    pebbles_core_2433
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2428),
       .in0_consume_en(vin0_consume_en_2433),
       .out_canPeek(vout_canPeek_2433),
       .out_peek(vout_peek_2433));
  assign v_2434 = mux_2434(v_2435);
  assign v_2435 = ~v_2430;
  assign v_2436 = v_2437 | v_2440;
  assign v_2437 = mux_2437(v_2438);
  assign v_2438 = vout_canPeek_2439 & 1'h1;
  pebbles_core
    pebbles_core_2439
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2436),
       .in0_consume_en(vin0_consume_en_2439),
       .out_canPeek(vout_canPeek_2439),
       .out_peek(vout_peek_2439));
  assign v_2440 = mux_2440(v_2441);
  assign v_2441 = ~v_2438;
  assign v_2442 = v_2443 | v_2448;
  assign v_2443 = mux_2443(v_2444);
  assign v_2444 = v_2445 & 1'h1;
  assign v_2445 = v_2446 & vout_canPeek_2447;
  assign v_2446 = ~vout_canPeek_2439;
  pebbles_core
    pebbles_core_2447
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2442),
       .in0_consume_en(vin0_consume_en_2447),
       .out_canPeek(vout_canPeek_2447),
       .out_peek(vout_peek_2447));
  assign v_2448 = mux_2448(v_2449);
  assign v_2449 = ~v_2444;
  assign v_2450 = v_2451 | v_2454;
  assign v_2451 = mux_2451(v_2452);
  assign v_2452 = vout_canPeek_2453 & 1'h1;
  pebbles_core
    pebbles_core_2453
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2450),
       .in0_consume_en(vin0_consume_en_2453),
       .out_canPeek(vout_canPeek_2453),
       .out_peek(vout_peek_2453));
  assign v_2454 = mux_2454(v_2455);
  assign v_2455 = ~v_2452;
  assign v_2456 = v_2457 | v_2462;
  assign v_2457 = mux_2457(v_2458);
  assign v_2458 = v_2459 & 1'h1;
  assign v_2459 = v_2460 & vout_canPeek_2461;
  assign v_2460 = ~vout_canPeek_2453;
  pebbles_core
    pebbles_core_2461
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2456),
       .in0_consume_en(vin0_consume_en_2461),
       .out_canPeek(vout_canPeek_2461),
       .out_peek(vout_peek_2461));
  assign v_2462 = mux_2462(v_2463);
  assign v_2463 = ~v_2458;
  assign v_2464 = v_2465 | v_2468;
  assign v_2465 = mux_2465(v_2466);
  assign v_2466 = vout_canPeek_2467 & 1'h1;
  pebbles_core
    pebbles_core_2467
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2464),
       .in0_consume_en(vin0_consume_en_2467),
       .out_canPeek(vout_canPeek_2467),
       .out_peek(vout_peek_2467));
  assign v_2468 = mux_2468(v_2469);
  assign v_2469 = ~v_2466;
  assign v_2470 = v_2471 | v_2476;
  assign v_2471 = mux_2471(v_2472);
  assign v_2472 = v_2473 & 1'h1;
  assign v_2473 = v_2474 & vout_canPeek_2475;
  assign v_2474 = ~vout_canPeek_2467;
  pebbles_core
    pebbles_core_2475
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2470),
       .in0_consume_en(vin0_consume_en_2475),
       .out_canPeek(vout_canPeek_2475),
       .out_peek(vout_peek_2475));
  assign v_2476 = mux_2476(v_2477);
  assign v_2477 = ~v_2472;
  assign v_2478 = v_2479 | v_2482;
  assign v_2479 = mux_2479(v_2480);
  assign v_2480 = vout_canPeek_2481 & 1'h1;
  pebbles_core
    pebbles_core_2481
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2478),
       .in0_consume_en(vin0_consume_en_2481),
       .out_canPeek(vout_canPeek_2481),
       .out_peek(vout_peek_2481));
  assign v_2482 = mux_2482(v_2483);
  assign v_2483 = ~v_2480;
  assign v_2484 = v_2485 | v_2490;
  assign v_2485 = mux_2485(v_2486);
  assign v_2486 = v_2487 & 1'h1;
  assign v_2487 = v_2488 & vout_canPeek_2489;
  assign v_2488 = ~vout_canPeek_2481;
  pebbles_core
    pebbles_core_2489
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2484),
       .in0_consume_en(vin0_consume_en_2489),
       .out_canPeek(vout_canPeek_2489),
       .out_peek(vout_peek_2489));
  assign v_2490 = mux_2490(v_2491);
  assign v_2491 = ~v_2486;
  assign v_2492 = v_2493 | v_2496;
  assign v_2493 = mux_2493(v_2494);
  assign v_2494 = vout_canPeek_2495 & 1'h1;
  pebbles_core
    pebbles_core_2495
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2492),
       .in0_consume_en(vin0_consume_en_2495),
       .out_canPeek(vout_canPeek_2495),
       .out_peek(vout_peek_2495));
  assign v_2496 = mux_2496(v_2497);
  assign v_2497 = ~v_2494;
  assign v_2498 = v_2499 | v_2504;
  assign v_2499 = mux_2499(v_2500);
  assign v_2500 = v_2501 & 1'h1;
  assign v_2501 = v_2502 & vout_canPeek_2503;
  assign v_2502 = ~vout_canPeek_2495;
  pebbles_core
    pebbles_core_2503
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2498),
       .in0_consume_en(vin0_consume_en_2503),
       .out_canPeek(vout_canPeek_2503),
       .out_peek(vout_peek_2503));
  assign v_2504 = mux_2504(v_2505);
  assign v_2505 = ~v_2500;
  assign v_2506 = v_2507 | v_2510;
  assign v_2507 = mux_2507(v_2508);
  assign v_2508 = vout_canPeek_2509 & 1'h1;
  pebbles_core
    pebbles_core_2509
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2506),
       .in0_consume_en(vin0_consume_en_2509),
       .out_canPeek(vout_canPeek_2509),
       .out_peek(vout_peek_2509));
  assign v_2510 = mux_2510(v_2511);
  assign v_2511 = ~v_2508;
  assign v_2512 = v_2513 | v_2518;
  assign v_2513 = mux_2513(v_2514);
  assign v_2514 = v_2515 & 1'h1;
  assign v_2515 = v_2516 & vout_canPeek_2517;
  assign v_2516 = ~vout_canPeek_2509;
  pebbles_core
    pebbles_core_2517
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2512),
       .in0_consume_en(vin0_consume_en_2517),
       .out_canPeek(vout_canPeek_2517),
       .out_peek(vout_peek_2517));
  assign v_2518 = mux_2518(v_2519);
  assign v_2519 = ~v_2514;
  assign v_2520 = v_2521 | v_2524;
  assign v_2521 = mux_2521(v_2522);
  assign v_2522 = vout_canPeek_2523 & 1'h1;
  pebbles_core
    pebbles_core_2523
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2520),
       .in0_consume_en(vin0_consume_en_2523),
       .out_canPeek(vout_canPeek_2523),
       .out_peek(vout_peek_2523));
  assign v_2524 = mux_2524(v_2525);
  assign v_2525 = ~v_2522;
  assign v_2526 = v_2527 | v_2532;
  assign v_2527 = mux_2527(v_2528);
  assign v_2528 = v_2529 & 1'h1;
  assign v_2529 = v_2530 & vout_canPeek_2531;
  assign v_2530 = ~vout_canPeek_2523;
  pebbles_core
    pebbles_core_2531
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2526),
       .in0_consume_en(vin0_consume_en_2531),
       .out_canPeek(vout_canPeek_2531),
       .out_peek(vout_peek_2531));
  assign v_2532 = mux_2532(v_2533);
  assign v_2533 = ~v_2528;
  assign v_2534 = v_2535 | v_2538;
  assign v_2535 = mux_2535(v_2536);
  assign v_2536 = vout_canPeek_2537 & 1'h1;
  pebbles_core
    pebbles_core_2537
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2534),
       .in0_consume_en(vin0_consume_en_2537),
       .out_canPeek(vout_canPeek_2537),
       .out_peek(vout_peek_2537));
  assign v_2538 = mux_2538(v_2539);
  assign v_2539 = ~v_2536;
  assign v_2540 = v_2541 | v_2546;
  assign v_2541 = mux_2541(v_2542);
  assign v_2542 = v_2543 & 1'h1;
  assign v_2543 = v_2544 & vout_canPeek_2545;
  assign v_2544 = ~vout_canPeek_2537;
  pebbles_core
    pebbles_core_2545
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2540),
       .in0_consume_en(vin0_consume_en_2545),
       .out_canPeek(vout_canPeek_2545),
       .out_peek(vout_peek_2545));
  assign v_2546 = mux_2546(v_2547);
  assign v_2547 = ~v_2542;
  assign v_2548 = v_2549 | v_2552;
  assign v_2549 = mux_2549(v_2550);
  assign v_2550 = vout_canPeek_2551 & 1'h1;
  pebbles_core
    pebbles_core_2551
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2548),
       .in0_consume_en(vin0_consume_en_2551),
       .out_canPeek(vout_canPeek_2551),
       .out_peek(vout_peek_2551));
  assign v_2552 = mux_2552(v_2553);
  assign v_2553 = ~v_2550;
  assign v_2554 = v_2555 | v_2560;
  assign v_2555 = mux_2555(v_2556);
  assign v_2556 = v_2557 & 1'h1;
  assign v_2557 = v_2558 & vout_canPeek_2559;
  assign v_2558 = ~vout_canPeek_2551;
  pebbles_core
    pebbles_core_2559
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2554),
       .in0_consume_en(vin0_consume_en_2559),
       .out_canPeek(vout_canPeek_2559),
       .out_peek(vout_peek_2559));
  assign v_2560 = mux_2560(v_2561);
  assign v_2561 = ~v_2556;
  assign v_2562 = v_2563 | v_2566;
  assign v_2563 = mux_2563(v_2564);
  assign v_2564 = vout_canPeek_2565 & 1'h1;
  pebbles_core
    pebbles_core_2565
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2562),
       .in0_consume_en(vin0_consume_en_2565),
       .out_canPeek(vout_canPeek_2565),
       .out_peek(vout_peek_2565));
  assign v_2566 = mux_2566(v_2567);
  assign v_2567 = ~v_2564;
  assign v_2568 = v_2569 | v_2574;
  assign v_2569 = mux_2569(v_2570);
  assign v_2570 = v_2571 & 1'h1;
  assign v_2571 = v_2572 & vout_canPeek_2573;
  assign v_2572 = ~vout_canPeek_2565;
  pebbles_core
    pebbles_core_2573
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2568),
       .in0_consume_en(vin0_consume_en_2573),
       .out_canPeek(vout_canPeek_2573),
       .out_peek(vout_peek_2573));
  assign v_2574 = mux_2574(v_2575);
  assign v_2575 = ~v_2570;
  assign v_2576 = v_2577 | v_2580;
  assign v_2577 = mux_2577(v_2578);
  assign v_2578 = vout_canPeek_2579 & 1'h1;
  pebbles_core
    pebbles_core_2579
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2576),
       .in0_consume_en(vin0_consume_en_2579),
       .out_canPeek(vout_canPeek_2579),
       .out_peek(vout_peek_2579));
  assign v_2580 = mux_2580(v_2581);
  assign v_2581 = ~v_2578;
  assign v_2582 = v_2583 | v_2588;
  assign v_2583 = mux_2583(v_2584);
  assign v_2584 = v_2585 & 1'h1;
  assign v_2585 = v_2586 & vout_canPeek_2587;
  assign v_2586 = ~vout_canPeek_2579;
  pebbles_core
    pebbles_core_2587
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2582),
       .in0_consume_en(vin0_consume_en_2587),
       .out_canPeek(vout_canPeek_2587),
       .out_peek(vout_peek_2587));
  assign v_2588 = mux_2588(v_2589);
  assign v_2589 = ~v_2584;
  assign v_2590 = v_2591 | v_2594;
  assign v_2591 = mux_2591(v_2592);
  assign v_2592 = vout_canPeek_2593 & 1'h1;
  pebbles_core
    pebbles_core_2593
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2590),
       .in0_consume_en(vin0_consume_en_2593),
       .out_canPeek(vout_canPeek_2593),
       .out_peek(vout_peek_2593));
  assign v_2594 = mux_2594(v_2595);
  assign v_2595 = ~v_2592;
  assign v_2596 = v_2597 | v_2602;
  assign v_2597 = mux_2597(v_2598);
  assign v_2598 = v_2599 & 1'h1;
  assign v_2599 = v_2600 & vout_canPeek_2601;
  assign v_2600 = ~vout_canPeek_2593;
  pebbles_core
    pebbles_core_2601
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2596),
       .in0_consume_en(vin0_consume_en_2601),
       .out_canPeek(vout_canPeek_2601),
       .out_peek(vout_peek_2601));
  assign v_2602 = mux_2602(v_2603);
  assign v_2603 = ~v_2598;
  assign v_2604 = v_2605 | v_2608;
  assign v_2605 = mux_2605(v_2606);
  assign v_2606 = vout_canPeek_2607 & 1'h1;
  pebbles_core
    pebbles_core_2607
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2604),
       .in0_consume_en(vin0_consume_en_2607),
       .out_canPeek(vout_canPeek_2607),
       .out_peek(vout_peek_2607));
  assign v_2608 = mux_2608(v_2609);
  assign v_2609 = ~v_2606;
  assign v_2610 = v_2611 | v_2616;
  assign v_2611 = mux_2611(v_2612);
  assign v_2612 = v_2613 & 1'h1;
  assign v_2613 = v_2614 & vout_canPeek_2615;
  assign v_2614 = ~vout_canPeek_2607;
  pebbles_core
    pebbles_core_2615
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2610),
       .in0_consume_en(vin0_consume_en_2615),
       .out_canPeek(vout_canPeek_2615),
       .out_peek(vout_peek_2615));
  assign v_2616 = mux_2616(v_2617);
  assign v_2617 = ~v_2612;
  assign v_2618 = v_2619 | v_2622;
  assign v_2619 = mux_2619(v_2620);
  assign v_2620 = vout_canPeek_2621 & 1'h1;
  pebbles_core
    pebbles_core_2621
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2618),
       .in0_consume_en(vin0_consume_en_2621),
       .out_canPeek(vout_canPeek_2621),
       .out_peek(vout_peek_2621));
  assign v_2622 = mux_2622(v_2623);
  assign v_2623 = ~v_2620;
  assign v_2624 = v_2625 | v_2630;
  assign v_2625 = mux_2625(v_2626);
  assign v_2626 = v_2627 & 1'h1;
  assign v_2627 = v_2628 & vout_canPeek_2629;
  assign v_2628 = ~vout_canPeek_2621;
  pebbles_core
    pebbles_core_2629
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2624),
       .in0_consume_en(vin0_consume_en_2629),
       .out_canPeek(vout_canPeek_2629),
       .out_peek(vout_peek_2629));
  assign v_2630 = mux_2630(v_2631);
  assign v_2631 = ~v_2626;
  assign v_2632 = v_2633 | v_2636;
  assign v_2633 = mux_2633(v_2634);
  assign v_2634 = vout_canPeek_2635 & 1'h1;
  pebbles_core
    pebbles_core_2635
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2632),
       .in0_consume_en(vin0_consume_en_2635),
       .out_canPeek(vout_canPeek_2635),
       .out_peek(vout_peek_2635));
  assign v_2636 = mux_2636(v_2637);
  assign v_2637 = ~v_2634;
  assign v_2638 = v_2639 | v_2644;
  assign v_2639 = mux_2639(v_2640);
  assign v_2640 = v_2641 & 1'h1;
  assign v_2641 = v_2642 & vout_canPeek_2643;
  assign v_2642 = ~vout_canPeek_2635;
  pebbles_core
    pebbles_core_2643
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2638),
       .in0_consume_en(vin0_consume_en_2643),
       .out_canPeek(vout_canPeek_2643),
       .out_peek(vout_peek_2643));
  assign v_2644 = mux_2644(v_2645);
  assign v_2645 = ~v_2640;
  assign v_2646 = v_2647 | v_2650;
  assign v_2647 = mux_2647(v_2648);
  assign v_2648 = vout_canPeek_2649 & 1'h1;
  pebbles_core
    pebbles_core_2649
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2646),
       .in0_consume_en(vin0_consume_en_2649),
       .out_canPeek(vout_canPeek_2649),
       .out_peek(vout_peek_2649));
  assign v_2650 = mux_2650(v_2651);
  assign v_2651 = ~v_2648;
  assign v_2652 = v_2653 | v_2658;
  assign v_2653 = mux_2653(v_2654);
  assign v_2654 = v_2655 & 1'h1;
  assign v_2655 = v_2656 & vout_canPeek_2657;
  assign v_2656 = ~vout_canPeek_2649;
  pebbles_core
    pebbles_core_2657
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2652),
       .in0_consume_en(vin0_consume_en_2657),
       .out_canPeek(vout_canPeek_2657),
       .out_peek(vout_peek_2657));
  assign v_2658 = mux_2658(v_2659);
  assign v_2659 = ~v_2654;
  assign v_2660 = v_2661 | v_2664;
  assign v_2661 = mux_2661(v_2662);
  assign v_2662 = vout_canPeek_2663 & 1'h1;
  pebbles_core
    pebbles_core_2663
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2660),
       .in0_consume_en(vin0_consume_en_2663),
       .out_canPeek(vout_canPeek_2663),
       .out_peek(vout_peek_2663));
  assign v_2664 = mux_2664(v_2665);
  assign v_2665 = ~v_2662;
  assign v_2666 = v_2667 | v_2672;
  assign v_2667 = mux_2667(v_2668);
  assign v_2668 = v_2669 & 1'h1;
  assign v_2669 = v_2670 & vout_canPeek_2671;
  assign v_2670 = ~vout_canPeek_2663;
  pebbles_core
    pebbles_core_2671
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2666),
       .in0_consume_en(vin0_consume_en_2671),
       .out_canPeek(vout_canPeek_2671),
       .out_peek(vout_peek_2671));
  assign v_2672 = mux_2672(v_2673);
  assign v_2673 = ~v_2668;
  assign v_2674 = v_2675 | v_2678;
  assign v_2675 = mux_2675(v_2676);
  assign v_2676 = vout_canPeek_2677 & 1'h1;
  pebbles_core
    pebbles_core_2677
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2674),
       .in0_consume_en(vin0_consume_en_2677),
       .out_canPeek(vout_canPeek_2677),
       .out_peek(vout_peek_2677));
  assign v_2678 = mux_2678(v_2679);
  assign v_2679 = ~v_2676;
  assign v_2680 = v_2681 | v_2686;
  assign v_2681 = mux_2681(v_2682);
  assign v_2682 = v_2683 & 1'h1;
  assign v_2683 = v_2684 & vout_canPeek_2685;
  assign v_2684 = ~vout_canPeek_2677;
  pebbles_core
    pebbles_core_2685
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2680),
       .in0_consume_en(vin0_consume_en_2685),
       .out_canPeek(vout_canPeek_2685),
       .out_peek(vout_peek_2685));
  assign v_2686 = mux_2686(v_2687);
  assign v_2687 = ~v_2682;
  assign v_2688 = v_2689 | v_2692;
  assign v_2689 = mux_2689(v_2690);
  assign v_2690 = vout_canPeek_2691 & 1'h1;
  pebbles_core
    pebbles_core_2691
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2688),
       .in0_consume_en(vin0_consume_en_2691),
       .out_canPeek(vout_canPeek_2691),
       .out_peek(vout_peek_2691));
  assign v_2692 = mux_2692(v_2693);
  assign v_2693 = ~v_2690;
  assign v_2694 = v_2695 | v_2700;
  assign v_2695 = mux_2695(v_2696);
  assign v_2696 = v_2697 & 1'h1;
  assign v_2697 = v_2698 & vout_canPeek_2699;
  assign v_2698 = ~vout_canPeek_2691;
  pebbles_core
    pebbles_core_2699
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2694),
       .in0_consume_en(vin0_consume_en_2699),
       .out_canPeek(vout_canPeek_2699),
       .out_peek(vout_peek_2699));
  assign v_2700 = mux_2700(v_2701);
  assign v_2701 = ~v_2696;
  assign v_2702 = v_2703 | v_2706;
  assign v_2703 = mux_2703(v_2704);
  assign v_2704 = vout_canPeek_2705 & 1'h1;
  pebbles_core
    pebbles_core_2705
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2702),
       .in0_consume_en(vin0_consume_en_2705),
       .out_canPeek(vout_canPeek_2705),
       .out_peek(vout_peek_2705));
  assign v_2706 = mux_2706(v_2707);
  assign v_2707 = ~v_2704;
  assign v_2708 = v_2709 | v_2714;
  assign v_2709 = mux_2709(v_2710);
  assign v_2710 = v_2711 & 1'h1;
  assign v_2711 = v_2712 & vout_canPeek_2713;
  assign v_2712 = ~vout_canPeek_2705;
  pebbles_core
    pebbles_core_2713
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2708),
       .in0_consume_en(vin0_consume_en_2713),
       .out_canPeek(vout_canPeek_2713),
       .out_peek(vout_peek_2713));
  assign v_2714 = mux_2714(v_2715);
  assign v_2715 = ~v_2710;
  assign v_2716 = v_2717 | v_2720;
  assign v_2717 = mux_2717(v_2718);
  assign v_2718 = vout_canPeek_2719 & 1'h1;
  pebbles_core
    pebbles_core_2719
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2716),
       .in0_consume_en(vin0_consume_en_2719),
       .out_canPeek(vout_canPeek_2719),
       .out_peek(vout_peek_2719));
  assign v_2720 = mux_2720(v_2721);
  assign v_2721 = ~v_2718;
  assign v_2722 = v_2723 | v_2728;
  assign v_2723 = mux_2723(v_2724);
  assign v_2724 = v_2725 & 1'h1;
  assign v_2725 = v_2726 & vout_canPeek_2727;
  assign v_2726 = ~vout_canPeek_2719;
  pebbles_core
    pebbles_core_2727
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2722),
       .in0_consume_en(vin0_consume_en_2727),
       .out_canPeek(vout_canPeek_2727),
       .out_peek(vout_peek_2727));
  assign v_2728 = mux_2728(v_2729);
  assign v_2729 = ~v_2724;
  assign v_2730 = v_2731 | v_2734;
  assign v_2731 = mux_2731(v_2732);
  assign v_2732 = vout_canPeek_2733 & 1'h1;
  pebbles_core
    pebbles_core_2733
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2730),
       .in0_consume_en(vin0_consume_en_2733),
       .out_canPeek(vout_canPeek_2733),
       .out_peek(vout_peek_2733));
  assign v_2734 = mux_2734(v_2735);
  assign v_2735 = ~v_2732;
  assign v_2736 = v_2737 | v_2742;
  assign v_2737 = mux_2737(v_2738);
  assign v_2738 = v_2739 & 1'h1;
  assign v_2739 = v_2740 & vout_canPeek_2741;
  assign v_2740 = ~vout_canPeek_2733;
  pebbles_core
    pebbles_core_2741
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2736),
       .in0_consume_en(vin0_consume_en_2741),
       .out_canPeek(vout_canPeek_2741),
       .out_peek(vout_peek_2741));
  assign v_2742 = mux_2742(v_2743);
  assign v_2743 = ~v_2738;
  assign v_2744 = v_2745 | v_2748;
  assign v_2745 = mux_2745(v_2746);
  assign v_2746 = vout_canPeek_2747 & 1'h1;
  pebbles_core
    pebbles_core_2747
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2744),
       .in0_consume_en(vin0_consume_en_2747),
       .out_canPeek(vout_canPeek_2747),
       .out_peek(vout_peek_2747));
  assign v_2748 = mux_2748(v_2749);
  assign v_2749 = ~v_2746;
  assign v_2750 = v_2751 | v_2756;
  assign v_2751 = mux_2751(v_2752);
  assign v_2752 = v_2753 & 1'h1;
  assign v_2753 = v_2754 & vout_canPeek_2755;
  assign v_2754 = ~vout_canPeek_2747;
  pebbles_core
    pebbles_core_2755
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2750),
       .in0_consume_en(vin0_consume_en_2755),
       .out_canPeek(vout_canPeek_2755),
       .out_peek(vout_peek_2755));
  assign v_2756 = mux_2756(v_2757);
  assign v_2757 = ~v_2752;
  assign v_2758 = v_2759 | v_2762;
  assign v_2759 = mux_2759(v_2760);
  assign v_2760 = vout_canPeek_2761 & 1'h1;
  pebbles_core
    pebbles_core_2761
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2758),
       .in0_consume_en(vin0_consume_en_2761),
       .out_canPeek(vout_canPeek_2761),
       .out_peek(vout_peek_2761));
  assign v_2762 = mux_2762(v_2763);
  assign v_2763 = ~v_2760;
  assign v_2764 = v_2765 | v_2770;
  assign v_2765 = mux_2765(v_2766);
  assign v_2766 = v_2767 & 1'h1;
  assign v_2767 = v_2768 & vout_canPeek_2769;
  assign v_2768 = ~vout_canPeek_2761;
  pebbles_core
    pebbles_core_2769
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2764),
       .in0_consume_en(vin0_consume_en_2769),
       .out_canPeek(vout_canPeek_2769),
       .out_peek(vout_peek_2769));
  assign v_2770 = mux_2770(v_2771);
  assign v_2771 = ~v_2766;
  assign v_2772 = v_2773 | v_2776;
  assign v_2773 = mux_2773(v_2774);
  assign v_2774 = vout_canPeek_2775 & 1'h1;
  pebbles_core
    pebbles_core_2775
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2772),
       .in0_consume_en(vin0_consume_en_2775),
       .out_canPeek(vout_canPeek_2775),
       .out_peek(vout_peek_2775));
  assign v_2776 = mux_2776(v_2777);
  assign v_2777 = ~v_2774;
  assign v_2778 = v_2779 | v_2784;
  assign v_2779 = mux_2779(v_2780);
  assign v_2780 = v_2781 & 1'h1;
  assign v_2781 = v_2782 & vout_canPeek_2783;
  assign v_2782 = ~vout_canPeek_2775;
  pebbles_core
    pebbles_core_2783
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2778),
       .in0_consume_en(vin0_consume_en_2783),
       .out_canPeek(vout_canPeek_2783),
       .out_peek(vout_peek_2783));
  assign v_2784 = mux_2784(v_2785);
  assign v_2785 = ~v_2780;
  assign v_2786 = v_2787 | v_2790;
  assign v_2787 = mux_2787(v_2788);
  assign v_2788 = vout_canPeek_2789 & 1'h1;
  pebbles_core
    pebbles_core_2789
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2786),
       .in0_consume_en(vin0_consume_en_2789),
       .out_canPeek(vout_canPeek_2789),
       .out_peek(vout_peek_2789));
  assign v_2790 = mux_2790(v_2791);
  assign v_2791 = ~v_2788;
  assign v_2792 = v_2793 | v_2798;
  assign v_2793 = mux_2793(v_2794);
  assign v_2794 = v_2795 & 1'h1;
  assign v_2795 = v_2796 & vout_canPeek_2797;
  assign v_2796 = ~vout_canPeek_2789;
  pebbles_core
    pebbles_core_2797
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(1'h0),
       .in0_peek(8'bxxxxxxxx),
       .out_consume_en(v_2792),
       .in0_consume_en(vin0_consume_en_2797),
       .out_canPeek(vout_canPeek_2797),
       .out_peek(vout_peek_2797));
  assign v_2798 = mux_2798(v_2799);
  assign v_2799 = ~v_2794;
  assign in0_consume_en = v_2801;
  assign v_2801 = mux_2801(v_2802);
  assign v_2802 = ~1'h0;
  assign out_canPeek = v_2804;
  assign v_2805 = v_2806 | v_9972;
  assign v_2806 = act_2807 & 1'h1;
  assign act_2807 = v_2808 | v_5377;
  assign v_2808 = v_2809 & 1'h1;
  assign v_2809 = v_2810 & v_5384;
  assign v_2810 = ~v_2811;
  assign v_2812 = v_2813 | v_5371;
  assign v_2813 = act_2814 & 1'h1;
  assign act_2814 = v_2815 | v_3944;
  assign v_2815 = v_2816 & 1'h1;
  assign v_2816 = v_2817 & v_3951;
  assign v_2817 = ~v_2818;
  assign v_2819 = v_2820 | v_3938;
  assign v_2820 = act_2821 & 1'h1;
  assign act_2821 = v_2822 | v_3375;
  assign v_2822 = v_2823 & 1'h1;
  assign v_2823 = v_2824 & v_3382;
  assign v_2824 = ~v_2825;
  assign v_2826 = v_2827 | v_3369;
  assign v_2827 = act_2828 & 1'h1;
  assign act_2828 = v_2829 | v_3094;
  assign v_2829 = v_2830 & 1'h1;
  assign v_2830 = v_2831 & v_3101;
  assign v_2831 = ~v_2832;
  assign v_2833 = v_2834 | v_3088;
  assign v_2834 = act_2835 & 1'h1;
  assign act_2835 = v_2836 | v_2957;
  assign v_2836 = v_2837 & 1'h1;
  assign v_2837 = v_2838 & v_2964;
  assign v_2838 = ~v_2839;
  assign v_2840 = v_2841 | v_2951;
  assign v_2841 = act_2842 & 1'h1;
  assign act_2842 = v_2843 | v_2892;
  assign v_2843 = v_2844 & 1'h1;
  assign v_2844 = v_2845 & v_2899;
  assign v_2845 = ~v_2846;
  assign v_2847 = v_2848 | v_2886;
  assign v_2848 = act_2849 & 1'h1;
  assign act_2849 = v_2850 | v_2863;
  assign v_2850 = v_2851 & 1'h1;
  assign v_2851 = v_2852 & v_2870;
  assign v_2852 = ~v_2853;
  assign v_2854 = v_2855 | v_2857;
  assign v_2855 = act_2856 & 1'h1;
  assign act_2856 = v_2024 | v_2018;
  assign v_2857 = v_2858 & 1'h1;
  assign v_2858 = v_2859 & v_2860;
  assign v_2859 = ~act_2856;
  assign v_2860 = v_2861 | v_2866;
  assign v_2861 = v_2862 | v_2864;
  assign v_2862 = mux_2862(v_2863);
  assign v_2863 = v_2853 & 1'h1;
  assign v_2864 = mux_2864(v_2865);
  assign v_2865 = ~v_2863;
  assign v_2866 = ~v_2853;
  assign v_2867 = v_2868 | v_2869;
  assign v_2868 = mux_2868(v_2855);
  assign v_2869 = mux_2869(v_2857);
  assign v_2871 = v_2872 | v_2874;
  assign v_2872 = act_2873 & 1'h1;
  assign act_2873 = v_2038 | v_2032;
  assign v_2874 = v_2875 & 1'h1;
  assign v_2875 = v_2876 & v_2877;
  assign v_2876 = ~act_2873;
  assign v_2877 = v_2878 | v_2882;
  assign v_2878 = v_2879 | v_2880;
  assign v_2879 = mux_2879(v_2850);
  assign v_2880 = mux_2880(v_2881);
  assign v_2881 = ~v_2850;
  assign v_2882 = ~v_2870;
  assign v_2883 = v_2884 | v_2885;
  assign v_2884 = mux_2884(v_2872);
  assign v_2885 = mux_2885(v_2874);
  assign v_2886 = v_2887 & 1'h1;
  assign v_2887 = v_2888 & v_2889;
  assign v_2888 = ~act_2849;
  assign v_2889 = v_2890 | v_2895;
  assign v_2890 = v_2891 | v_2893;
  assign v_2891 = mux_2891(v_2892);
  assign v_2892 = v_2846 & 1'h1;
  assign v_2893 = mux_2893(v_2894);
  assign v_2894 = ~v_2892;
  assign v_2895 = ~v_2846;
  assign v_2896 = v_2897 | v_2898;
  assign v_2897 = mux_2897(v_2848);
  assign v_2898 = mux_2898(v_2886);
  assign v_2900 = v_2901 | v_2939;
  assign v_2901 = act_2902 & 1'h1;
  assign act_2902 = v_2903 | v_2916;
  assign v_2903 = v_2904 & 1'h1;
  assign v_2904 = v_2905 & v_2923;
  assign v_2905 = ~v_2906;
  assign v_2907 = v_2908 | v_2910;
  assign v_2908 = act_2909 & 1'h1;
  assign act_2909 = v_2052 | v_2046;
  assign v_2910 = v_2911 & 1'h1;
  assign v_2911 = v_2912 & v_2913;
  assign v_2912 = ~act_2909;
  assign v_2913 = v_2914 | v_2919;
  assign v_2914 = v_2915 | v_2917;
  assign v_2915 = mux_2915(v_2916);
  assign v_2916 = v_2906 & 1'h1;
  assign v_2917 = mux_2917(v_2918);
  assign v_2918 = ~v_2916;
  assign v_2919 = ~v_2906;
  assign v_2920 = v_2921 | v_2922;
  assign v_2921 = mux_2921(v_2908);
  assign v_2922 = mux_2922(v_2910);
  assign v_2924 = v_2925 | v_2927;
  assign v_2925 = act_2926 & 1'h1;
  assign act_2926 = v_2066 | v_2060;
  assign v_2927 = v_2928 & 1'h1;
  assign v_2928 = v_2929 & v_2930;
  assign v_2929 = ~act_2926;
  assign v_2930 = v_2931 | v_2935;
  assign v_2931 = v_2932 | v_2933;
  assign v_2932 = mux_2932(v_2903);
  assign v_2933 = mux_2933(v_2934);
  assign v_2934 = ~v_2903;
  assign v_2935 = ~v_2923;
  assign v_2936 = v_2937 | v_2938;
  assign v_2937 = mux_2937(v_2925);
  assign v_2938 = mux_2938(v_2927);
  assign v_2939 = v_2940 & 1'h1;
  assign v_2940 = v_2941 & v_2942;
  assign v_2941 = ~act_2902;
  assign v_2942 = v_2943 | v_2947;
  assign v_2943 = v_2944 | v_2945;
  assign v_2944 = mux_2944(v_2843);
  assign v_2945 = mux_2945(v_2946);
  assign v_2946 = ~v_2843;
  assign v_2947 = ~v_2899;
  assign v_2948 = v_2949 | v_2950;
  assign v_2949 = mux_2949(v_2901);
  assign v_2950 = mux_2950(v_2939);
  assign v_2951 = v_2952 & 1'h1;
  assign v_2952 = v_2953 & v_2954;
  assign v_2953 = ~act_2842;
  assign v_2954 = v_2955 | v_2960;
  assign v_2955 = v_2956 | v_2958;
  assign v_2956 = mux_2956(v_2957);
  assign v_2957 = v_2839 & 1'h1;
  assign v_2958 = mux_2958(v_2959);
  assign v_2959 = ~v_2957;
  assign v_2960 = ~v_2839;
  assign v_2961 = v_2962 | v_2963;
  assign v_2962 = mux_2962(v_2841);
  assign v_2963 = mux_2963(v_2951);
  assign v_2965 = v_2966 | v_3076;
  assign v_2966 = act_2967 & 1'h1;
  assign act_2967 = v_2968 | v_3017;
  assign v_2968 = v_2969 & 1'h1;
  assign v_2969 = v_2970 & v_3024;
  assign v_2970 = ~v_2971;
  assign v_2972 = v_2973 | v_3011;
  assign v_2973 = act_2974 & 1'h1;
  assign act_2974 = v_2975 | v_2988;
  assign v_2975 = v_2976 & 1'h1;
  assign v_2976 = v_2977 & v_2995;
  assign v_2977 = ~v_2978;
  assign v_2979 = v_2980 | v_2982;
  assign v_2980 = act_2981 & 1'h1;
  assign act_2981 = v_2080 | v_2074;
  assign v_2982 = v_2983 & 1'h1;
  assign v_2983 = v_2984 & v_2985;
  assign v_2984 = ~act_2981;
  assign v_2985 = v_2986 | v_2991;
  assign v_2986 = v_2987 | v_2989;
  assign v_2987 = mux_2987(v_2988);
  assign v_2988 = v_2978 & 1'h1;
  assign v_2989 = mux_2989(v_2990);
  assign v_2990 = ~v_2988;
  assign v_2991 = ~v_2978;
  assign v_2992 = v_2993 | v_2994;
  assign v_2993 = mux_2993(v_2980);
  assign v_2994 = mux_2994(v_2982);
  assign v_2996 = v_2997 | v_2999;
  assign v_2997 = act_2998 & 1'h1;
  assign act_2998 = v_2094 | v_2088;
  assign v_2999 = v_3000 & 1'h1;
  assign v_3000 = v_3001 & v_3002;
  assign v_3001 = ~act_2998;
  assign v_3002 = v_3003 | v_3007;
  assign v_3003 = v_3004 | v_3005;
  assign v_3004 = mux_3004(v_2975);
  assign v_3005 = mux_3005(v_3006);
  assign v_3006 = ~v_2975;
  assign v_3007 = ~v_2995;
  assign v_3008 = v_3009 | v_3010;
  assign v_3009 = mux_3009(v_2997);
  assign v_3010 = mux_3010(v_2999);
  assign v_3011 = v_3012 & 1'h1;
  assign v_3012 = v_3013 & v_3014;
  assign v_3013 = ~act_2974;
  assign v_3014 = v_3015 | v_3020;
  assign v_3015 = v_3016 | v_3018;
  assign v_3016 = mux_3016(v_3017);
  assign v_3017 = v_2971 & 1'h1;
  assign v_3018 = mux_3018(v_3019);
  assign v_3019 = ~v_3017;
  assign v_3020 = ~v_2971;
  assign v_3021 = v_3022 | v_3023;
  assign v_3022 = mux_3022(v_2973);
  assign v_3023 = mux_3023(v_3011);
  assign v_3025 = v_3026 | v_3064;
  assign v_3026 = act_3027 & 1'h1;
  assign act_3027 = v_3028 | v_3041;
  assign v_3028 = v_3029 & 1'h1;
  assign v_3029 = v_3030 & v_3048;
  assign v_3030 = ~v_3031;
  assign v_3032 = v_3033 | v_3035;
  assign v_3033 = act_3034 & 1'h1;
  assign act_3034 = v_2108 | v_2102;
  assign v_3035 = v_3036 & 1'h1;
  assign v_3036 = v_3037 & v_3038;
  assign v_3037 = ~act_3034;
  assign v_3038 = v_3039 | v_3044;
  assign v_3039 = v_3040 | v_3042;
  assign v_3040 = mux_3040(v_3041);
  assign v_3041 = v_3031 & 1'h1;
  assign v_3042 = mux_3042(v_3043);
  assign v_3043 = ~v_3041;
  assign v_3044 = ~v_3031;
  assign v_3045 = v_3046 | v_3047;
  assign v_3046 = mux_3046(v_3033);
  assign v_3047 = mux_3047(v_3035);
  assign v_3049 = v_3050 | v_3052;
  assign v_3050 = act_3051 & 1'h1;
  assign act_3051 = v_2122 | v_2116;
  assign v_3052 = v_3053 & 1'h1;
  assign v_3053 = v_3054 & v_3055;
  assign v_3054 = ~act_3051;
  assign v_3055 = v_3056 | v_3060;
  assign v_3056 = v_3057 | v_3058;
  assign v_3057 = mux_3057(v_3028);
  assign v_3058 = mux_3058(v_3059);
  assign v_3059 = ~v_3028;
  assign v_3060 = ~v_3048;
  assign v_3061 = v_3062 | v_3063;
  assign v_3062 = mux_3062(v_3050);
  assign v_3063 = mux_3063(v_3052);
  assign v_3064 = v_3065 & 1'h1;
  assign v_3065 = v_3066 & v_3067;
  assign v_3066 = ~act_3027;
  assign v_3067 = v_3068 | v_3072;
  assign v_3068 = v_3069 | v_3070;
  assign v_3069 = mux_3069(v_2968);
  assign v_3070 = mux_3070(v_3071);
  assign v_3071 = ~v_2968;
  assign v_3072 = ~v_3024;
  assign v_3073 = v_3074 | v_3075;
  assign v_3074 = mux_3074(v_3026);
  assign v_3075 = mux_3075(v_3064);
  assign v_3076 = v_3077 & 1'h1;
  assign v_3077 = v_3078 & v_3079;
  assign v_3078 = ~act_2967;
  assign v_3079 = v_3080 | v_3084;
  assign v_3080 = v_3081 | v_3082;
  assign v_3081 = mux_3081(v_2836);
  assign v_3082 = mux_3082(v_3083);
  assign v_3083 = ~v_2836;
  assign v_3084 = ~v_2964;
  assign v_3085 = v_3086 | v_3087;
  assign v_3086 = mux_3086(v_2966);
  assign v_3087 = mux_3087(v_3076);
  assign v_3088 = v_3089 & 1'h1;
  assign v_3089 = v_3090 & v_3091;
  assign v_3090 = ~act_2835;
  assign v_3091 = v_3092 | v_3097;
  assign v_3092 = v_3093 | v_3095;
  assign v_3093 = mux_3093(v_3094);
  assign v_3094 = v_2832 & 1'h1;
  assign v_3095 = mux_3095(v_3096);
  assign v_3096 = ~v_3094;
  assign v_3097 = ~v_2832;
  assign v_3098 = v_3099 | v_3100;
  assign v_3099 = mux_3099(v_2834);
  assign v_3100 = mux_3100(v_3088);
  assign v_3102 = v_3103 | v_3357;
  assign v_3103 = act_3104 & 1'h1;
  assign act_3104 = v_3105 | v_3226;
  assign v_3105 = v_3106 & 1'h1;
  assign v_3106 = v_3107 & v_3233;
  assign v_3107 = ~v_3108;
  assign v_3109 = v_3110 | v_3220;
  assign v_3110 = act_3111 & 1'h1;
  assign act_3111 = v_3112 | v_3161;
  assign v_3112 = v_3113 & 1'h1;
  assign v_3113 = v_3114 & v_3168;
  assign v_3114 = ~v_3115;
  assign v_3116 = v_3117 | v_3155;
  assign v_3117 = act_3118 & 1'h1;
  assign act_3118 = v_3119 | v_3132;
  assign v_3119 = v_3120 & 1'h1;
  assign v_3120 = v_3121 & v_3139;
  assign v_3121 = ~v_3122;
  assign v_3123 = v_3124 | v_3126;
  assign v_3124 = act_3125 & 1'h1;
  assign act_3125 = v_2136 | v_2130;
  assign v_3126 = v_3127 & 1'h1;
  assign v_3127 = v_3128 & v_3129;
  assign v_3128 = ~act_3125;
  assign v_3129 = v_3130 | v_3135;
  assign v_3130 = v_3131 | v_3133;
  assign v_3131 = mux_3131(v_3132);
  assign v_3132 = v_3122 & 1'h1;
  assign v_3133 = mux_3133(v_3134);
  assign v_3134 = ~v_3132;
  assign v_3135 = ~v_3122;
  assign v_3136 = v_3137 | v_3138;
  assign v_3137 = mux_3137(v_3124);
  assign v_3138 = mux_3138(v_3126);
  assign v_3140 = v_3141 | v_3143;
  assign v_3141 = act_3142 & 1'h1;
  assign act_3142 = v_2150 | v_2144;
  assign v_3143 = v_3144 & 1'h1;
  assign v_3144 = v_3145 & v_3146;
  assign v_3145 = ~act_3142;
  assign v_3146 = v_3147 | v_3151;
  assign v_3147 = v_3148 | v_3149;
  assign v_3148 = mux_3148(v_3119);
  assign v_3149 = mux_3149(v_3150);
  assign v_3150 = ~v_3119;
  assign v_3151 = ~v_3139;
  assign v_3152 = v_3153 | v_3154;
  assign v_3153 = mux_3153(v_3141);
  assign v_3154 = mux_3154(v_3143);
  assign v_3155 = v_3156 & 1'h1;
  assign v_3156 = v_3157 & v_3158;
  assign v_3157 = ~act_3118;
  assign v_3158 = v_3159 | v_3164;
  assign v_3159 = v_3160 | v_3162;
  assign v_3160 = mux_3160(v_3161);
  assign v_3161 = v_3115 & 1'h1;
  assign v_3162 = mux_3162(v_3163);
  assign v_3163 = ~v_3161;
  assign v_3164 = ~v_3115;
  assign v_3165 = v_3166 | v_3167;
  assign v_3166 = mux_3166(v_3117);
  assign v_3167 = mux_3167(v_3155);
  assign v_3169 = v_3170 | v_3208;
  assign v_3170 = act_3171 & 1'h1;
  assign act_3171 = v_3172 | v_3185;
  assign v_3172 = v_3173 & 1'h1;
  assign v_3173 = v_3174 & v_3192;
  assign v_3174 = ~v_3175;
  assign v_3176 = v_3177 | v_3179;
  assign v_3177 = act_3178 & 1'h1;
  assign act_3178 = v_2164 | v_2158;
  assign v_3179 = v_3180 & 1'h1;
  assign v_3180 = v_3181 & v_3182;
  assign v_3181 = ~act_3178;
  assign v_3182 = v_3183 | v_3188;
  assign v_3183 = v_3184 | v_3186;
  assign v_3184 = mux_3184(v_3185);
  assign v_3185 = v_3175 & 1'h1;
  assign v_3186 = mux_3186(v_3187);
  assign v_3187 = ~v_3185;
  assign v_3188 = ~v_3175;
  assign v_3189 = v_3190 | v_3191;
  assign v_3190 = mux_3190(v_3177);
  assign v_3191 = mux_3191(v_3179);
  assign v_3193 = v_3194 | v_3196;
  assign v_3194 = act_3195 & 1'h1;
  assign act_3195 = v_2178 | v_2172;
  assign v_3196 = v_3197 & 1'h1;
  assign v_3197 = v_3198 & v_3199;
  assign v_3198 = ~act_3195;
  assign v_3199 = v_3200 | v_3204;
  assign v_3200 = v_3201 | v_3202;
  assign v_3201 = mux_3201(v_3172);
  assign v_3202 = mux_3202(v_3203);
  assign v_3203 = ~v_3172;
  assign v_3204 = ~v_3192;
  assign v_3205 = v_3206 | v_3207;
  assign v_3206 = mux_3206(v_3194);
  assign v_3207 = mux_3207(v_3196);
  assign v_3208 = v_3209 & 1'h1;
  assign v_3209 = v_3210 & v_3211;
  assign v_3210 = ~act_3171;
  assign v_3211 = v_3212 | v_3216;
  assign v_3212 = v_3213 | v_3214;
  assign v_3213 = mux_3213(v_3112);
  assign v_3214 = mux_3214(v_3215);
  assign v_3215 = ~v_3112;
  assign v_3216 = ~v_3168;
  assign v_3217 = v_3218 | v_3219;
  assign v_3218 = mux_3218(v_3170);
  assign v_3219 = mux_3219(v_3208);
  assign v_3220 = v_3221 & 1'h1;
  assign v_3221 = v_3222 & v_3223;
  assign v_3222 = ~act_3111;
  assign v_3223 = v_3224 | v_3229;
  assign v_3224 = v_3225 | v_3227;
  assign v_3225 = mux_3225(v_3226);
  assign v_3226 = v_3108 & 1'h1;
  assign v_3227 = mux_3227(v_3228);
  assign v_3228 = ~v_3226;
  assign v_3229 = ~v_3108;
  assign v_3230 = v_3231 | v_3232;
  assign v_3231 = mux_3231(v_3110);
  assign v_3232 = mux_3232(v_3220);
  assign v_3234 = v_3235 | v_3345;
  assign v_3235 = act_3236 & 1'h1;
  assign act_3236 = v_3237 | v_3286;
  assign v_3237 = v_3238 & 1'h1;
  assign v_3238 = v_3239 & v_3293;
  assign v_3239 = ~v_3240;
  assign v_3241 = v_3242 | v_3280;
  assign v_3242 = act_3243 & 1'h1;
  assign act_3243 = v_3244 | v_3257;
  assign v_3244 = v_3245 & 1'h1;
  assign v_3245 = v_3246 & v_3264;
  assign v_3246 = ~v_3247;
  assign v_3248 = v_3249 | v_3251;
  assign v_3249 = act_3250 & 1'h1;
  assign act_3250 = v_2192 | v_2186;
  assign v_3251 = v_3252 & 1'h1;
  assign v_3252 = v_3253 & v_3254;
  assign v_3253 = ~act_3250;
  assign v_3254 = v_3255 | v_3260;
  assign v_3255 = v_3256 | v_3258;
  assign v_3256 = mux_3256(v_3257);
  assign v_3257 = v_3247 & 1'h1;
  assign v_3258 = mux_3258(v_3259);
  assign v_3259 = ~v_3257;
  assign v_3260 = ~v_3247;
  assign v_3261 = v_3262 | v_3263;
  assign v_3262 = mux_3262(v_3249);
  assign v_3263 = mux_3263(v_3251);
  assign v_3265 = v_3266 | v_3268;
  assign v_3266 = act_3267 & 1'h1;
  assign act_3267 = v_2206 | v_2200;
  assign v_3268 = v_3269 & 1'h1;
  assign v_3269 = v_3270 & v_3271;
  assign v_3270 = ~act_3267;
  assign v_3271 = v_3272 | v_3276;
  assign v_3272 = v_3273 | v_3274;
  assign v_3273 = mux_3273(v_3244);
  assign v_3274 = mux_3274(v_3275);
  assign v_3275 = ~v_3244;
  assign v_3276 = ~v_3264;
  assign v_3277 = v_3278 | v_3279;
  assign v_3278 = mux_3278(v_3266);
  assign v_3279 = mux_3279(v_3268);
  assign v_3280 = v_3281 & 1'h1;
  assign v_3281 = v_3282 & v_3283;
  assign v_3282 = ~act_3243;
  assign v_3283 = v_3284 | v_3289;
  assign v_3284 = v_3285 | v_3287;
  assign v_3285 = mux_3285(v_3286);
  assign v_3286 = v_3240 & 1'h1;
  assign v_3287 = mux_3287(v_3288);
  assign v_3288 = ~v_3286;
  assign v_3289 = ~v_3240;
  assign v_3290 = v_3291 | v_3292;
  assign v_3291 = mux_3291(v_3242);
  assign v_3292 = mux_3292(v_3280);
  assign v_3294 = v_3295 | v_3333;
  assign v_3295 = act_3296 & 1'h1;
  assign act_3296 = v_3297 | v_3310;
  assign v_3297 = v_3298 & 1'h1;
  assign v_3298 = v_3299 & v_3317;
  assign v_3299 = ~v_3300;
  assign v_3301 = v_3302 | v_3304;
  assign v_3302 = act_3303 & 1'h1;
  assign act_3303 = v_2220 | v_2214;
  assign v_3304 = v_3305 & 1'h1;
  assign v_3305 = v_3306 & v_3307;
  assign v_3306 = ~act_3303;
  assign v_3307 = v_3308 | v_3313;
  assign v_3308 = v_3309 | v_3311;
  assign v_3309 = mux_3309(v_3310);
  assign v_3310 = v_3300 & 1'h1;
  assign v_3311 = mux_3311(v_3312);
  assign v_3312 = ~v_3310;
  assign v_3313 = ~v_3300;
  assign v_3314 = v_3315 | v_3316;
  assign v_3315 = mux_3315(v_3302);
  assign v_3316 = mux_3316(v_3304);
  assign v_3318 = v_3319 | v_3321;
  assign v_3319 = act_3320 & 1'h1;
  assign act_3320 = v_2234 | v_2228;
  assign v_3321 = v_3322 & 1'h1;
  assign v_3322 = v_3323 & v_3324;
  assign v_3323 = ~act_3320;
  assign v_3324 = v_3325 | v_3329;
  assign v_3325 = v_3326 | v_3327;
  assign v_3326 = mux_3326(v_3297);
  assign v_3327 = mux_3327(v_3328);
  assign v_3328 = ~v_3297;
  assign v_3329 = ~v_3317;
  assign v_3330 = v_3331 | v_3332;
  assign v_3331 = mux_3331(v_3319);
  assign v_3332 = mux_3332(v_3321);
  assign v_3333 = v_3334 & 1'h1;
  assign v_3334 = v_3335 & v_3336;
  assign v_3335 = ~act_3296;
  assign v_3336 = v_3337 | v_3341;
  assign v_3337 = v_3338 | v_3339;
  assign v_3338 = mux_3338(v_3237);
  assign v_3339 = mux_3339(v_3340);
  assign v_3340 = ~v_3237;
  assign v_3341 = ~v_3293;
  assign v_3342 = v_3343 | v_3344;
  assign v_3343 = mux_3343(v_3295);
  assign v_3344 = mux_3344(v_3333);
  assign v_3345 = v_3346 & 1'h1;
  assign v_3346 = v_3347 & v_3348;
  assign v_3347 = ~act_3236;
  assign v_3348 = v_3349 | v_3353;
  assign v_3349 = v_3350 | v_3351;
  assign v_3350 = mux_3350(v_3105);
  assign v_3351 = mux_3351(v_3352);
  assign v_3352 = ~v_3105;
  assign v_3353 = ~v_3233;
  assign v_3354 = v_3355 | v_3356;
  assign v_3355 = mux_3355(v_3235);
  assign v_3356 = mux_3356(v_3345);
  assign v_3357 = v_3358 & 1'h1;
  assign v_3358 = v_3359 & v_3360;
  assign v_3359 = ~act_3104;
  assign v_3360 = v_3361 | v_3365;
  assign v_3361 = v_3362 | v_3363;
  assign v_3362 = mux_3362(v_2829);
  assign v_3363 = mux_3363(v_3364);
  assign v_3364 = ~v_2829;
  assign v_3365 = ~v_3101;
  assign v_3366 = v_3367 | v_3368;
  assign v_3367 = mux_3367(v_3103);
  assign v_3368 = mux_3368(v_3357);
  assign v_3369 = v_3370 & 1'h1;
  assign v_3370 = v_3371 & v_3372;
  assign v_3371 = ~act_2828;
  assign v_3372 = v_3373 | v_3378;
  assign v_3373 = v_3374 | v_3376;
  assign v_3374 = mux_3374(v_3375);
  assign v_3375 = v_2825 & 1'h1;
  assign v_3376 = mux_3376(v_3377);
  assign v_3377 = ~v_3375;
  assign v_3378 = ~v_2825;
  assign v_3379 = v_3380 | v_3381;
  assign v_3380 = mux_3380(v_2827);
  assign v_3381 = mux_3381(v_3369);
  assign v_3383 = v_3384 | v_3926;
  assign v_3384 = act_3385 & 1'h1;
  assign act_3385 = v_3386 | v_3651;
  assign v_3386 = v_3387 & 1'h1;
  assign v_3387 = v_3388 & v_3658;
  assign v_3388 = ~v_3389;
  assign v_3390 = v_3391 | v_3645;
  assign v_3391 = act_3392 & 1'h1;
  assign act_3392 = v_3393 | v_3514;
  assign v_3393 = v_3394 & 1'h1;
  assign v_3394 = v_3395 & v_3521;
  assign v_3395 = ~v_3396;
  assign v_3397 = v_3398 | v_3508;
  assign v_3398 = act_3399 & 1'h1;
  assign act_3399 = v_3400 | v_3449;
  assign v_3400 = v_3401 & 1'h1;
  assign v_3401 = v_3402 & v_3456;
  assign v_3402 = ~v_3403;
  assign v_3404 = v_3405 | v_3443;
  assign v_3405 = act_3406 & 1'h1;
  assign act_3406 = v_3407 | v_3420;
  assign v_3407 = v_3408 & 1'h1;
  assign v_3408 = v_3409 & v_3427;
  assign v_3409 = ~v_3410;
  assign v_3411 = v_3412 | v_3414;
  assign v_3412 = act_3413 & 1'h1;
  assign act_3413 = v_2248 | v_2242;
  assign v_3414 = v_3415 & 1'h1;
  assign v_3415 = v_3416 & v_3417;
  assign v_3416 = ~act_3413;
  assign v_3417 = v_3418 | v_3423;
  assign v_3418 = v_3419 | v_3421;
  assign v_3419 = mux_3419(v_3420);
  assign v_3420 = v_3410 & 1'h1;
  assign v_3421 = mux_3421(v_3422);
  assign v_3422 = ~v_3420;
  assign v_3423 = ~v_3410;
  assign v_3424 = v_3425 | v_3426;
  assign v_3425 = mux_3425(v_3412);
  assign v_3426 = mux_3426(v_3414);
  assign v_3428 = v_3429 | v_3431;
  assign v_3429 = act_3430 & 1'h1;
  assign act_3430 = v_2262 | v_2256;
  assign v_3431 = v_3432 & 1'h1;
  assign v_3432 = v_3433 & v_3434;
  assign v_3433 = ~act_3430;
  assign v_3434 = v_3435 | v_3439;
  assign v_3435 = v_3436 | v_3437;
  assign v_3436 = mux_3436(v_3407);
  assign v_3437 = mux_3437(v_3438);
  assign v_3438 = ~v_3407;
  assign v_3439 = ~v_3427;
  assign v_3440 = v_3441 | v_3442;
  assign v_3441 = mux_3441(v_3429);
  assign v_3442 = mux_3442(v_3431);
  assign v_3443 = v_3444 & 1'h1;
  assign v_3444 = v_3445 & v_3446;
  assign v_3445 = ~act_3406;
  assign v_3446 = v_3447 | v_3452;
  assign v_3447 = v_3448 | v_3450;
  assign v_3448 = mux_3448(v_3449);
  assign v_3449 = v_3403 & 1'h1;
  assign v_3450 = mux_3450(v_3451);
  assign v_3451 = ~v_3449;
  assign v_3452 = ~v_3403;
  assign v_3453 = v_3454 | v_3455;
  assign v_3454 = mux_3454(v_3405);
  assign v_3455 = mux_3455(v_3443);
  assign v_3457 = v_3458 | v_3496;
  assign v_3458 = act_3459 & 1'h1;
  assign act_3459 = v_3460 | v_3473;
  assign v_3460 = v_3461 & 1'h1;
  assign v_3461 = v_3462 & v_3480;
  assign v_3462 = ~v_3463;
  assign v_3464 = v_3465 | v_3467;
  assign v_3465 = act_3466 & 1'h1;
  assign act_3466 = v_2276 | v_2270;
  assign v_3467 = v_3468 & 1'h1;
  assign v_3468 = v_3469 & v_3470;
  assign v_3469 = ~act_3466;
  assign v_3470 = v_3471 | v_3476;
  assign v_3471 = v_3472 | v_3474;
  assign v_3472 = mux_3472(v_3473);
  assign v_3473 = v_3463 & 1'h1;
  assign v_3474 = mux_3474(v_3475);
  assign v_3475 = ~v_3473;
  assign v_3476 = ~v_3463;
  assign v_3477 = v_3478 | v_3479;
  assign v_3478 = mux_3478(v_3465);
  assign v_3479 = mux_3479(v_3467);
  assign v_3481 = v_3482 | v_3484;
  assign v_3482 = act_3483 & 1'h1;
  assign act_3483 = v_2290 | v_2284;
  assign v_3484 = v_3485 & 1'h1;
  assign v_3485 = v_3486 & v_3487;
  assign v_3486 = ~act_3483;
  assign v_3487 = v_3488 | v_3492;
  assign v_3488 = v_3489 | v_3490;
  assign v_3489 = mux_3489(v_3460);
  assign v_3490 = mux_3490(v_3491);
  assign v_3491 = ~v_3460;
  assign v_3492 = ~v_3480;
  assign v_3493 = v_3494 | v_3495;
  assign v_3494 = mux_3494(v_3482);
  assign v_3495 = mux_3495(v_3484);
  assign v_3496 = v_3497 & 1'h1;
  assign v_3497 = v_3498 & v_3499;
  assign v_3498 = ~act_3459;
  assign v_3499 = v_3500 | v_3504;
  assign v_3500 = v_3501 | v_3502;
  assign v_3501 = mux_3501(v_3400);
  assign v_3502 = mux_3502(v_3503);
  assign v_3503 = ~v_3400;
  assign v_3504 = ~v_3456;
  assign v_3505 = v_3506 | v_3507;
  assign v_3506 = mux_3506(v_3458);
  assign v_3507 = mux_3507(v_3496);
  assign v_3508 = v_3509 & 1'h1;
  assign v_3509 = v_3510 & v_3511;
  assign v_3510 = ~act_3399;
  assign v_3511 = v_3512 | v_3517;
  assign v_3512 = v_3513 | v_3515;
  assign v_3513 = mux_3513(v_3514);
  assign v_3514 = v_3396 & 1'h1;
  assign v_3515 = mux_3515(v_3516);
  assign v_3516 = ~v_3514;
  assign v_3517 = ~v_3396;
  assign v_3518 = v_3519 | v_3520;
  assign v_3519 = mux_3519(v_3398);
  assign v_3520 = mux_3520(v_3508);
  assign v_3522 = v_3523 | v_3633;
  assign v_3523 = act_3524 & 1'h1;
  assign act_3524 = v_3525 | v_3574;
  assign v_3525 = v_3526 & 1'h1;
  assign v_3526 = v_3527 & v_3581;
  assign v_3527 = ~v_3528;
  assign v_3529 = v_3530 | v_3568;
  assign v_3530 = act_3531 & 1'h1;
  assign act_3531 = v_3532 | v_3545;
  assign v_3532 = v_3533 & 1'h1;
  assign v_3533 = v_3534 & v_3552;
  assign v_3534 = ~v_3535;
  assign v_3536 = v_3537 | v_3539;
  assign v_3537 = act_3538 & 1'h1;
  assign act_3538 = v_2304 | v_2298;
  assign v_3539 = v_3540 & 1'h1;
  assign v_3540 = v_3541 & v_3542;
  assign v_3541 = ~act_3538;
  assign v_3542 = v_3543 | v_3548;
  assign v_3543 = v_3544 | v_3546;
  assign v_3544 = mux_3544(v_3545);
  assign v_3545 = v_3535 & 1'h1;
  assign v_3546 = mux_3546(v_3547);
  assign v_3547 = ~v_3545;
  assign v_3548 = ~v_3535;
  assign v_3549 = v_3550 | v_3551;
  assign v_3550 = mux_3550(v_3537);
  assign v_3551 = mux_3551(v_3539);
  assign v_3553 = v_3554 | v_3556;
  assign v_3554 = act_3555 & 1'h1;
  assign act_3555 = v_2318 | v_2312;
  assign v_3556 = v_3557 & 1'h1;
  assign v_3557 = v_3558 & v_3559;
  assign v_3558 = ~act_3555;
  assign v_3559 = v_3560 | v_3564;
  assign v_3560 = v_3561 | v_3562;
  assign v_3561 = mux_3561(v_3532);
  assign v_3562 = mux_3562(v_3563);
  assign v_3563 = ~v_3532;
  assign v_3564 = ~v_3552;
  assign v_3565 = v_3566 | v_3567;
  assign v_3566 = mux_3566(v_3554);
  assign v_3567 = mux_3567(v_3556);
  assign v_3568 = v_3569 & 1'h1;
  assign v_3569 = v_3570 & v_3571;
  assign v_3570 = ~act_3531;
  assign v_3571 = v_3572 | v_3577;
  assign v_3572 = v_3573 | v_3575;
  assign v_3573 = mux_3573(v_3574);
  assign v_3574 = v_3528 & 1'h1;
  assign v_3575 = mux_3575(v_3576);
  assign v_3576 = ~v_3574;
  assign v_3577 = ~v_3528;
  assign v_3578 = v_3579 | v_3580;
  assign v_3579 = mux_3579(v_3530);
  assign v_3580 = mux_3580(v_3568);
  assign v_3582 = v_3583 | v_3621;
  assign v_3583 = act_3584 & 1'h1;
  assign act_3584 = v_3585 | v_3598;
  assign v_3585 = v_3586 & 1'h1;
  assign v_3586 = v_3587 & v_3605;
  assign v_3587 = ~v_3588;
  assign v_3589 = v_3590 | v_3592;
  assign v_3590 = act_3591 & 1'h1;
  assign act_3591 = v_2332 | v_2326;
  assign v_3592 = v_3593 & 1'h1;
  assign v_3593 = v_3594 & v_3595;
  assign v_3594 = ~act_3591;
  assign v_3595 = v_3596 | v_3601;
  assign v_3596 = v_3597 | v_3599;
  assign v_3597 = mux_3597(v_3598);
  assign v_3598 = v_3588 & 1'h1;
  assign v_3599 = mux_3599(v_3600);
  assign v_3600 = ~v_3598;
  assign v_3601 = ~v_3588;
  assign v_3602 = v_3603 | v_3604;
  assign v_3603 = mux_3603(v_3590);
  assign v_3604 = mux_3604(v_3592);
  assign v_3606 = v_3607 | v_3609;
  assign v_3607 = act_3608 & 1'h1;
  assign act_3608 = v_2346 | v_2340;
  assign v_3609 = v_3610 & 1'h1;
  assign v_3610 = v_3611 & v_3612;
  assign v_3611 = ~act_3608;
  assign v_3612 = v_3613 | v_3617;
  assign v_3613 = v_3614 | v_3615;
  assign v_3614 = mux_3614(v_3585);
  assign v_3615 = mux_3615(v_3616);
  assign v_3616 = ~v_3585;
  assign v_3617 = ~v_3605;
  assign v_3618 = v_3619 | v_3620;
  assign v_3619 = mux_3619(v_3607);
  assign v_3620 = mux_3620(v_3609);
  assign v_3621 = v_3622 & 1'h1;
  assign v_3622 = v_3623 & v_3624;
  assign v_3623 = ~act_3584;
  assign v_3624 = v_3625 | v_3629;
  assign v_3625 = v_3626 | v_3627;
  assign v_3626 = mux_3626(v_3525);
  assign v_3627 = mux_3627(v_3628);
  assign v_3628 = ~v_3525;
  assign v_3629 = ~v_3581;
  assign v_3630 = v_3631 | v_3632;
  assign v_3631 = mux_3631(v_3583);
  assign v_3632 = mux_3632(v_3621);
  assign v_3633 = v_3634 & 1'h1;
  assign v_3634 = v_3635 & v_3636;
  assign v_3635 = ~act_3524;
  assign v_3636 = v_3637 | v_3641;
  assign v_3637 = v_3638 | v_3639;
  assign v_3638 = mux_3638(v_3393);
  assign v_3639 = mux_3639(v_3640);
  assign v_3640 = ~v_3393;
  assign v_3641 = ~v_3521;
  assign v_3642 = v_3643 | v_3644;
  assign v_3643 = mux_3643(v_3523);
  assign v_3644 = mux_3644(v_3633);
  assign v_3645 = v_3646 & 1'h1;
  assign v_3646 = v_3647 & v_3648;
  assign v_3647 = ~act_3392;
  assign v_3648 = v_3649 | v_3654;
  assign v_3649 = v_3650 | v_3652;
  assign v_3650 = mux_3650(v_3651);
  assign v_3651 = v_3389 & 1'h1;
  assign v_3652 = mux_3652(v_3653);
  assign v_3653 = ~v_3651;
  assign v_3654 = ~v_3389;
  assign v_3655 = v_3656 | v_3657;
  assign v_3656 = mux_3656(v_3391);
  assign v_3657 = mux_3657(v_3645);
  assign v_3659 = v_3660 | v_3914;
  assign v_3660 = act_3661 & 1'h1;
  assign act_3661 = v_3662 | v_3783;
  assign v_3662 = v_3663 & 1'h1;
  assign v_3663 = v_3664 & v_3790;
  assign v_3664 = ~v_3665;
  assign v_3666 = v_3667 | v_3777;
  assign v_3667 = act_3668 & 1'h1;
  assign act_3668 = v_3669 | v_3718;
  assign v_3669 = v_3670 & 1'h1;
  assign v_3670 = v_3671 & v_3725;
  assign v_3671 = ~v_3672;
  assign v_3673 = v_3674 | v_3712;
  assign v_3674 = act_3675 & 1'h1;
  assign act_3675 = v_3676 | v_3689;
  assign v_3676 = v_3677 & 1'h1;
  assign v_3677 = v_3678 & v_3696;
  assign v_3678 = ~v_3679;
  assign v_3680 = v_3681 | v_3683;
  assign v_3681 = act_3682 & 1'h1;
  assign act_3682 = v_2360 | v_2354;
  assign v_3683 = v_3684 & 1'h1;
  assign v_3684 = v_3685 & v_3686;
  assign v_3685 = ~act_3682;
  assign v_3686 = v_3687 | v_3692;
  assign v_3687 = v_3688 | v_3690;
  assign v_3688 = mux_3688(v_3689);
  assign v_3689 = v_3679 & 1'h1;
  assign v_3690 = mux_3690(v_3691);
  assign v_3691 = ~v_3689;
  assign v_3692 = ~v_3679;
  assign v_3693 = v_3694 | v_3695;
  assign v_3694 = mux_3694(v_3681);
  assign v_3695 = mux_3695(v_3683);
  assign v_3697 = v_3698 | v_3700;
  assign v_3698 = act_3699 & 1'h1;
  assign act_3699 = v_2374 | v_2368;
  assign v_3700 = v_3701 & 1'h1;
  assign v_3701 = v_3702 & v_3703;
  assign v_3702 = ~act_3699;
  assign v_3703 = v_3704 | v_3708;
  assign v_3704 = v_3705 | v_3706;
  assign v_3705 = mux_3705(v_3676);
  assign v_3706 = mux_3706(v_3707);
  assign v_3707 = ~v_3676;
  assign v_3708 = ~v_3696;
  assign v_3709 = v_3710 | v_3711;
  assign v_3710 = mux_3710(v_3698);
  assign v_3711 = mux_3711(v_3700);
  assign v_3712 = v_3713 & 1'h1;
  assign v_3713 = v_3714 & v_3715;
  assign v_3714 = ~act_3675;
  assign v_3715 = v_3716 | v_3721;
  assign v_3716 = v_3717 | v_3719;
  assign v_3717 = mux_3717(v_3718);
  assign v_3718 = v_3672 & 1'h1;
  assign v_3719 = mux_3719(v_3720);
  assign v_3720 = ~v_3718;
  assign v_3721 = ~v_3672;
  assign v_3722 = v_3723 | v_3724;
  assign v_3723 = mux_3723(v_3674);
  assign v_3724 = mux_3724(v_3712);
  assign v_3726 = v_3727 | v_3765;
  assign v_3727 = act_3728 & 1'h1;
  assign act_3728 = v_3729 | v_3742;
  assign v_3729 = v_3730 & 1'h1;
  assign v_3730 = v_3731 & v_3749;
  assign v_3731 = ~v_3732;
  assign v_3733 = v_3734 | v_3736;
  assign v_3734 = act_3735 & 1'h1;
  assign act_3735 = v_2388 | v_2382;
  assign v_3736 = v_3737 & 1'h1;
  assign v_3737 = v_3738 & v_3739;
  assign v_3738 = ~act_3735;
  assign v_3739 = v_3740 | v_3745;
  assign v_3740 = v_3741 | v_3743;
  assign v_3741 = mux_3741(v_3742);
  assign v_3742 = v_3732 & 1'h1;
  assign v_3743 = mux_3743(v_3744);
  assign v_3744 = ~v_3742;
  assign v_3745 = ~v_3732;
  assign v_3746 = v_3747 | v_3748;
  assign v_3747 = mux_3747(v_3734);
  assign v_3748 = mux_3748(v_3736);
  assign v_3750 = v_3751 | v_3753;
  assign v_3751 = act_3752 & 1'h1;
  assign act_3752 = v_2402 | v_2396;
  assign v_3753 = v_3754 & 1'h1;
  assign v_3754 = v_3755 & v_3756;
  assign v_3755 = ~act_3752;
  assign v_3756 = v_3757 | v_3761;
  assign v_3757 = v_3758 | v_3759;
  assign v_3758 = mux_3758(v_3729);
  assign v_3759 = mux_3759(v_3760);
  assign v_3760 = ~v_3729;
  assign v_3761 = ~v_3749;
  assign v_3762 = v_3763 | v_3764;
  assign v_3763 = mux_3763(v_3751);
  assign v_3764 = mux_3764(v_3753);
  assign v_3765 = v_3766 & 1'h1;
  assign v_3766 = v_3767 & v_3768;
  assign v_3767 = ~act_3728;
  assign v_3768 = v_3769 | v_3773;
  assign v_3769 = v_3770 | v_3771;
  assign v_3770 = mux_3770(v_3669);
  assign v_3771 = mux_3771(v_3772);
  assign v_3772 = ~v_3669;
  assign v_3773 = ~v_3725;
  assign v_3774 = v_3775 | v_3776;
  assign v_3775 = mux_3775(v_3727);
  assign v_3776 = mux_3776(v_3765);
  assign v_3777 = v_3778 & 1'h1;
  assign v_3778 = v_3779 & v_3780;
  assign v_3779 = ~act_3668;
  assign v_3780 = v_3781 | v_3786;
  assign v_3781 = v_3782 | v_3784;
  assign v_3782 = mux_3782(v_3783);
  assign v_3783 = v_3665 & 1'h1;
  assign v_3784 = mux_3784(v_3785);
  assign v_3785 = ~v_3783;
  assign v_3786 = ~v_3665;
  assign v_3787 = v_3788 | v_3789;
  assign v_3788 = mux_3788(v_3667);
  assign v_3789 = mux_3789(v_3777);
  assign v_3791 = v_3792 | v_3902;
  assign v_3792 = act_3793 & 1'h1;
  assign act_3793 = v_3794 | v_3843;
  assign v_3794 = v_3795 & 1'h1;
  assign v_3795 = v_3796 & v_3850;
  assign v_3796 = ~v_3797;
  assign v_3798 = v_3799 | v_3837;
  assign v_3799 = act_3800 & 1'h1;
  assign act_3800 = v_3801 | v_3814;
  assign v_3801 = v_3802 & 1'h1;
  assign v_3802 = v_3803 & v_3821;
  assign v_3803 = ~v_3804;
  assign v_3805 = v_3806 | v_3808;
  assign v_3806 = act_3807 & 1'h1;
  assign act_3807 = v_2416 | v_2410;
  assign v_3808 = v_3809 & 1'h1;
  assign v_3809 = v_3810 & v_3811;
  assign v_3810 = ~act_3807;
  assign v_3811 = v_3812 | v_3817;
  assign v_3812 = v_3813 | v_3815;
  assign v_3813 = mux_3813(v_3814);
  assign v_3814 = v_3804 & 1'h1;
  assign v_3815 = mux_3815(v_3816);
  assign v_3816 = ~v_3814;
  assign v_3817 = ~v_3804;
  assign v_3818 = v_3819 | v_3820;
  assign v_3819 = mux_3819(v_3806);
  assign v_3820 = mux_3820(v_3808);
  assign v_3822 = v_3823 | v_3825;
  assign v_3823 = act_3824 & 1'h1;
  assign act_3824 = v_2430 | v_2424;
  assign v_3825 = v_3826 & 1'h1;
  assign v_3826 = v_3827 & v_3828;
  assign v_3827 = ~act_3824;
  assign v_3828 = v_3829 | v_3833;
  assign v_3829 = v_3830 | v_3831;
  assign v_3830 = mux_3830(v_3801);
  assign v_3831 = mux_3831(v_3832);
  assign v_3832 = ~v_3801;
  assign v_3833 = ~v_3821;
  assign v_3834 = v_3835 | v_3836;
  assign v_3835 = mux_3835(v_3823);
  assign v_3836 = mux_3836(v_3825);
  assign v_3837 = v_3838 & 1'h1;
  assign v_3838 = v_3839 & v_3840;
  assign v_3839 = ~act_3800;
  assign v_3840 = v_3841 | v_3846;
  assign v_3841 = v_3842 | v_3844;
  assign v_3842 = mux_3842(v_3843);
  assign v_3843 = v_3797 & 1'h1;
  assign v_3844 = mux_3844(v_3845);
  assign v_3845 = ~v_3843;
  assign v_3846 = ~v_3797;
  assign v_3847 = v_3848 | v_3849;
  assign v_3848 = mux_3848(v_3799);
  assign v_3849 = mux_3849(v_3837);
  assign v_3851 = v_3852 | v_3890;
  assign v_3852 = act_3853 & 1'h1;
  assign act_3853 = v_3854 | v_3867;
  assign v_3854 = v_3855 & 1'h1;
  assign v_3855 = v_3856 & v_3874;
  assign v_3856 = ~v_3857;
  assign v_3858 = v_3859 | v_3861;
  assign v_3859 = act_3860 & 1'h1;
  assign act_3860 = v_2444 | v_2438;
  assign v_3861 = v_3862 & 1'h1;
  assign v_3862 = v_3863 & v_3864;
  assign v_3863 = ~act_3860;
  assign v_3864 = v_3865 | v_3870;
  assign v_3865 = v_3866 | v_3868;
  assign v_3866 = mux_3866(v_3867);
  assign v_3867 = v_3857 & 1'h1;
  assign v_3868 = mux_3868(v_3869);
  assign v_3869 = ~v_3867;
  assign v_3870 = ~v_3857;
  assign v_3871 = v_3872 | v_3873;
  assign v_3872 = mux_3872(v_3859);
  assign v_3873 = mux_3873(v_3861);
  assign v_3875 = v_3876 | v_3878;
  assign v_3876 = act_3877 & 1'h1;
  assign act_3877 = v_2458 | v_2452;
  assign v_3878 = v_3879 & 1'h1;
  assign v_3879 = v_3880 & v_3881;
  assign v_3880 = ~act_3877;
  assign v_3881 = v_3882 | v_3886;
  assign v_3882 = v_3883 | v_3884;
  assign v_3883 = mux_3883(v_3854);
  assign v_3884 = mux_3884(v_3885);
  assign v_3885 = ~v_3854;
  assign v_3886 = ~v_3874;
  assign v_3887 = v_3888 | v_3889;
  assign v_3888 = mux_3888(v_3876);
  assign v_3889 = mux_3889(v_3878);
  assign v_3890 = v_3891 & 1'h1;
  assign v_3891 = v_3892 & v_3893;
  assign v_3892 = ~act_3853;
  assign v_3893 = v_3894 | v_3898;
  assign v_3894 = v_3895 | v_3896;
  assign v_3895 = mux_3895(v_3794);
  assign v_3896 = mux_3896(v_3897);
  assign v_3897 = ~v_3794;
  assign v_3898 = ~v_3850;
  assign v_3899 = v_3900 | v_3901;
  assign v_3900 = mux_3900(v_3852);
  assign v_3901 = mux_3901(v_3890);
  assign v_3902 = v_3903 & 1'h1;
  assign v_3903 = v_3904 & v_3905;
  assign v_3904 = ~act_3793;
  assign v_3905 = v_3906 | v_3910;
  assign v_3906 = v_3907 | v_3908;
  assign v_3907 = mux_3907(v_3662);
  assign v_3908 = mux_3908(v_3909);
  assign v_3909 = ~v_3662;
  assign v_3910 = ~v_3790;
  assign v_3911 = v_3912 | v_3913;
  assign v_3912 = mux_3912(v_3792);
  assign v_3913 = mux_3913(v_3902);
  assign v_3914 = v_3915 & 1'h1;
  assign v_3915 = v_3916 & v_3917;
  assign v_3916 = ~act_3661;
  assign v_3917 = v_3918 | v_3922;
  assign v_3918 = v_3919 | v_3920;
  assign v_3919 = mux_3919(v_3386);
  assign v_3920 = mux_3920(v_3921);
  assign v_3921 = ~v_3386;
  assign v_3922 = ~v_3658;
  assign v_3923 = v_3924 | v_3925;
  assign v_3924 = mux_3924(v_3660);
  assign v_3925 = mux_3925(v_3914);
  assign v_3926 = v_3927 & 1'h1;
  assign v_3927 = v_3928 & v_3929;
  assign v_3928 = ~act_3385;
  assign v_3929 = v_3930 | v_3934;
  assign v_3930 = v_3931 | v_3932;
  assign v_3931 = mux_3931(v_2822);
  assign v_3932 = mux_3932(v_3933);
  assign v_3933 = ~v_2822;
  assign v_3934 = ~v_3382;
  assign v_3935 = v_3936 | v_3937;
  assign v_3936 = mux_3936(v_3384);
  assign v_3937 = mux_3937(v_3926);
  assign v_3938 = v_3939 & 1'h1;
  assign v_3939 = v_3940 & v_3941;
  assign v_3940 = ~act_2821;
  assign v_3941 = v_3942 | v_3947;
  assign v_3942 = v_3943 | v_3945;
  assign v_3943 = mux_3943(v_3944);
  assign v_3944 = v_2818 & 1'h1;
  assign v_3945 = mux_3945(v_3946);
  assign v_3946 = ~v_3944;
  assign v_3947 = ~v_2818;
  assign v_3948 = v_3949 | v_3950;
  assign v_3949 = mux_3949(v_2820);
  assign v_3950 = mux_3950(v_3938);
  assign v_3952 = v_3953 | v_5359;
  assign v_3953 = act_3954 & 1'h1;
  assign act_3954 = v_3955 | v_4508;
  assign v_3955 = v_3956 & 1'h1;
  assign v_3956 = v_3957 & v_4515;
  assign v_3957 = ~v_3958;
  assign v_3959 = v_3960 | v_4502;
  assign v_3960 = act_3961 & 1'h1;
  assign act_3961 = v_3962 | v_4227;
  assign v_3962 = v_3963 & 1'h1;
  assign v_3963 = v_3964 & v_4234;
  assign v_3964 = ~v_3965;
  assign v_3966 = v_3967 | v_4221;
  assign v_3967 = act_3968 & 1'h1;
  assign act_3968 = v_3969 | v_4090;
  assign v_3969 = v_3970 & 1'h1;
  assign v_3970 = v_3971 & v_4097;
  assign v_3971 = ~v_3972;
  assign v_3973 = v_3974 | v_4084;
  assign v_3974 = act_3975 & 1'h1;
  assign act_3975 = v_3976 | v_4025;
  assign v_3976 = v_3977 & 1'h1;
  assign v_3977 = v_3978 & v_4032;
  assign v_3978 = ~v_3979;
  assign v_3980 = v_3981 | v_4019;
  assign v_3981 = act_3982 & 1'h1;
  assign act_3982 = v_3983 | v_3996;
  assign v_3983 = v_3984 & 1'h1;
  assign v_3984 = v_3985 & v_4003;
  assign v_3985 = ~v_3986;
  assign v_3987 = v_3988 | v_3990;
  assign v_3988 = act_3989 & 1'h1;
  assign act_3989 = v_2472 | v_2466;
  assign v_3990 = v_3991 & 1'h1;
  assign v_3991 = v_3992 & v_3993;
  assign v_3992 = ~act_3989;
  assign v_3993 = v_3994 | v_3999;
  assign v_3994 = v_3995 | v_3997;
  assign v_3995 = mux_3995(v_3996);
  assign v_3996 = v_3986 & 1'h1;
  assign v_3997 = mux_3997(v_3998);
  assign v_3998 = ~v_3996;
  assign v_3999 = ~v_3986;
  assign v_4000 = v_4001 | v_4002;
  assign v_4001 = mux_4001(v_3988);
  assign v_4002 = mux_4002(v_3990);
  assign v_4004 = v_4005 | v_4007;
  assign v_4005 = act_4006 & 1'h1;
  assign act_4006 = v_2486 | v_2480;
  assign v_4007 = v_4008 & 1'h1;
  assign v_4008 = v_4009 & v_4010;
  assign v_4009 = ~act_4006;
  assign v_4010 = v_4011 | v_4015;
  assign v_4011 = v_4012 | v_4013;
  assign v_4012 = mux_4012(v_3983);
  assign v_4013 = mux_4013(v_4014);
  assign v_4014 = ~v_3983;
  assign v_4015 = ~v_4003;
  assign v_4016 = v_4017 | v_4018;
  assign v_4017 = mux_4017(v_4005);
  assign v_4018 = mux_4018(v_4007);
  assign v_4019 = v_4020 & 1'h1;
  assign v_4020 = v_4021 & v_4022;
  assign v_4021 = ~act_3982;
  assign v_4022 = v_4023 | v_4028;
  assign v_4023 = v_4024 | v_4026;
  assign v_4024 = mux_4024(v_4025);
  assign v_4025 = v_3979 & 1'h1;
  assign v_4026 = mux_4026(v_4027);
  assign v_4027 = ~v_4025;
  assign v_4028 = ~v_3979;
  assign v_4029 = v_4030 | v_4031;
  assign v_4030 = mux_4030(v_3981);
  assign v_4031 = mux_4031(v_4019);
  assign v_4033 = v_4034 | v_4072;
  assign v_4034 = act_4035 & 1'h1;
  assign act_4035 = v_4036 | v_4049;
  assign v_4036 = v_4037 & 1'h1;
  assign v_4037 = v_4038 & v_4056;
  assign v_4038 = ~v_4039;
  assign v_4040 = v_4041 | v_4043;
  assign v_4041 = act_4042 & 1'h1;
  assign act_4042 = v_2500 | v_2494;
  assign v_4043 = v_4044 & 1'h1;
  assign v_4044 = v_4045 & v_4046;
  assign v_4045 = ~act_4042;
  assign v_4046 = v_4047 | v_4052;
  assign v_4047 = v_4048 | v_4050;
  assign v_4048 = mux_4048(v_4049);
  assign v_4049 = v_4039 & 1'h1;
  assign v_4050 = mux_4050(v_4051);
  assign v_4051 = ~v_4049;
  assign v_4052 = ~v_4039;
  assign v_4053 = v_4054 | v_4055;
  assign v_4054 = mux_4054(v_4041);
  assign v_4055 = mux_4055(v_4043);
  assign v_4057 = v_4058 | v_4060;
  assign v_4058 = act_4059 & 1'h1;
  assign act_4059 = v_2514 | v_2508;
  assign v_4060 = v_4061 & 1'h1;
  assign v_4061 = v_4062 & v_4063;
  assign v_4062 = ~act_4059;
  assign v_4063 = v_4064 | v_4068;
  assign v_4064 = v_4065 | v_4066;
  assign v_4065 = mux_4065(v_4036);
  assign v_4066 = mux_4066(v_4067);
  assign v_4067 = ~v_4036;
  assign v_4068 = ~v_4056;
  assign v_4069 = v_4070 | v_4071;
  assign v_4070 = mux_4070(v_4058);
  assign v_4071 = mux_4071(v_4060);
  assign v_4072 = v_4073 & 1'h1;
  assign v_4073 = v_4074 & v_4075;
  assign v_4074 = ~act_4035;
  assign v_4075 = v_4076 | v_4080;
  assign v_4076 = v_4077 | v_4078;
  assign v_4077 = mux_4077(v_3976);
  assign v_4078 = mux_4078(v_4079);
  assign v_4079 = ~v_3976;
  assign v_4080 = ~v_4032;
  assign v_4081 = v_4082 | v_4083;
  assign v_4082 = mux_4082(v_4034);
  assign v_4083 = mux_4083(v_4072);
  assign v_4084 = v_4085 & 1'h1;
  assign v_4085 = v_4086 & v_4087;
  assign v_4086 = ~act_3975;
  assign v_4087 = v_4088 | v_4093;
  assign v_4088 = v_4089 | v_4091;
  assign v_4089 = mux_4089(v_4090);
  assign v_4090 = v_3972 & 1'h1;
  assign v_4091 = mux_4091(v_4092);
  assign v_4092 = ~v_4090;
  assign v_4093 = ~v_3972;
  assign v_4094 = v_4095 | v_4096;
  assign v_4095 = mux_4095(v_3974);
  assign v_4096 = mux_4096(v_4084);
  assign v_4098 = v_4099 | v_4209;
  assign v_4099 = act_4100 & 1'h1;
  assign act_4100 = v_4101 | v_4150;
  assign v_4101 = v_4102 & 1'h1;
  assign v_4102 = v_4103 & v_4157;
  assign v_4103 = ~v_4104;
  assign v_4105 = v_4106 | v_4144;
  assign v_4106 = act_4107 & 1'h1;
  assign act_4107 = v_4108 | v_4121;
  assign v_4108 = v_4109 & 1'h1;
  assign v_4109 = v_4110 & v_4128;
  assign v_4110 = ~v_4111;
  assign v_4112 = v_4113 | v_4115;
  assign v_4113 = act_4114 & 1'h1;
  assign act_4114 = v_2528 | v_2522;
  assign v_4115 = v_4116 & 1'h1;
  assign v_4116 = v_4117 & v_4118;
  assign v_4117 = ~act_4114;
  assign v_4118 = v_4119 | v_4124;
  assign v_4119 = v_4120 | v_4122;
  assign v_4120 = mux_4120(v_4121);
  assign v_4121 = v_4111 & 1'h1;
  assign v_4122 = mux_4122(v_4123);
  assign v_4123 = ~v_4121;
  assign v_4124 = ~v_4111;
  assign v_4125 = v_4126 | v_4127;
  assign v_4126 = mux_4126(v_4113);
  assign v_4127 = mux_4127(v_4115);
  assign v_4129 = v_4130 | v_4132;
  assign v_4130 = act_4131 & 1'h1;
  assign act_4131 = v_2542 | v_2536;
  assign v_4132 = v_4133 & 1'h1;
  assign v_4133 = v_4134 & v_4135;
  assign v_4134 = ~act_4131;
  assign v_4135 = v_4136 | v_4140;
  assign v_4136 = v_4137 | v_4138;
  assign v_4137 = mux_4137(v_4108);
  assign v_4138 = mux_4138(v_4139);
  assign v_4139 = ~v_4108;
  assign v_4140 = ~v_4128;
  assign v_4141 = v_4142 | v_4143;
  assign v_4142 = mux_4142(v_4130);
  assign v_4143 = mux_4143(v_4132);
  assign v_4144 = v_4145 & 1'h1;
  assign v_4145 = v_4146 & v_4147;
  assign v_4146 = ~act_4107;
  assign v_4147 = v_4148 | v_4153;
  assign v_4148 = v_4149 | v_4151;
  assign v_4149 = mux_4149(v_4150);
  assign v_4150 = v_4104 & 1'h1;
  assign v_4151 = mux_4151(v_4152);
  assign v_4152 = ~v_4150;
  assign v_4153 = ~v_4104;
  assign v_4154 = v_4155 | v_4156;
  assign v_4155 = mux_4155(v_4106);
  assign v_4156 = mux_4156(v_4144);
  assign v_4158 = v_4159 | v_4197;
  assign v_4159 = act_4160 & 1'h1;
  assign act_4160 = v_4161 | v_4174;
  assign v_4161 = v_4162 & 1'h1;
  assign v_4162 = v_4163 & v_4181;
  assign v_4163 = ~v_4164;
  assign v_4165 = v_4166 | v_4168;
  assign v_4166 = act_4167 & 1'h1;
  assign act_4167 = v_2556 | v_2550;
  assign v_4168 = v_4169 & 1'h1;
  assign v_4169 = v_4170 & v_4171;
  assign v_4170 = ~act_4167;
  assign v_4171 = v_4172 | v_4177;
  assign v_4172 = v_4173 | v_4175;
  assign v_4173 = mux_4173(v_4174);
  assign v_4174 = v_4164 & 1'h1;
  assign v_4175 = mux_4175(v_4176);
  assign v_4176 = ~v_4174;
  assign v_4177 = ~v_4164;
  assign v_4178 = v_4179 | v_4180;
  assign v_4179 = mux_4179(v_4166);
  assign v_4180 = mux_4180(v_4168);
  assign v_4182 = v_4183 | v_4185;
  assign v_4183 = act_4184 & 1'h1;
  assign act_4184 = v_2570 | v_2564;
  assign v_4185 = v_4186 & 1'h1;
  assign v_4186 = v_4187 & v_4188;
  assign v_4187 = ~act_4184;
  assign v_4188 = v_4189 | v_4193;
  assign v_4189 = v_4190 | v_4191;
  assign v_4190 = mux_4190(v_4161);
  assign v_4191 = mux_4191(v_4192);
  assign v_4192 = ~v_4161;
  assign v_4193 = ~v_4181;
  assign v_4194 = v_4195 | v_4196;
  assign v_4195 = mux_4195(v_4183);
  assign v_4196 = mux_4196(v_4185);
  assign v_4197 = v_4198 & 1'h1;
  assign v_4198 = v_4199 & v_4200;
  assign v_4199 = ~act_4160;
  assign v_4200 = v_4201 | v_4205;
  assign v_4201 = v_4202 | v_4203;
  assign v_4202 = mux_4202(v_4101);
  assign v_4203 = mux_4203(v_4204);
  assign v_4204 = ~v_4101;
  assign v_4205 = ~v_4157;
  assign v_4206 = v_4207 | v_4208;
  assign v_4207 = mux_4207(v_4159);
  assign v_4208 = mux_4208(v_4197);
  assign v_4209 = v_4210 & 1'h1;
  assign v_4210 = v_4211 & v_4212;
  assign v_4211 = ~act_4100;
  assign v_4212 = v_4213 | v_4217;
  assign v_4213 = v_4214 | v_4215;
  assign v_4214 = mux_4214(v_3969);
  assign v_4215 = mux_4215(v_4216);
  assign v_4216 = ~v_3969;
  assign v_4217 = ~v_4097;
  assign v_4218 = v_4219 | v_4220;
  assign v_4219 = mux_4219(v_4099);
  assign v_4220 = mux_4220(v_4209);
  assign v_4221 = v_4222 & 1'h1;
  assign v_4222 = v_4223 & v_4224;
  assign v_4223 = ~act_3968;
  assign v_4224 = v_4225 | v_4230;
  assign v_4225 = v_4226 | v_4228;
  assign v_4226 = mux_4226(v_4227);
  assign v_4227 = v_3965 & 1'h1;
  assign v_4228 = mux_4228(v_4229);
  assign v_4229 = ~v_4227;
  assign v_4230 = ~v_3965;
  assign v_4231 = v_4232 | v_4233;
  assign v_4232 = mux_4232(v_3967);
  assign v_4233 = mux_4233(v_4221);
  assign v_4235 = v_4236 | v_4490;
  assign v_4236 = act_4237 & 1'h1;
  assign act_4237 = v_4238 | v_4359;
  assign v_4238 = v_4239 & 1'h1;
  assign v_4239 = v_4240 & v_4366;
  assign v_4240 = ~v_4241;
  assign v_4242 = v_4243 | v_4353;
  assign v_4243 = act_4244 & 1'h1;
  assign act_4244 = v_4245 | v_4294;
  assign v_4245 = v_4246 & 1'h1;
  assign v_4246 = v_4247 & v_4301;
  assign v_4247 = ~v_4248;
  assign v_4249 = v_4250 | v_4288;
  assign v_4250 = act_4251 & 1'h1;
  assign act_4251 = v_4252 | v_4265;
  assign v_4252 = v_4253 & 1'h1;
  assign v_4253 = v_4254 & v_4272;
  assign v_4254 = ~v_4255;
  assign v_4256 = v_4257 | v_4259;
  assign v_4257 = act_4258 & 1'h1;
  assign act_4258 = v_2584 | v_2578;
  assign v_4259 = v_4260 & 1'h1;
  assign v_4260 = v_4261 & v_4262;
  assign v_4261 = ~act_4258;
  assign v_4262 = v_4263 | v_4268;
  assign v_4263 = v_4264 | v_4266;
  assign v_4264 = mux_4264(v_4265);
  assign v_4265 = v_4255 & 1'h1;
  assign v_4266 = mux_4266(v_4267);
  assign v_4267 = ~v_4265;
  assign v_4268 = ~v_4255;
  assign v_4269 = v_4270 | v_4271;
  assign v_4270 = mux_4270(v_4257);
  assign v_4271 = mux_4271(v_4259);
  assign v_4273 = v_4274 | v_4276;
  assign v_4274 = act_4275 & 1'h1;
  assign act_4275 = v_2598 | v_2592;
  assign v_4276 = v_4277 & 1'h1;
  assign v_4277 = v_4278 & v_4279;
  assign v_4278 = ~act_4275;
  assign v_4279 = v_4280 | v_4284;
  assign v_4280 = v_4281 | v_4282;
  assign v_4281 = mux_4281(v_4252);
  assign v_4282 = mux_4282(v_4283);
  assign v_4283 = ~v_4252;
  assign v_4284 = ~v_4272;
  assign v_4285 = v_4286 | v_4287;
  assign v_4286 = mux_4286(v_4274);
  assign v_4287 = mux_4287(v_4276);
  assign v_4288 = v_4289 & 1'h1;
  assign v_4289 = v_4290 & v_4291;
  assign v_4290 = ~act_4251;
  assign v_4291 = v_4292 | v_4297;
  assign v_4292 = v_4293 | v_4295;
  assign v_4293 = mux_4293(v_4294);
  assign v_4294 = v_4248 & 1'h1;
  assign v_4295 = mux_4295(v_4296);
  assign v_4296 = ~v_4294;
  assign v_4297 = ~v_4248;
  assign v_4298 = v_4299 | v_4300;
  assign v_4299 = mux_4299(v_4250);
  assign v_4300 = mux_4300(v_4288);
  assign v_4302 = v_4303 | v_4341;
  assign v_4303 = act_4304 & 1'h1;
  assign act_4304 = v_4305 | v_4318;
  assign v_4305 = v_4306 & 1'h1;
  assign v_4306 = v_4307 & v_4325;
  assign v_4307 = ~v_4308;
  assign v_4309 = v_4310 | v_4312;
  assign v_4310 = act_4311 & 1'h1;
  assign act_4311 = v_2612 | v_2606;
  assign v_4312 = v_4313 & 1'h1;
  assign v_4313 = v_4314 & v_4315;
  assign v_4314 = ~act_4311;
  assign v_4315 = v_4316 | v_4321;
  assign v_4316 = v_4317 | v_4319;
  assign v_4317 = mux_4317(v_4318);
  assign v_4318 = v_4308 & 1'h1;
  assign v_4319 = mux_4319(v_4320);
  assign v_4320 = ~v_4318;
  assign v_4321 = ~v_4308;
  assign v_4322 = v_4323 | v_4324;
  assign v_4323 = mux_4323(v_4310);
  assign v_4324 = mux_4324(v_4312);
  assign v_4326 = v_4327 | v_4329;
  assign v_4327 = act_4328 & 1'h1;
  assign act_4328 = v_2626 | v_2620;
  assign v_4329 = v_4330 & 1'h1;
  assign v_4330 = v_4331 & v_4332;
  assign v_4331 = ~act_4328;
  assign v_4332 = v_4333 | v_4337;
  assign v_4333 = v_4334 | v_4335;
  assign v_4334 = mux_4334(v_4305);
  assign v_4335 = mux_4335(v_4336);
  assign v_4336 = ~v_4305;
  assign v_4337 = ~v_4325;
  assign v_4338 = v_4339 | v_4340;
  assign v_4339 = mux_4339(v_4327);
  assign v_4340 = mux_4340(v_4329);
  assign v_4341 = v_4342 & 1'h1;
  assign v_4342 = v_4343 & v_4344;
  assign v_4343 = ~act_4304;
  assign v_4344 = v_4345 | v_4349;
  assign v_4345 = v_4346 | v_4347;
  assign v_4346 = mux_4346(v_4245);
  assign v_4347 = mux_4347(v_4348);
  assign v_4348 = ~v_4245;
  assign v_4349 = ~v_4301;
  assign v_4350 = v_4351 | v_4352;
  assign v_4351 = mux_4351(v_4303);
  assign v_4352 = mux_4352(v_4341);
  assign v_4353 = v_4354 & 1'h1;
  assign v_4354 = v_4355 & v_4356;
  assign v_4355 = ~act_4244;
  assign v_4356 = v_4357 | v_4362;
  assign v_4357 = v_4358 | v_4360;
  assign v_4358 = mux_4358(v_4359);
  assign v_4359 = v_4241 & 1'h1;
  assign v_4360 = mux_4360(v_4361);
  assign v_4361 = ~v_4359;
  assign v_4362 = ~v_4241;
  assign v_4363 = v_4364 | v_4365;
  assign v_4364 = mux_4364(v_4243);
  assign v_4365 = mux_4365(v_4353);
  assign v_4367 = v_4368 | v_4478;
  assign v_4368 = act_4369 & 1'h1;
  assign act_4369 = v_4370 | v_4419;
  assign v_4370 = v_4371 & 1'h1;
  assign v_4371 = v_4372 & v_4426;
  assign v_4372 = ~v_4373;
  assign v_4374 = v_4375 | v_4413;
  assign v_4375 = act_4376 & 1'h1;
  assign act_4376 = v_4377 | v_4390;
  assign v_4377 = v_4378 & 1'h1;
  assign v_4378 = v_4379 & v_4397;
  assign v_4379 = ~v_4380;
  assign v_4381 = v_4382 | v_4384;
  assign v_4382 = act_4383 & 1'h1;
  assign act_4383 = v_2640 | v_2634;
  assign v_4384 = v_4385 & 1'h1;
  assign v_4385 = v_4386 & v_4387;
  assign v_4386 = ~act_4383;
  assign v_4387 = v_4388 | v_4393;
  assign v_4388 = v_4389 | v_4391;
  assign v_4389 = mux_4389(v_4390);
  assign v_4390 = v_4380 & 1'h1;
  assign v_4391 = mux_4391(v_4392);
  assign v_4392 = ~v_4390;
  assign v_4393 = ~v_4380;
  assign v_4394 = v_4395 | v_4396;
  assign v_4395 = mux_4395(v_4382);
  assign v_4396 = mux_4396(v_4384);
  assign v_4398 = v_4399 | v_4401;
  assign v_4399 = act_4400 & 1'h1;
  assign act_4400 = v_2654 | v_2648;
  assign v_4401 = v_4402 & 1'h1;
  assign v_4402 = v_4403 & v_4404;
  assign v_4403 = ~act_4400;
  assign v_4404 = v_4405 | v_4409;
  assign v_4405 = v_4406 | v_4407;
  assign v_4406 = mux_4406(v_4377);
  assign v_4407 = mux_4407(v_4408);
  assign v_4408 = ~v_4377;
  assign v_4409 = ~v_4397;
  assign v_4410 = v_4411 | v_4412;
  assign v_4411 = mux_4411(v_4399);
  assign v_4412 = mux_4412(v_4401);
  assign v_4413 = v_4414 & 1'h1;
  assign v_4414 = v_4415 & v_4416;
  assign v_4415 = ~act_4376;
  assign v_4416 = v_4417 | v_4422;
  assign v_4417 = v_4418 | v_4420;
  assign v_4418 = mux_4418(v_4419);
  assign v_4419 = v_4373 & 1'h1;
  assign v_4420 = mux_4420(v_4421);
  assign v_4421 = ~v_4419;
  assign v_4422 = ~v_4373;
  assign v_4423 = v_4424 | v_4425;
  assign v_4424 = mux_4424(v_4375);
  assign v_4425 = mux_4425(v_4413);
  assign v_4427 = v_4428 | v_4466;
  assign v_4428 = act_4429 & 1'h1;
  assign act_4429 = v_4430 | v_4443;
  assign v_4430 = v_4431 & 1'h1;
  assign v_4431 = v_4432 & v_4450;
  assign v_4432 = ~v_4433;
  assign v_4434 = v_4435 | v_4437;
  assign v_4435 = act_4436 & 1'h1;
  assign act_4436 = v_2668 | v_2662;
  assign v_4437 = v_4438 & 1'h1;
  assign v_4438 = v_4439 & v_4440;
  assign v_4439 = ~act_4436;
  assign v_4440 = v_4441 | v_4446;
  assign v_4441 = v_4442 | v_4444;
  assign v_4442 = mux_4442(v_4443);
  assign v_4443 = v_4433 & 1'h1;
  assign v_4444 = mux_4444(v_4445);
  assign v_4445 = ~v_4443;
  assign v_4446 = ~v_4433;
  assign v_4447 = v_4448 | v_4449;
  assign v_4448 = mux_4448(v_4435);
  assign v_4449 = mux_4449(v_4437);
  assign v_4451 = v_4452 | v_4454;
  assign v_4452 = act_4453 & 1'h1;
  assign act_4453 = v_2682 | v_2676;
  assign v_4454 = v_4455 & 1'h1;
  assign v_4455 = v_4456 & v_4457;
  assign v_4456 = ~act_4453;
  assign v_4457 = v_4458 | v_4462;
  assign v_4458 = v_4459 | v_4460;
  assign v_4459 = mux_4459(v_4430);
  assign v_4460 = mux_4460(v_4461);
  assign v_4461 = ~v_4430;
  assign v_4462 = ~v_4450;
  assign v_4463 = v_4464 | v_4465;
  assign v_4464 = mux_4464(v_4452);
  assign v_4465 = mux_4465(v_4454);
  assign v_4466 = v_4467 & 1'h1;
  assign v_4467 = v_4468 & v_4469;
  assign v_4468 = ~act_4429;
  assign v_4469 = v_4470 | v_4474;
  assign v_4470 = v_4471 | v_4472;
  assign v_4471 = mux_4471(v_4370);
  assign v_4472 = mux_4472(v_4473);
  assign v_4473 = ~v_4370;
  assign v_4474 = ~v_4426;
  assign v_4475 = v_4476 | v_4477;
  assign v_4476 = mux_4476(v_4428);
  assign v_4477 = mux_4477(v_4466);
  assign v_4478 = v_4479 & 1'h1;
  assign v_4479 = v_4480 & v_4481;
  assign v_4480 = ~act_4369;
  assign v_4481 = v_4482 | v_4486;
  assign v_4482 = v_4483 | v_4484;
  assign v_4483 = mux_4483(v_4238);
  assign v_4484 = mux_4484(v_4485);
  assign v_4485 = ~v_4238;
  assign v_4486 = ~v_4366;
  assign v_4487 = v_4488 | v_4489;
  assign v_4488 = mux_4488(v_4368);
  assign v_4489 = mux_4489(v_4478);
  assign v_4490 = v_4491 & 1'h1;
  assign v_4491 = v_4492 & v_4493;
  assign v_4492 = ~act_4237;
  assign v_4493 = v_4494 | v_4498;
  assign v_4494 = v_4495 | v_4496;
  assign v_4495 = mux_4495(v_3962);
  assign v_4496 = mux_4496(v_4497);
  assign v_4497 = ~v_3962;
  assign v_4498 = ~v_4234;
  assign v_4499 = v_4500 | v_4501;
  assign v_4500 = mux_4500(v_4236);
  assign v_4501 = mux_4501(v_4490);
  assign v_4502 = v_4503 & 1'h1;
  assign v_4503 = v_4504 & v_4505;
  assign v_4504 = ~act_3961;
  assign v_4505 = v_4506 | v_4511;
  assign v_4506 = v_4507 | v_4509;
  assign v_4507 = mux_4507(v_4508);
  assign v_4508 = v_3958 & 1'h1;
  assign v_4509 = mux_4509(v_4510);
  assign v_4510 = ~v_4508;
  assign v_4511 = ~v_3958;
  assign v_4512 = v_4513 | v_4514;
  assign v_4513 = mux_4513(v_3960);
  assign v_4514 = mux_4514(v_4502);
  assign v_4516 = v_4517 | v_5347;
  assign v_4517 = act_4518 & 1'h1;
  assign act_4518 = v_4519 | v_4784;
  assign v_4519 = v_4520 & 1'h1;
  assign v_4520 = v_4521 & v_4791;
  assign v_4521 = ~v_4522;
  assign v_4523 = v_4524 | v_4778;
  assign v_4524 = act_4525 & 1'h1;
  assign act_4525 = v_4526 | v_4647;
  assign v_4526 = v_4527 & 1'h1;
  assign v_4527 = v_4528 & v_4654;
  assign v_4528 = ~v_4529;
  assign v_4530 = v_4531 | v_4641;
  assign v_4531 = act_4532 & 1'h1;
  assign act_4532 = v_4533 | v_4582;
  assign v_4533 = v_4534 & 1'h1;
  assign v_4534 = v_4535 & v_4589;
  assign v_4535 = ~v_4536;
  assign v_4537 = v_4538 | v_4576;
  assign v_4538 = act_4539 & 1'h1;
  assign act_4539 = v_4540 | v_4553;
  assign v_4540 = v_4541 & 1'h1;
  assign v_4541 = v_4542 & v_4560;
  assign v_4542 = ~v_4543;
  assign v_4544 = v_4545 | v_4547;
  assign v_4545 = act_4546 & 1'h1;
  assign act_4546 = v_2696 | v_2690;
  assign v_4547 = v_4548 & 1'h1;
  assign v_4548 = v_4549 & v_4550;
  assign v_4549 = ~act_4546;
  assign v_4550 = v_4551 | v_4556;
  assign v_4551 = v_4552 | v_4554;
  assign v_4552 = mux_4552(v_4553);
  assign v_4553 = v_4543 & 1'h1;
  assign v_4554 = mux_4554(v_4555);
  assign v_4555 = ~v_4553;
  assign v_4556 = ~v_4543;
  assign v_4557 = v_4558 | v_4559;
  assign v_4558 = mux_4558(v_4545);
  assign v_4559 = mux_4559(v_4547);
  assign v_4561 = v_4562 | v_4564;
  assign v_4562 = act_4563 & 1'h1;
  assign act_4563 = v_2710 | v_2704;
  assign v_4564 = v_4565 & 1'h1;
  assign v_4565 = v_4566 & v_4567;
  assign v_4566 = ~act_4563;
  assign v_4567 = v_4568 | v_4572;
  assign v_4568 = v_4569 | v_4570;
  assign v_4569 = mux_4569(v_4540);
  assign v_4570 = mux_4570(v_4571);
  assign v_4571 = ~v_4540;
  assign v_4572 = ~v_4560;
  assign v_4573 = v_4574 | v_4575;
  assign v_4574 = mux_4574(v_4562);
  assign v_4575 = mux_4575(v_4564);
  assign v_4576 = v_4577 & 1'h1;
  assign v_4577 = v_4578 & v_4579;
  assign v_4578 = ~act_4539;
  assign v_4579 = v_4580 | v_4585;
  assign v_4580 = v_4581 | v_4583;
  assign v_4581 = mux_4581(v_4582);
  assign v_4582 = v_4536 & 1'h1;
  assign v_4583 = mux_4583(v_4584);
  assign v_4584 = ~v_4582;
  assign v_4585 = ~v_4536;
  assign v_4586 = v_4587 | v_4588;
  assign v_4587 = mux_4587(v_4538);
  assign v_4588 = mux_4588(v_4576);
  assign v_4590 = v_4591 | v_4629;
  assign v_4591 = act_4592 & 1'h1;
  assign act_4592 = v_4593 | v_4606;
  assign v_4593 = v_4594 & 1'h1;
  assign v_4594 = v_4595 & v_4613;
  assign v_4595 = ~v_4596;
  assign v_4597 = v_4598 | v_4600;
  assign v_4598 = act_4599 & 1'h1;
  assign act_4599 = v_2724 | v_2718;
  assign v_4600 = v_4601 & 1'h1;
  assign v_4601 = v_4602 & v_4603;
  assign v_4602 = ~act_4599;
  assign v_4603 = v_4604 | v_4609;
  assign v_4604 = v_4605 | v_4607;
  assign v_4605 = mux_4605(v_4606);
  assign v_4606 = v_4596 & 1'h1;
  assign v_4607 = mux_4607(v_4608);
  assign v_4608 = ~v_4606;
  assign v_4609 = ~v_4596;
  assign v_4610 = v_4611 | v_4612;
  assign v_4611 = mux_4611(v_4598);
  assign v_4612 = mux_4612(v_4600);
  assign v_4614 = v_4615 | v_4617;
  assign v_4615 = act_4616 & 1'h1;
  assign act_4616 = v_2738 | v_2732;
  assign v_4617 = v_4618 & 1'h1;
  assign v_4618 = v_4619 & v_4620;
  assign v_4619 = ~act_4616;
  assign v_4620 = v_4621 | v_4625;
  assign v_4621 = v_4622 | v_4623;
  assign v_4622 = mux_4622(v_4593);
  assign v_4623 = mux_4623(v_4624);
  assign v_4624 = ~v_4593;
  assign v_4625 = ~v_4613;
  assign v_4626 = v_4627 | v_4628;
  assign v_4627 = mux_4627(v_4615);
  assign v_4628 = mux_4628(v_4617);
  assign v_4629 = v_4630 & 1'h1;
  assign v_4630 = v_4631 & v_4632;
  assign v_4631 = ~act_4592;
  assign v_4632 = v_4633 | v_4637;
  assign v_4633 = v_4634 | v_4635;
  assign v_4634 = mux_4634(v_4533);
  assign v_4635 = mux_4635(v_4636);
  assign v_4636 = ~v_4533;
  assign v_4637 = ~v_4589;
  assign v_4638 = v_4639 | v_4640;
  assign v_4639 = mux_4639(v_4591);
  assign v_4640 = mux_4640(v_4629);
  assign v_4641 = v_4642 & 1'h1;
  assign v_4642 = v_4643 & v_4644;
  assign v_4643 = ~act_4532;
  assign v_4644 = v_4645 | v_4650;
  assign v_4645 = v_4646 | v_4648;
  assign v_4646 = mux_4646(v_4647);
  assign v_4647 = v_4529 & 1'h1;
  assign v_4648 = mux_4648(v_4649);
  assign v_4649 = ~v_4647;
  assign v_4650 = ~v_4529;
  assign v_4651 = v_4652 | v_4653;
  assign v_4652 = mux_4652(v_4531);
  assign v_4653 = mux_4653(v_4641);
  assign v_4655 = v_4656 | v_4766;
  assign v_4656 = act_4657 & 1'h1;
  assign act_4657 = v_4658 | v_4707;
  assign v_4658 = v_4659 & 1'h1;
  assign v_4659 = v_4660 & v_4714;
  assign v_4660 = ~v_4661;
  assign v_4662 = v_4663 | v_4701;
  assign v_4663 = act_4664 & 1'h1;
  assign act_4664 = v_4665 | v_4678;
  assign v_4665 = v_4666 & 1'h1;
  assign v_4666 = v_4667 & v_4685;
  assign v_4667 = ~v_4668;
  assign v_4669 = v_4670 | v_4672;
  assign v_4670 = act_4671 & 1'h1;
  assign act_4671 = v_2752 | v_2746;
  assign v_4672 = v_4673 & 1'h1;
  assign v_4673 = v_4674 & v_4675;
  assign v_4674 = ~act_4671;
  assign v_4675 = v_4676 | v_4681;
  assign v_4676 = v_4677 | v_4679;
  assign v_4677 = mux_4677(v_4678);
  assign v_4678 = v_4668 & 1'h1;
  assign v_4679 = mux_4679(v_4680);
  assign v_4680 = ~v_4678;
  assign v_4681 = ~v_4668;
  assign v_4682 = v_4683 | v_4684;
  assign v_4683 = mux_4683(v_4670);
  assign v_4684 = mux_4684(v_4672);
  assign v_4686 = v_4687 | v_4689;
  assign v_4687 = act_4688 & 1'h1;
  assign act_4688 = v_2766 | v_2760;
  assign v_4689 = v_4690 & 1'h1;
  assign v_4690 = v_4691 & v_4692;
  assign v_4691 = ~act_4688;
  assign v_4692 = v_4693 | v_4697;
  assign v_4693 = v_4694 | v_4695;
  assign v_4694 = mux_4694(v_4665);
  assign v_4695 = mux_4695(v_4696);
  assign v_4696 = ~v_4665;
  assign v_4697 = ~v_4685;
  assign v_4698 = v_4699 | v_4700;
  assign v_4699 = mux_4699(v_4687);
  assign v_4700 = mux_4700(v_4689);
  assign v_4701 = v_4702 & 1'h1;
  assign v_4702 = v_4703 & v_4704;
  assign v_4703 = ~act_4664;
  assign v_4704 = v_4705 | v_4710;
  assign v_4705 = v_4706 | v_4708;
  assign v_4706 = mux_4706(v_4707);
  assign v_4707 = v_4661 & 1'h1;
  assign v_4708 = mux_4708(v_4709);
  assign v_4709 = ~v_4707;
  assign v_4710 = ~v_4661;
  assign v_4711 = v_4712 | v_4713;
  assign v_4712 = mux_4712(v_4663);
  assign v_4713 = mux_4713(v_4701);
  assign v_4715 = v_4716 | v_4754;
  assign v_4716 = act_4717 & 1'h1;
  assign act_4717 = v_4718 | v_4731;
  assign v_4718 = v_4719 & 1'h1;
  assign v_4719 = v_4720 & v_4738;
  assign v_4720 = ~v_4721;
  assign v_4722 = v_4723 | v_4725;
  assign v_4723 = act_4724 & 1'h1;
  assign act_4724 = v_2780 | v_2774;
  assign v_4725 = v_4726 & 1'h1;
  assign v_4726 = v_4727 & v_4728;
  assign v_4727 = ~act_4724;
  assign v_4728 = v_4729 | v_4734;
  assign v_4729 = v_4730 | v_4732;
  assign v_4730 = mux_4730(v_4731);
  assign v_4731 = v_4721 & 1'h1;
  assign v_4732 = mux_4732(v_4733);
  assign v_4733 = ~v_4731;
  assign v_4734 = ~v_4721;
  assign v_4735 = v_4736 | v_4737;
  assign v_4736 = mux_4736(v_4723);
  assign v_4737 = mux_4737(v_4725);
  assign v_4739 = v_4740 | v_4742;
  assign v_4740 = act_4741 & 1'h1;
  assign act_4741 = v_2794 | v_2788;
  assign v_4742 = v_4743 & 1'h1;
  assign v_4743 = v_4744 & v_4745;
  assign v_4744 = ~act_4741;
  assign v_4745 = v_4746 | v_4750;
  assign v_4746 = v_4747 | v_4748;
  assign v_4747 = mux_4747(v_4718);
  assign v_4748 = mux_4748(v_4749);
  assign v_4749 = ~v_4718;
  assign v_4750 = ~v_4738;
  assign v_4751 = v_4752 | v_4753;
  assign v_4752 = mux_4752(v_4740);
  assign v_4753 = mux_4753(v_4742);
  assign v_4754 = v_4755 & 1'h1;
  assign v_4755 = v_4756 & v_4757;
  assign v_4756 = ~act_4717;
  assign v_4757 = v_4758 | v_4762;
  assign v_4758 = v_4759 | v_4760;
  assign v_4759 = mux_4759(v_4658);
  assign v_4760 = mux_4760(v_4761);
  assign v_4761 = ~v_4658;
  assign v_4762 = ~v_4714;
  assign v_4763 = v_4764 | v_4765;
  assign v_4764 = mux_4764(v_4716);
  assign v_4765 = mux_4765(v_4754);
  assign v_4766 = v_4767 & 1'h1;
  assign v_4767 = v_4768 & v_4769;
  assign v_4768 = ~act_4657;
  assign v_4769 = v_4770 | v_4774;
  assign v_4770 = v_4771 | v_4772;
  assign v_4771 = mux_4771(v_4526);
  assign v_4772 = mux_4772(v_4773);
  assign v_4773 = ~v_4526;
  assign v_4774 = ~v_4654;
  assign v_4775 = v_4776 | v_4777;
  assign v_4776 = mux_4776(v_4656);
  assign v_4777 = mux_4777(v_4766);
  assign v_4778 = v_4779 & 1'h1;
  assign v_4779 = v_4780 & v_4781;
  assign v_4780 = ~act_4525;
  assign v_4781 = v_4782 | v_4787;
  assign v_4782 = v_4783 | v_4785;
  assign v_4783 = mux_4783(v_4784);
  assign v_4784 = v_4522 & 1'h1;
  assign v_4785 = mux_4785(v_4786);
  assign v_4786 = ~v_4784;
  assign v_4787 = ~v_4522;
  assign v_4788 = v_4789 | v_4790;
  assign v_4789 = mux_4789(v_4524);
  assign v_4790 = mux_4790(v_4778);
  assign v_4792 = v_4793 | v_5335;
  assign v_4793 = act_4794 & 1'h1;
  assign act_4794 = v_4795 | v_5060;
  assign v_4795 = v_4796 & 1'h1;
  assign v_4796 = v_4797 & v_5067;
  assign v_4797 = ~v_4798;
  assign v_4799 = v_4800 | v_5054;
  assign v_4800 = act_4801 & 1'h1;
  assign act_4801 = v_4802 | v_4923;
  assign v_4802 = v_4803 & 1'h1;
  assign v_4803 = v_4804 & v_4930;
  assign v_4804 = ~v_4805;
  assign v_4806 = v_4807 | v_4917;
  assign v_4807 = act_4808 & 1'h1;
  assign act_4808 = v_4809 | v_4858;
  assign v_4809 = v_4810 & 1'h1;
  assign v_4810 = v_4811 & v_4865;
  assign v_4811 = ~v_4812;
  assign v_4813 = v_4814 | v_4852;
  assign v_4814 = act_4815 & 1'h1;
  assign act_4815 = v_4816 | v_4829;
  assign v_4816 = v_4817 & 1'h1;
  assign v_4817 = v_4818 & v_4836;
  assign v_4818 = ~v_4819;
  assign v_4820 = v_4821 | v_4823;
  assign v_4821 = act_4822 & 1'h1;
  assign act_4822 = v_8 | v_2;
  assign v_4823 = v_4824 & 1'h1;
  assign v_4824 = v_4825 & v_4826;
  assign v_4825 = ~act_4822;
  assign v_4826 = v_4827 | v_4832;
  assign v_4827 = v_4828 | v_4830;
  assign v_4828 = mux_4828(v_4829);
  assign v_4829 = v_4819 & 1'h1;
  assign v_4830 = mux_4830(v_4831);
  assign v_4831 = ~v_4829;
  assign v_4832 = ~v_4819;
  assign v_4833 = v_4834 | v_4835;
  assign v_4834 = mux_4834(v_4821);
  assign v_4835 = mux_4835(v_4823);
  assign v_4837 = v_4838 | v_4840;
  assign v_4838 = act_4839 & 1'h1;
  assign act_4839 = v_22 | v_16;
  assign v_4840 = v_4841 & 1'h1;
  assign v_4841 = v_4842 & v_4843;
  assign v_4842 = ~act_4839;
  assign v_4843 = v_4844 | v_4848;
  assign v_4844 = v_4845 | v_4846;
  assign v_4845 = mux_4845(v_4816);
  assign v_4846 = mux_4846(v_4847);
  assign v_4847 = ~v_4816;
  assign v_4848 = ~v_4836;
  assign v_4849 = v_4850 | v_4851;
  assign v_4850 = mux_4850(v_4838);
  assign v_4851 = mux_4851(v_4840);
  assign v_4852 = v_4853 & 1'h1;
  assign v_4853 = v_4854 & v_4855;
  assign v_4854 = ~act_4815;
  assign v_4855 = v_4856 | v_4861;
  assign v_4856 = v_4857 | v_4859;
  assign v_4857 = mux_4857(v_4858);
  assign v_4858 = v_4812 & 1'h1;
  assign v_4859 = mux_4859(v_4860);
  assign v_4860 = ~v_4858;
  assign v_4861 = ~v_4812;
  assign v_4862 = v_4863 | v_4864;
  assign v_4863 = mux_4863(v_4814);
  assign v_4864 = mux_4864(v_4852);
  assign v_4866 = v_4867 | v_4905;
  assign v_4867 = act_4868 & 1'h1;
  assign act_4868 = v_4869 | v_4882;
  assign v_4869 = v_4870 & 1'h1;
  assign v_4870 = v_4871 & v_4889;
  assign v_4871 = ~v_4872;
  assign v_4873 = v_4874 | v_4876;
  assign v_4874 = act_4875 & 1'h1;
  assign act_4875 = v_36 | v_30;
  assign v_4876 = v_4877 & 1'h1;
  assign v_4877 = v_4878 & v_4879;
  assign v_4878 = ~act_4875;
  assign v_4879 = v_4880 | v_4885;
  assign v_4880 = v_4881 | v_4883;
  assign v_4881 = mux_4881(v_4882);
  assign v_4882 = v_4872 & 1'h1;
  assign v_4883 = mux_4883(v_4884);
  assign v_4884 = ~v_4882;
  assign v_4885 = ~v_4872;
  assign v_4886 = v_4887 | v_4888;
  assign v_4887 = mux_4887(v_4874);
  assign v_4888 = mux_4888(v_4876);
  assign v_4890 = v_4891 | v_4893;
  assign v_4891 = act_4892 & 1'h1;
  assign act_4892 = v_50 | v_44;
  assign v_4893 = v_4894 & 1'h1;
  assign v_4894 = v_4895 & v_4896;
  assign v_4895 = ~act_4892;
  assign v_4896 = v_4897 | v_4901;
  assign v_4897 = v_4898 | v_4899;
  assign v_4898 = mux_4898(v_4869);
  assign v_4899 = mux_4899(v_4900);
  assign v_4900 = ~v_4869;
  assign v_4901 = ~v_4889;
  assign v_4902 = v_4903 | v_4904;
  assign v_4903 = mux_4903(v_4891);
  assign v_4904 = mux_4904(v_4893);
  assign v_4905 = v_4906 & 1'h1;
  assign v_4906 = v_4907 & v_4908;
  assign v_4907 = ~act_4868;
  assign v_4908 = v_4909 | v_4913;
  assign v_4909 = v_4910 | v_4911;
  assign v_4910 = mux_4910(v_4809);
  assign v_4911 = mux_4911(v_4912);
  assign v_4912 = ~v_4809;
  assign v_4913 = ~v_4865;
  assign v_4914 = v_4915 | v_4916;
  assign v_4915 = mux_4915(v_4867);
  assign v_4916 = mux_4916(v_4905);
  assign v_4917 = v_4918 & 1'h1;
  assign v_4918 = v_4919 & v_4920;
  assign v_4919 = ~act_4808;
  assign v_4920 = v_4921 | v_4926;
  assign v_4921 = v_4922 | v_4924;
  assign v_4922 = mux_4922(v_4923);
  assign v_4923 = v_4805 & 1'h1;
  assign v_4924 = mux_4924(v_4925);
  assign v_4925 = ~v_4923;
  assign v_4926 = ~v_4805;
  assign v_4927 = v_4928 | v_4929;
  assign v_4928 = mux_4928(v_4807);
  assign v_4929 = mux_4929(v_4917);
  assign v_4931 = v_4932 | v_5042;
  assign v_4932 = act_4933 & 1'h1;
  assign act_4933 = v_4934 | v_4983;
  assign v_4934 = v_4935 & 1'h1;
  assign v_4935 = v_4936 & v_4990;
  assign v_4936 = ~v_4937;
  assign v_4938 = v_4939 | v_4977;
  assign v_4939 = act_4940 & 1'h1;
  assign act_4940 = v_4941 | v_4954;
  assign v_4941 = v_4942 & 1'h1;
  assign v_4942 = v_4943 & v_4961;
  assign v_4943 = ~v_4944;
  assign v_4945 = v_4946 | v_4948;
  assign v_4946 = act_4947 & 1'h1;
  assign act_4947 = v_64 | v_58;
  assign v_4948 = v_4949 & 1'h1;
  assign v_4949 = v_4950 & v_4951;
  assign v_4950 = ~act_4947;
  assign v_4951 = v_4952 | v_4957;
  assign v_4952 = v_4953 | v_4955;
  assign v_4953 = mux_4953(v_4954);
  assign v_4954 = v_4944 & 1'h1;
  assign v_4955 = mux_4955(v_4956);
  assign v_4956 = ~v_4954;
  assign v_4957 = ~v_4944;
  assign v_4958 = v_4959 | v_4960;
  assign v_4959 = mux_4959(v_4946);
  assign v_4960 = mux_4960(v_4948);
  assign v_4962 = v_4963 | v_4965;
  assign v_4963 = act_4964 & 1'h1;
  assign act_4964 = v_78 | v_72;
  assign v_4965 = v_4966 & 1'h1;
  assign v_4966 = v_4967 & v_4968;
  assign v_4967 = ~act_4964;
  assign v_4968 = v_4969 | v_4973;
  assign v_4969 = v_4970 | v_4971;
  assign v_4970 = mux_4970(v_4941);
  assign v_4971 = mux_4971(v_4972);
  assign v_4972 = ~v_4941;
  assign v_4973 = ~v_4961;
  assign v_4974 = v_4975 | v_4976;
  assign v_4975 = mux_4975(v_4963);
  assign v_4976 = mux_4976(v_4965);
  assign v_4977 = v_4978 & 1'h1;
  assign v_4978 = v_4979 & v_4980;
  assign v_4979 = ~act_4940;
  assign v_4980 = v_4981 | v_4986;
  assign v_4981 = v_4982 | v_4984;
  assign v_4982 = mux_4982(v_4983);
  assign v_4983 = v_4937 & 1'h1;
  assign v_4984 = mux_4984(v_4985);
  assign v_4985 = ~v_4983;
  assign v_4986 = ~v_4937;
  assign v_4987 = v_4988 | v_4989;
  assign v_4988 = mux_4988(v_4939);
  assign v_4989 = mux_4989(v_4977);
  assign v_4991 = v_4992 | v_5030;
  assign v_4992 = act_4993 & 1'h1;
  assign act_4993 = v_4994 | v_5007;
  assign v_4994 = v_4995 & 1'h1;
  assign v_4995 = v_4996 & v_5014;
  assign v_4996 = ~v_4997;
  assign v_4998 = v_4999 | v_5001;
  assign v_4999 = act_5000 & 1'h1;
  assign act_5000 = v_92 | v_86;
  assign v_5001 = v_5002 & 1'h1;
  assign v_5002 = v_5003 & v_5004;
  assign v_5003 = ~act_5000;
  assign v_5004 = v_5005 | v_5010;
  assign v_5005 = v_5006 | v_5008;
  assign v_5006 = mux_5006(v_5007);
  assign v_5007 = v_4997 & 1'h1;
  assign v_5008 = mux_5008(v_5009);
  assign v_5009 = ~v_5007;
  assign v_5010 = ~v_4997;
  assign v_5011 = v_5012 | v_5013;
  assign v_5012 = mux_5012(v_4999);
  assign v_5013 = mux_5013(v_5001);
  assign v_5015 = v_5016 | v_5018;
  assign v_5016 = act_5017 & 1'h1;
  assign act_5017 = v_106 | v_100;
  assign v_5018 = v_5019 & 1'h1;
  assign v_5019 = v_5020 & v_5021;
  assign v_5020 = ~act_5017;
  assign v_5021 = v_5022 | v_5026;
  assign v_5022 = v_5023 | v_5024;
  assign v_5023 = mux_5023(v_4994);
  assign v_5024 = mux_5024(v_5025);
  assign v_5025 = ~v_4994;
  assign v_5026 = ~v_5014;
  assign v_5027 = v_5028 | v_5029;
  assign v_5028 = mux_5028(v_5016);
  assign v_5029 = mux_5029(v_5018);
  assign v_5030 = v_5031 & 1'h1;
  assign v_5031 = v_5032 & v_5033;
  assign v_5032 = ~act_4993;
  assign v_5033 = v_5034 | v_5038;
  assign v_5034 = v_5035 | v_5036;
  assign v_5035 = mux_5035(v_4934);
  assign v_5036 = mux_5036(v_5037);
  assign v_5037 = ~v_4934;
  assign v_5038 = ~v_4990;
  assign v_5039 = v_5040 | v_5041;
  assign v_5040 = mux_5040(v_4992);
  assign v_5041 = mux_5041(v_5030);
  assign v_5042 = v_5043 & 1'h1;
  assign v_5043 = v_5044 & v_5045;
  assign v_5044 = ~act_4933;
  assign v_5045 = v_5046 | v_5050;
  assign v_5046 = v_5047 | v_5048;
  assign v_5047 = mux_5047(v_4802);
  assign v_5048 = mux_5048(v_5049);
  assign v_5049 = ~v_4802;
  assign v_5050 = ~v_4930;
  assign v_5051 = v_5052 | v_5053;
  assign v_5052 = mux_5052(v_4932);
  assign v_5053 = mux_5053(v_5042);
  assign v_5054 = v_5055 & 1'h1;
  assign v_5055 = v_5056 & v_5057;
  assign v_5056 = ~act_4801;
  assign v_5057 = v_5058 | v_5063;
  assign v_5058 = v_5059 | v_5061;
  assign v_5059 = mux_5059(v_5060);
  assign v_5060 = v_4798 & 1'h1;
  assign v_5061 = mux_5061(v_5062);
  assign v_5062 = ~v_5060;
  assign v_5063 = ~v_4798;
  assign v_5064 = v_5065 | v_5066;
  assign v_5065 = mux_5065(v_4800);
  assign v_5066 = mux_5066(v_5054);
  assign v_5068 = v_5069 | v_5323;
  assign v_5069 = act_5070 & 1'h1;
  assign act_5070 = v_5071 | v_5192;
  assign v_5071 = v_5072 & 1'h1;
  assign v_5072 = v_5073 & v_5199;
  assign v_5073 = ~v_5074;
  assign v_5075 = v_5076 | v_5186;
  assign v_5076 = act_5077 & 1'h1;
  assign act_5077 = v_5078 | v_5127;
  assign v_5078 = v_5079 & 1'h1;
  assign v_5079 = v_5080 & v_5134;
  assign v_5080 = ~v_5081;
  assign v_5082 = v_5083 | v_5121;
  assign v_5083 = act_5084 & 1'h1;
  assign act_5084 = v_5085 | v_5098;
  assign v_5085 = v_5086 & 1'h1;
  assign v_5086 = v_5087 & v_5105;
  assign v_5087 = ~v_5088;
  assign v_5089 = v_5090 | v_5092;
  assign v_5090 = act_5091 & 1'h1;
  assign act_5091 = v_120 | v_114;
  assign v_5092 = v_5093 & 1'h1;
  assign v_5093 = v_5094 & v_5095;
  assign v_5094 = ~act_5091;
  assign v_5095 = v_5096 | v_5101;
  assign v_5096 = v_5097 | v_5099;
  assign v_5097 = mux_5097(v_5098);
  assign v_5098 = v_5088 & 1'h1;
  assign v_5099 = mux_5099(v_5100);
  assign v_5100 = ~v_5098;
  assign v_5101 = ~v_5088;
  assign v_5102 = v_5103 | v_5104;
  assign v_5103 = mux_5103(v_5090);
  assign v_5104 = mux_5104(v_5092);
  assign v_5106 = v_5107 | v_5109;
  assign v_5107 = act_5108 & 1'h1;
  assign act_5108 = v_134 | v_128;
  assign v_5109 = v_5110 & 1'h1;
  assign v_5110 = v_5111 & v_5112;
  assign v_5111 = ~act_5108;
  assign v_5112 = v_5113 | v_5117;
  assign v_5113 = v_5114 | v_5115;
  assign v_5114 = mux_5114(v_5085);
  assign v_5115 = mux_5115(v_5116);
  assign v_5116 = ~v_5085;
  assign v_5117 = ~v_5105;
  assign v_5118 = v_5119 | v_5120;
  assign v_5119 = mux_5119(v_5107);
  assign v_5120 = mux_5120(v_5109);
  assign v_5121 = v_5122 & 1'h1;
  assign v_5122 = v_5123 & v_5124;
  assign v_5123 = ~act_5084;
  assign v_5124 = v_5125 | v_5130;
  assign v_5125 = v_5126 | v_5128;
  assign v_5126 = mux_5126(v_5127);
  assign v_5127 = v_5081 & 1'h1;
  assign v_5128 = mux_5128(v_5129);
  assign v_5129 = ~v_5127;
  assign v_5130 = ~v_5081;
  assign v_5131 = v_5132 | v_5133;
  assign v_5132 = mux_5132(v_5083);
  assign v_5133 = mux_5133(v_5121);
  assign v_5135 = v_5136 | v_5174;
  assign v_5136 = act_5137 & 1'h1;
  assign act_5137 = v_5138 | v_5151;
  assign v_5138 = v_5139 & 1'h1;
  assign v_5139 = v_5140 & v_5158;
  assign v_5140 = ~v_5141;
  assign v_5142 = v_5143 | v_5145;
  assign v_5143 = act_5144 & 1'h1;
  assign act_5144 = v_148 | v_142;
  assign v_5145 = v_5146 & 1'h1;
  assign v_5146 = v_5147 & v_5148;
  assign v_5147 = ~act_5144;
  assign v_5148 = v_5149 | v_5154;
  assign v_5149 = v_5150 | v_5152;
  assign v_5150 = mux_5150(v_5151);
  assign v_5151 = v_5141 & 1'h1;
  assign v_5152 = mux_5152(v_5153);
  assign v_5153 = ~v_5151;
  assign v_5154 = ~v_5141;
  assign v_5155 = v_5156 | v_5157;
  assign v_5156 = mux_5156(v_5143);
  assign v_5157 = mux_5157(v_5145);
  assign v_5159 = v_5160 | v_5162;
  assign v_5160 = act_5161 & 1'h1;
  assign act_5161 = v_162 | v_156;
  assign v_5162 = v_5163 & 1'h1;
  assign v_5163 = v_5164 & v_5165;
  assign v_5164 = ~act_5161;
  assign v_5165 = v_5166 | v_5170;
  assign v_5166 = v_5167 | v_5168;
  assign v_5167 = mux_5167(v_5138);
  assign v_5168 = mux_5168(v_5169);
  assign v_5169 = ~v_5138;
  assign v_5170 = ~v_5158;
  assign v_5171 = v_5172 | v_5173;
  assign v_5172 = mux_5172(v_5160);
  assign v_5173 = mux_5173(v_5162);
  assign v_5174 = v_5175 & 1'h1;
  assign v_5175 = v_5176 & v_5177;
  assign v_5176 = ~act_5137;
  assign v_5177 = v_5178 | v_5182;
  assign v_5178 = v_5179 | v_5180;
  assign v_5179 = mux_5179(v_5078);
  assign v_5180 = mux_5180(v_5181);
  assign v_5181 = ~v_5078;
  assign v_5182 = ~v_5134;
  assign v_5183 = v_5184 | v_5185;
  assign v_5184 = mux_5184(v_5136);
  assign v_5185 = mux_5185(v_5174);
  assign v_5186 = v_5187 & 1'h1;
  assign v_5187 = v_5188 & v_5189;
  assign v_5188 = ~act_5077;
  assign v_5189 = v_5190 | v_5195;
  assign v_5190 = v_5191 | v_5193;
  assign v_5191 = mux_5191(v_5192);
  assign v_5192 = v_5074 & 1'h1;
  assign v_5193 = mux_5193(v_5194);
  assign v_5194 = ~v_5192;
  assign v_5195 = ~v_5074;
  assign v_5196 = v_5197 | v_5198;
  assign v_5197 = mux_5197(v_5076);
  assign v_5198 = mux_5198(v_5186);
  assign v_5200 = v_5201 | v_5311;
  assign v_5201 = act_5202 & 1'h1;
  assign act_5202 = v_5203 | v_5252;
  assign v_5203 = v_5204 & 1'h1;
  assign v_5204 = v_5205 & v_5259;
  assign v_5205 = ~v_5206;
  assign v_5207 = v_5208 | v_5246;
  assign v_5208 = act_5209 & 1'h1;
  assign act_5209 = v_5210 | v_5223;
  assign v_5210 = v_5211 & 1'h1;
  assign v_5211 = v_5212 & v_5230;
  assign v_5212 = ~v_5213;
  assign v_5214 = v_5215 | v_5217;
  assign v_5215 = act_5216 & 1'h1;
  assign act_5216 = v_176 | v_170;
  assign v_5217 = v_5218 & 1'h1;
  assign v_5218 = v_5219 & v_5220;
  assign v_5219 = ~act_5216;
  assign v_5220 = v_5221 | v_5226;
  assign v_5221 = v_5222 | v_5224;
  assign v_5222 = mux_5222(v_5223);
  assign v_5223 = v_5213 & 1'h1;
  assign v_5224 = mux_5224(v_5225);
  assign v_5225 = ~v_5223;
  assign v_5226 = ~v_5213;
  assign v_5227 = v_5228 | v_5229;
  assign v_5228 = mux_5228(v_5215);
  assign v_5229 = mux_5229(v_5217);
  assign v_5231 = v_5232 | v_5234;
  assign v_5232 = act_5233 & 1'h1;
  assign act_5233 = v_190 | v_184;
  assign v_5234 = v_5235 & 1'h1;
  assign v_5235 = v_5236 & v_5237;
  assign v_5236 = ~act_5233;
  assign v_5237 = v_5238 | v_5242;
  assign v_5238 = v_5239 | v_5240;
  assign v_5239 = mux_5239(v_5210);
  assign v_5240 = mux_5240(v_5241);
  assign v_5241 = ~v_5210;
  assign v_5242 = ~v_5230;
  assign v_5243 = v_5244 | v_5245;
  assign v_5244 = mux_5244(v_5232);
  assign v_5245 = mux_5245(v_5234);
  assign v_5246 = v_5247 & 1'h1;
  assign v_5247 = v_5248 & v_5249;
  assign v_5248 = ~act_5209;
  assign v_5249 = v_5250 | v_5255;
  assign v_5250 = v_5251 | v_5253;
  assign v_5251 = mux_5251(v_5252);
  assign v_5252 = v_5206 & 1'h1;
  assign v_5253 = mux_5253(v_5254);
  assign v_5254 = ~v_5252;
  assign v_5255 = ~v_5206;
  assign v_5256 = v_5257 | v_5258;
  assign v_5257 = mux_5257(v_5208);
  assign v_5258 = mux_5258(v_5246);
  assign v_5260 = v_5261 | v_5299;
  assign v_5261 = act_5262 & 1'h1;
  assign act_5262 = v_5263 | v_5276;
  assign v_5263 = v_5264 & 1'h1;
  assign v_5264 = v_5265 & v_5283;
  assign v_5265 = ~v_5266;
  assign v_5267 = v_5268 | v_5270;
  assign v_5268 = act_5269 & 1'h1;
  assign act_5269 = v_204 | v_198;
  assign v_5270 = v_5271 & 1'h1;
  assign v_5271 = v_5272 & v_5273;
  assign v_5272 = ~act_5269;
  assign v_5273 = v_5274 | v_5279;
  assign v_5274 = v_5275 | v_5277;
  assign v_5275 = mux_5275(v_5276);
  assign v_5276 = v_5266 & 1'h1;
  assign v_5277 = mux_5277(v_5278);
  assign v_5278 = ~v_5276;
  assign v_5279 = ~v_5266;
  assign v_5280 = v_5281 | v_5282;
  assign v_5281 = mux_5281(v_5268);
  assign v_5282 = mux_5282(v_5270);
  assign v_5284 = v_5285 | v_5287;
  assign v_5285 = act_5286 & 1'h1;
  assign act_5286 = v_218 | v_212;
  assign v_5287 = v_5288 & 1'h1;
  assign v_5288 = v_5289 & v_5290;
  assign v_5289 = ~act_5286;
  assign v_5290 = v_5291 | v_5295;
  assign v_5291 = v_5292 | v_5293;
  assign v_5292 = mux_5292(v_5263);
  assign v_5293 = mux_5293(v_5294);
  assign v_5294 = ~v_5263;
  assign v_5295 = ~v_5283;
  assign v_5296 = v_5297 | v_5298;
  assign v_5297 = mux_5297(v_5285);
  assign v_5298 = mux_5298(v_5287);
  assign v_5299 = v_5300 & 1'h1;
  assign v_5300 = v_5301 & v_5302;
  assign v_5301 = ~act_5262;
  assign v_5302 = v_5303 | v_5307;
  assign v_5303 = v_5304 | v_5305;
  assign v_5304 = mux_5304(v_5203);
  assign v_5305 = mux_5305(v_5306);
  assign v_5306 = ~v_5203;
  assign v_5307 = ~v_5259;
  assign v_5308 = v_5309 | v_5310;
  assign v_5309 = mux_5309(v_5261);
  assign v_5310 = mux_5310(v_5299);
  assign v_5311 = v_5312 & 1'h1;
  assign v_5312 = v_5313 & v_5314;
  assign v_5313 = ~act_5202;
  assign v_5314 = v_5315 | v_5319;
  assign v_5315 = v_5316 | v_5317;
  assign v_5316 = mux_5316(v_5071);
  assign v_5317 = mux_5317(v_5318);
  assign v_5318 = ~v_5071;
  assign v_5319 = ~v_5199;
  assign v_5320 = v_5321 | v_5322;
  assign v_5321 = mux_5321(v_5201);
  assign v_5322 = mux_5322(v_5311);
  assign v_5323 = v_5324 & 1'h1;
  assign v_5324 = v_5325 & v_5326;
  assign v_5325 = ~act_5070;
  assign v_5326 = v_5327 | v_5331;
  assign v_5327 = v_5328 | v_5329;
  assign v_5328 = mux_5328(v_4795);
  assign v_5329 = mux_5329(v_5330);
  assign v_5330 = ~v_4795;
  assign v_5331 = ~v_5067;
  assign v_5332 = v_5333 | v_5334;
  assign v_5333 = mux_5333(v_5069);
  assign v_5334 = mux_5334(v_5323);
  assign v_5335 = v_5336 & 1'h1;
  assign v_5336 = v_5337 & v_5338;
  assign v_5337 = ~act_4794;
  assign v_5338 = v_5339 | v_5343;
  assign v_5339 = v_5340 | v_5341;
  assign v_5340 = mux_5340(v_4519);
  assign v_5341 = mux_5341(v_5342);
  assign v_5342 = ~v_4519;
  assign v_5343 = ~v_4791;
  assign v_5344 = v_5345 | v_5346;
  assign v_5345 = mux_5345(v_4793);
  assign v_5346 = mux_5346(v_5335);
  assign v_5347 = v_5348 & 1'h1;
  assign v_5348 = v_5349 & v_5350;
  assign v_5349 = ~act_4518;
  assign v_5350 = v_5351 | v_5355;
  assign v_5351 = v_5352 | v_5353;
  assign v_5352 = mux_5352(v_3955);
  assign v_5353 = mux_5353(v_5354);
  assign v_5354 = ~v_3955;
  assign v_5355 = ~v_4515;
  assign v_5356 = v_5357 | v_5358;
  assign v_5357 = mux_5357(v_4517);
  assign v_5358 = mux_5358(v_5347);
  assign v_5359 = v_5360 & 1'h1;
  assign v_5360 = v_5361 & v_5362;
  assign v_5361 = ~act_3954;
  assign v_5362 = v_5363 | v_5367;
  assign v_5363 = v_5364 | v_5365;
  assign v_5364 = mux_5364(v_2815);
  assign v_5365 = mux_5365(v_5366);
  assign v_5366 = ~v_2815;
  assign v_5367 = ~v_3951;
  assign v_5368 = v_5369 | v_5370;
  assign v_5369 = mux_5369(v_3953);
  assign v_5370 = mux_5370(v_5359);
  assign v_5371 = v_5372 & 1'h1;
  assign v_5372 = v_5373 & v_5374;
  assign v_5373 = ~act_2814;
  assign v_5374 = v_5375 | v_5380;
  assign v_5375 = v_5376 | v_5378;
  assign v_5376 = mux_5376(v_5377);
  assign v_5377 = v_2811 & 1'h1;
  assign v_5378 = mux_5378(v_5379);
  assign v_5379 = ~v_5377;
  assign v_5380 = ~v_2811;
  assign v_5381 = v_5382 | v_5383;
  assign v_5382 = mux_5382(v_2813);
  assign v_5383 = mux_5383(v_5371);
  assign v_5385 = v_5386 | v_9960;
  assign v_5386 = act_5387 & 1'h1;
  assign act_5387 = v_5388 | v_7669;
  assign v_5388 = v_5389 & 1'h1;
  assign v_5389 = v_5390 & v_7676;
  assign v_5390 = ~v_5391;
  assign v_5392 = v_5393 | v_7663;
  assign v_5393 = act_5394 & 1'h1;
  assign act_5394 = v_5395 | v_6524;
  assign v_5395 = v_5396 & 1'h1;
  assign v_5396 = v_5397 & v_6531;
  assign v_5397 = ~v_5398;
  assign v_5399 = v_5400 | v_6518;
  assign v_5400 = act_5401 & 1'h1;
  assign act_5401 = v_5402 | v_5955;
  assign v_5402 = v_5403 & 1'h1;
  assign v_5403 = v_5404 & v_5962;
  assign v_5404 = ~v_5405;
  assign v_5406 = v_5407 | v_5949;
  assign v_5407 = act_5408 & 1'h1;
  assign act_5408 = v_5409 | v_5674;
  assign v_5409 = v_5410 & 1'h1;
  assign v_5410 = v_5411 & v_5681;
  assign v_5411 = ~v_5412;
  assign v_5413 = v_5414 | v_5668;
  assign v_5414 = act_5415 & 1'h1;
  assign act_5415 = v_5416 | v_5537;
  assign v_5416 = v_5417 & 1'h1;
  assign v_5417 = v_5418 & v_5544;
  assign v_5418 = ~v_5419;
  assign v_5420 = v_5421 | v_5531;
  assign v_5421 = act_5422 & 1'h1;
  assign act_5422 = v_5423 | v_5472;
  assign v_5423 = v_5424 & 1'h1;
  assign v_5424 = v_5425 & v_5479;
  assign v_5425 = ~v_5426;
  assign v_5427 = v_5428 | v_5466;
  assign v_5428 = act_5429 & 1'h1;
  assign act_5429 = v_5430 | v_5443;
  assign v_5430 = v_5431 & 1'h1;
  assign v_5431 = v_5432 & v_5450;
  assign v_5432 = ~v_5433;
  assign v_5434 = v_5435 | v_5437;
  assign v_5435 = act_5436 & 1'h1;
  assign act_5436 = v_232 | v_226;
  assign v_5437 = v_5438 & 1'h1;
  assign v_5438 = v_5439 & v_5440;
  assign v_5439 = ~act_5436;
  assign v_5440 = v_5441 | v_5446;
  assign v_5441 = v_5442 | v_5444;
  assign v_5442 = mux_5442(v_5443);
  assign v_5443 = v_5433 & 1'h1;
  assign v_5444 = mux_5444(v_5445);
  assign v_5445 = ~v_5443;
  assign v_5446 = ~v_5433;
  assign v_5447 = v_5448 | v_5449;
  assign v_5448 = mux_5448(v_5435);
  assign v_5449 = mux_5449(v_5437);
  assign v_5451 = v_5452 | v_5454;
  assign v_5452 = act_5453 & 1'h1;
  assign act_5453 = v_246 | v_240;
  assign v_5454 = v_5455 & 1'h1;
  assign v_5455 = v_5456 & v_5457;
  assign v_5456 = ~act_5453;
  assign v_5457 = v_5458 | v_5462;
  assign v_5458 = v_5459 | v_5460;
  assign v_5459 = mux_5459(v_5430);
  assign v_5460 = mux_5460(v_5461);
  assign v_5461 = ~v_5430;
  assign v_5462 = ~v_5450;
  assign v_5463 = v_5464 | v_5465;
  assign v_5464 = mux_5464(v_5452);
  assign v_5465 = mux_5465(v_5454);
  assign v_5466 = v_5467 & 1'h1;
  assign v_5467 = v_5468 & v_5469;
  assign v_5468 = ~act_5429;
  assign v_5469 = v_5470 | v_5475;
  assign v_5470 = v_5471 | v_5473;
  assign v_5471 = mux_5471(v_5472);
  assign v_5472 = v_5426 & 1'h1;
  assign v_5473 = mux_5473(v_5474);
  assign v_5474 = ~v_5472;
  assign v_5475 = ~v_5426;
  assign v_5476 = v_5477 | v_5478;
  assign v_5477 = mux_5477(v_5428);
  assign v_5478 = mux_5478(v_5466);
  assign v_5480 = v_5481 | v_5519;
  assign v_5481 = act_5482 & 1'h1;
  assign act_5482 = v_5483 | v_5496;
  assign v_5483 = v_5484 & 1'h1;
  assign v_5484 = v_5485 & v_5503;
  assign v_5485 = ~v_5486;
  assign v_5487 = v_5488 | v_5490;
  assign v_5488 = act_5489 & 1'h1;
  assign act_5489 = v_260 | v_254;
  assign v_5490 = v_5491 & 1'h1;
  assign v_5491 = v_5492 & v_5493;
  assign v_5492 = ~act_5489;
  assign v_5493 = v_5494 | v_5499;
  assign v_5494 = v_5495 | v_5497;
  assign v_5495 = mux_5495(v_5496);
  assign v_5496 = v_5486 & 1'h1;
  assign v_5497 = mux_5497(v_5498);
  assign v_5498 = ~v_5496;
  assign v_5499 = ~v_5486;
  assign v_5500 = v_5501 | v_5502;
  assign v_5501 = mux_5501(v_5488);
  assign v_5502 = mux_5502(v_5490);
  assign v_5504 = v_5505 | v_5507;
  assign v_5505 = act_5506 & 1'h1;
  assign act_5506 = v_274 | v_268;
  assign v_5507 = v_5508 & 1'h1;
  assign v_5508 = v_5509 & v_5510;
  assign v_5509 = ~act_5506;
  assign v_5510 = v_5511 | v_5515;
  assign v_5511 = v_5512 | v_5513;
  assign v_5512 = mux_5512(v_5483);
  assign v_5513 = mux_5513(v_5514);
  assign v_5514 = ~v_5483;
  assign v_5515 = ~v_5503;
  assign v_5516 = v_5517 | v_5518;
  assign v_5517 = mux_5517(v_5505);
  assign v_5518 = mux_5518(v_5507);
  assign v_5519 = v_5520 & 1'h1;
  assign v_5520 = v_5521 & v_5522;
  assign v_5521 = ~act_5482;
  assign v_5522 = v_5523 | v_5527;
  assign v_5523 = v_5524 | v_5525;
  assign v_5524 = mux_5524(v_5423);
  assign v_5525 = mux_5525(v_5526);
  assign v_5526 = ~v_5423;
  assign v_5527 = ~v_5479;
  assign v_5528 = v_5529 | v_5530;
  assign v_5529 = mux_5529(v_5481);
  assign v_5530 = mux_5530(v_5519);
  assign v_5531 = v_5532 & 1'h1;
  assign v_5532 = v_5533 & v_5534;
  assign v_5533 = ~act_5422;
  assign v_5534 = v_5535 | v_5540;
  assign v_5535 = v_5536 | v_5538;
  assign v_5536 = mux_5536(v_5537);
  assign v_5537 = v_5419 & 1'h1;
  assign v_5538 = mux_5538(v_5539);
  assign v_5539 = ~v_5537;
  assign v_5540 = ~v_5419;
  assign v_5541 = v_5542 | v_5543;
  assign v_5542 = mux_5542(v_5421);
  assign v_5543 = mux_5543(v_5531);
  assign v_5545 = v_5546 | v_5656;
  assign v_5546 = act_5547 & 1'h1;
  assign act_5547 = v_5548 | v_5597;
  assign v_5548 = v_5549 & 1'h1;
  assign v_5549 = v_5550 & v_5604;
  assign v_5550 = ~v_5551;
  assign v_5552 = v_5553 | v_5591;
  assign v_5553 = act_5554 & 1'h1;
  assign act_5554 = v_5555 | v_5568;
  assign v_5555 = v_5556 & 1'h1;
  assign v_5556 = v_5557 & v_5575;
  assign v_5557 = ~v_5558;
  assign v_5559 = v_5560 | v_5562;
  assign v_5560 = act_5561 & 1'h1;
  assign act_5561 = v_288 | v_282;
  assign v_5562 = v_5563 & 1'h1;
  assign v_5563 = v_5564 & v_5565;
  assign v_5564 = ~act_5561;
  assign v_5565 = v_5566 | v_5571;
  assign v_5566 = v_5567 | v_5569;
  assign v_5567 = mux_5567(v_5568);
  assign v_5568 = v_5558 & 1'h1;
  assign v_5569 = mux_5569(v_5570);
  assign v_5570 = ~v_5568;
  assign v_5571 = ~v_5558;
  assign v_5572 = v_5573 | v_5574;
  assign v_5573 = mux_5573(v_5560);
  assign v_5574 = mux_5574(v_5562);
  assign v_5576 = v_5577 | v_5579;
  assign v_5577 = act_5578 & 1'h1;
  assign act_5578 = v_302 | v_296;
  assign v_5579 = v_5580 & 1'h1;
  assign v_5580 = v_5581 & v_5582;
  assign v_5581 = ~act_5578;
  assign v_5582 = v_5583 | v_5587;
  assign v_5583 = v_5584 | v_5585;
  assign v_5584 = mux_5584(v_5555);
  assign v_5585 = mux_5585(v_5586);
  assign v_5586 = ~v_5555;
  assign v_5587 = ~v_5575;
  assign v_5588 = v_5589 | v_5590;
  assign v_5589 = mux_5589(v_5577);
  assign v_5590 = mux_5590(v_5579);
  assign v_5591 = v_5592 & 1'h1;
  assign v_5592 = v_5593 & v_5594;
  assign v_5593 = ~act_5554;
  assign v_5594 = v_5595 | v_5600;
  assign v_5595 = v_5596 | v_5598;
  assign v_5596 = mux_5596(v_5597);
  assign v_5597 = v_5551 & 1'h1;
  assign v_5598 = mux_5598(v_5599);
  assign v_5599 = ~v_5597;
  assign v_5600 = ~v_5551;
  assign v_5601 = v_5602 | v_5603;
  assign v_5602 = mux_5602(v_5553);
  assign v_5603 = mux_5603(v_5591);
  assign v_5605 = v_5606 | v_5644;
  assign v_5606 = act_5607 & 1'h1;
  assign act_5607 = v_5608 | v_5621;
  assign v_5608 = v_5609 & 1'h1;
  assign v_5609 = v_5610 & v_5628;
  assign v_5610 = ~v_5611;
  assign v_5612 = v_5613 | v_5615;
  assign v_5613 = act_5614 & 1'h1;
  assign act_5614 = v_316 | v_310;
  assign v_5615 = v_5616 & 1'h1;
  assign v_5616 = v_5617 & v_5618;
  assign v_5617 = ~act_5614;
  assign v_5618 = v_5619 | v_5624;
  assign v_5619 = v_5620 | v_5622;
  assign v_5620 = mux_5620(v_5621);
  assign v_5621 = v_5611 & 1'h1;
  assign v_5622 = mux_5622(v_5623);
  assign v_5623 = ~v_5621;
  assign v_5624 = ~v_5611;
  assign v_5625 = v_5626 | v_5627;
  assign v_5626 = mux_5626(v_5613);
  assign v_5627 = mux_5627(v_5615);
  assign v_5629 = v_5630 | v_5632;
  assign v_5630 = act_5631 & 1'h1;
  assign act_5631 = v_330 | v_324;
  assign v_5632 = v_5633 & 1'h1;
  assign v_5633 = v_5634 & v_5635;
  assign v_5634 = ~act_5631;
  assign v_5635 = v_5636 | v_5640;
  assign v_5636 = v_5637 | v_5638;
  assign v_5637 = mux_5637(v_5608);
  assign v_5638 = mux_5638(v_5639);
  assign v_5639 = ~v_5608;
  assign v_5640 = ~v_5628;
  assign v_5641 = v_5642 | v_5643;
  assign v_5642 = mux_5642(v_5630);
  assign v_5643 = mux_5643(v_5632);
  assign v_5644 = v_5645 & 1'h1;
  assign v_5645 = v_5646 & v_5647;
  assign v_5646 = ~act_5607;
  assign v_5647 = v_5648 | v_5652;
  assign v_5648 = v_5649 | v_5650;
  assign v_5649 = mux_5649(v_5548);
  assign v_5650 = mux_5650(v_5651);
  assign v_5651 = ~v_5548;
  assign v_5652 = ~v_5604;
  assign v_5653 = v_5654 | v_5655;
  assign v_5654 = mux_5654(v_5606);
  assign v_5655 = mux_5655(v_5644);
  assign v_5656 = v_5657 & 1'h1;
  assign v_5657 = v_5658 & v_5659;
  assign v_5658 = ~act_5547;
  assign v_5659 = v_5660 | v_5664;
  assign v_5660 = v_5661 | v_5662;
  assign v_5661 = mux_5661(v_5416);
  assign v_5662 = mux_5662(v_5663);
  assign v_5663 = ~v_5416;
  assign v_5664 = ~v_5544;
  assign v_5665 = v_5666 | v_5667;
  assign v_5666 = mux_5666(v_5546);
  assign v_5667 = mux_5667(v_5656);
  assign v_5668 = v_5669 & 1'h1;
  assign v_5669 = v_5670 & v_5671;
  assign v_5670 = ~act_5415;
  assign v_5671 = v_5672 | v_5677;
  assign v_5672 = v_5673 | v_5675;
  assign v_5673 = mux_5673(v_5674);
  assign v_5674 = v_5412 & 1'h1;
  assign v_5675 = mux_5675(v_5676);
  assign v_5676 = ~v_5674;
  assign v_5677 = ~v_5412;
  assign v_5678 = v_5679 | v_5680;
  assign v_5679 = mux_5679(v_5414);
  assign v_5680 = mux_5680(v_5668);
  assign v_5682 = v_5683 | v_5937;
  assign v_5683 = act_5684 & 1'h1;
  assign act_5684 = v_5685 | v_5806;
  assign v_5685 = v_5686 & 1'h1;
  assign v_5686 = v_5687 & v_5813;
  assign v_5687 = ~v_5688;
  assign v_5689 = v_5690 | v_5800;
  assign v_5690 = act_5691 & 1'h1;
  assign act_5691 = v_5692 | v_5741;
  assign v_5692 = v_5693 & 1'h1;
  assign v_5693 = v_5694 & v_5748;
  assign v_5694 = ~v_5695;
  assign v_5696 = v_5697 | v_5735;
  assign v_5697 = act_5698 & 1'h1;
  assign act_5698 = v_5699 | v_5712;
  assign v_5699 = v_5700 & 1'h1;
  assign v_5700 = v_5701 & v_5719;
  assign v_5701 = ~v_5702;
  assign v_5703 = v_5704 | v_5706;
  assign v_5704 = act_5705 & 1'h1;
  assign act_5705 = v_344 | v_338;
  assign v_5706 = v_5707 & 1'h1;
  assign v_5707 = v_5708 & v_5709;
  assign v_5708 = ~act_5705;
  assign v_5709 = v_5710 | v_5715;
  assign v_5710 = v_5711 | v_5713;
  assign v_5711 = mux_5711(v_5712);
  assign v_5712 = v_5702 & 1'h1;
  assign v_5713 = mux_5713(v_5714);
  assign v_5714 = ~v_5712;
  assign v_5715 = ~v_5702;
  assign v_5716 = v_5717 | v_5718;
  assign v_5717 = mux_5717(v_5704);
  assign v_5718 = mux_5718(v_5706);
  assign v_5720 = v_5721 | v_5723;
  assign v_5721 = act_5722 & 1'h1;
  assign act_5722 = v_358 | v_352;
  assign v_5723 = v_5724 & 1'h1;
  assign v_5724 = v_5725 & v_5726;
  assign v_5725 = ~act_5722;
  assign v_5726 = v_5727 | v_5731;
  assign v_5727 = v_5728 | v_5729;
  assign v_5728 = mux_5728(v_5699);
  assign v_5729 = mux_5729(v_5730);
  assign v_5730 = ~v_5699;
  assign v_5731 = ~v_5719;
  assign v_5732 = v_5733 | v_5734;
  assign v_5733 = mux_5733(v_5721);
  assign v_5734 = mux_5734(v_5723);
  assign v_5735 = v_5736 & 1'h1;
  assign v_5736 = v_5737 & v_5738;
  assign v_5737 = ~act_5698;
  assign v_5738 = v_5739 | v_5744;
  assign v_5739 = v_5740 | v_5742;
  assign v_5740 = mux_5740(v_5741);
  assign v_5741 = v_5695 & 1'h1;
  assign v_5742 = mux_5742(v_5743);
  assign v_5743 = ~v_5741;
  assign v_5744 = ~v_5695;
  assign v_5745 = v_5746 | v_5747;
  assign v_5746 = mux_5746(v_5697);
  assign v_5747 = mux_5747(v_5735);
  assign v_5749 = v_5750 | v_5788;
  assign v_5750 = act_5751 & 1'h1;
  assign act_5751 = v_5752 | v_5765;
  assign v_5752 = v_5753 & 1'h1;
  assign v_5753 = v_5754 & v_5772;
  assign v_5754 = ~v_5755;
  assign v_5756 = v_5757 | v_5759;
  assign v_5757 = act_5758 & 1'h1;
  assign act_5758 = v_372 | v_366;
  assign v_5759 = v_5760 & 1'h1;
  assign v_5760 = v_5761 & v_5762;
  assign v_5761 = ~act_5758;
  assign v_5762 = v_5763 | v_5768;
  assign v_5763 = v_5764 | v_5766;
  assign v_5764 = mux_5764(v_5765);
  assign v_5765 = v_5755 & 1'h1;
  assign v_5766 = mux_5766(v_5767);
  assign v_5767 = ~v_5765;
  assign v_5768 = ~v_5755;
  assign v_5769 = v_5770 | v_5771;
  assign v_5770 = mux_5770(v_5757);
  assign v_5771 = mux_5771(v_5759);
  assign v_5773 = v_5774 | v_5776;
  assign v_5774 = act_5775 & 1'h1;
  assign act_5775 = v_386 | v_380;
  assign v_5776 = v_5777 & 1'h1;
  assign v_5777 = v_5778 & v_5779;
  assign v_5778 = ~act_5775;
  assign v_5779 = v_5780 | v_5784;
  assign v_5780 = v_5781 | v_5782;
  assign v_5781 = mux_5781(v_5752);
  assign v_5782 = mux_5782(v_5783);
  assign v_5783 = ~v_5752;
  assign v_5784 = ~v_5772;
  assign v_5785 = v_5786 | v_5787;
  assign v_5786 = mux_5786(v_5774);
  assign v_5787 = mux_5787(v_5776);
  assign v_5788 = v_5789 & 1'h1;
  assign v_5789 = v_5790 & v_5791;
  assign v_5790 = ~act_5751;
  assign v_5791 = v_5792 | v_5796;
  assign v_5792 = v_5793 | v_5794;
  assign v_5793 = mux_5793(v_5692);
  assign v_5794 = mux_5794(v_5795);
  assign v_5795 = ~v_5692;
  assign v_5796 = ~v_5748;
  assign v_5797 = v_5798 | v_5799;
  assign v_5798 = mux_5798(v_5750);
  assign v_5799 = mux_5799(v_5788);
  assign v_5800 = v_5801 & 1'h1;
  assign v_5801 = v_5802 & v_5803;
  assign v_5802 = ~act_5691;
  assign v_5803 = v_5804 | v_5809;
  assign v_5804 = v_5805 | v_5807;
  assign v_5805 = mux_5805(v_5806);
  assign v_5806 = v_5688 & 1'h1;
  assign v_5807 = mux_5807(v_5808);
  assign v_5808 = ~v_5806;
  assign v_5809 = ~v_5688;
  assign v_5810 = v_5811 | v_5812;
  assign v_5811 = mux_5811(v_5690);
  assign v_5812 = mux_5812(v_5800);
  assign v_5814 = v_5815 | v_5925;
  assign v_5815 = act_5816 & 1'h1;
  assign act_5816 = v_5817 | v_5866;
  assign v_5817 = v_5818 & 1'h1;
  assign v_5818 = v_5819 & v_5873;
  assign v_5819 = ~v_5820;
  assign v_5821 = v_5822 | v_5860;
  assign v_5822 = act_5823 & 1'h1;
  assign act_5823 = v_5824 | v_5837;
  assign v_5824 = v_5825 & 1'h1;
  assign v_5825 = v_5826 & v_5844;
  assign v_5826 = ~v_5827;
  assign v_5828 = v_5829 | v_5831;
  assign v_5829 = act_5830 & 1'h1;
  assign act_5830 = v_400 | v_394;
  assign v_5831 = v_5832 & 1'h1;
  assign v_5832 = v_5833 & v_5834;
  assign v_5833 = ~act_5830;
  assign v_5834 = v_5835 | v_5840;
  assign v_5835 = v_5836 | v_5838;
  assign v_5836 = mux_5836(v_5837);
  assign v_5837 = v_5827 & 1'h1;
  assign v_5838 = mux_5838(v_5839);
  assign v_5839 = ~v_5837;
  assign v_5840 = ~v_5827;
  assign v_5841 = v_5842 | v_5843;
  assign v_5842 = mux_5842(v_5829);
  assign v_5843 = mux_5843(v_5831);
  assign v_5845 = v_5846 | v_5848;
  assign v_5846 = act_5847 & 1'h1;
  assign act_5847 = v_414 | v_408;
  assign v_5848 = v_5849 & 1'h1;
  assign v_5849 = v_5850 & v_5851;
  assign v_5850 = ~act_5847;
  assign v_5851 = v_5852 | v_5856;
  assign v_5852 = v_5853 | v_5854;
  assign v_5853 = mux_5853(v_5824);
  assign v_5854 = mux_5854(v_5855);
  assign v_5855 = ~v_5824;
  assign v_5856 = ~v_5844;
  assign v_5857 = v_5858 | v_5859;
  assign v_5858 = mux_5858(v_5846);
  assign v_5859 = mux_5859(v_5848);
  assign v_5860 = v_5861 & 1'h1;
  assign v_5861 = v_5862 & v_5863;
  assign v_5862 = ~act_5823;
  assign v_5863 = v_5864 | v_5869;
  assign v_5864 = v_5865 | v_5867;
  assign v_5865 = mux_5865(v_5866);
  assign v_5866 = v_5820 & 1'h1;
  assign v_5867 = mux_5867(v_5868);
  assign v_5868 = ~v_5866;
  assign v_5869 = ~v_5820;
  assign v_5870 = v_5871 | v_5872;
  assign v_5871 = mux_5871(v_5822);
  assign v_5872 = mux_5872(v_5860);
  assign v_5874 = v_5875 | v_5913;
  assign v_5875 = act_5876 & 1'h1;
  assign act_5876 = v_5877 | v_5890;
  assign v_5877 = v_5878 & 1'h1;
  assign v_5878 = v_5879 & v_5897;
  assign v_5879 = ~v_5880;
  assign v_5881 = v_5882 | v_5884;
  assign v_5882 = act_5883 & 1'h1;
  assign act_5883 = v_428 | v_422;
  assign v_5884 = v_5885 & 1'h1;
  assign v_5885 = v_5886 & v_5887;
  assign v_5886 = ~act_5883;
  assign v_5887 = v_5888 | v_5893;
  assign v_5888 = v_5889 | v_5891;
  assign v_5889 = mux_5889(v_5890);
  assign v_5890 = v_5880 & 1'h1;
  assign v_5891 = mux_5891(v_5892);
  assign v_5892 = ~v_5890;
  assign v_5893 = ~v_5880;
  assign v_5894 = v_5895 | v_5896;
  assign v_5895 = mux_5895(v_5882);
  assign v_5896 = mux_5896(v_5884);
  assign v_5898 = v_5899 | v_5901;
  assign v_5899 = act_5900 & 1'h1;
  assign act_5900 = v_442 | v_436;
  assign v_5901 = v_5902 & 1'h1;
  assign v_5902 = v_5903 & v_5904;
  assign v_5903 = ~act_5900;
  assign v_5904 = v_5905 | v_5909;
  assign v_5905 = v_5906 | v_5907;
  assign v_5906 = mux_5906(v_5877);
  assign v_5907 = mux_5907(v_5908);
  assign v_5908 = ~v_5877;
  assign v_5909 = ~v_5897;
  assign v_5910 = v_5911 | v_5912;
  assign v_5911 = mux_5911(v_5899);
  assign v_5912 = mux_5912(v_5901);
  assign v_5913 = v_5914 & 1'h1;
  assign v_5914 = v_5915 & v_5916;
  assign v_5915 = ~act_5876;
  assign v_5916 = v_5917 | v_5921;
  assign v_5917 = v_5918 | v_5919;
  assign v_5918 = mux_5918(v_5817);
  assign v_5919 = mux_5919(v_5920);
  assign v_5920 = ~v_5817;
  assign v_5921 = ~v_5873;
  assign v_5922 = v_5923 | v_5924;
  assign v_5923 = mux_5923(v_5875);
  assign v_5924 = mux_5924(v_5913);
  assign v_5925 = v_5926 & 1'h1;
  assign v_5926 = v_5927 & v_5928;
  assign v_5927 = ~act_5816;
  assign v_5928 = v_5929 | v_5933;
  assign v_5929 = v_5930 | v_5931;
  assign v_5930 = mux_5930(v_5685);
  assign v_5931 = mux_5931(v_5932);
  assign v_5932 = ~v_5685;
  assign v_5933 = ~v_5813;
  assign v_5934 = v_5935 | v_5936;
  assign v_5935 = mux_5935(v_5815);
  assign v_5936 = mux_5936(v_5925);
  assign v_5937 = v_5938 & 1'h1;
  assign v_5938 = v_5939 & v_5940;
  assign v_5939 = ~act_5684;
  assign v_5940 = v_5941 | v_5945;
  assign v_5941 = v_5942 | v_5943;
  assign v_5942 = mux_5942(v_5409);
  assign v_5943 = mux_5943(v_5944);
  assign v_5944 = ~v_5409;
  assign v_5945 = ~v_5681;
  assign v_5946 = v_5947 | v_5948;
  assign v_5947 = mux_5947(v_5683);
  assign v_5948 = mux_5948(v_5937);
  assign v_5949 = v_5950 & 1'h1;
  assign v_5950 = v_5951 & v_5952;
  assign v_5951 = ~act_5408;
  assign v_5952 = v_5953 | v_5958;
  assign v_5953 = v_5954 | v_5956;
  assign v_5954 = mux_5954(v_5955);
  assign v_5955 = v_5405 & 1'h1;
  assign v_5956 = mux_5956(v_5957);
  assign v_5957 = ~v_5955;
  assign v_5958 = ~v_5405;
  assign v_5959 = v_5960 | v_5961;
  assign v_5960 = mux_5960(v_5407);
  assign v_5961 = mux_5961(v_5949);
  assign v_5963 = v_5964 | v_6506;
  assign v_5964 = act_5965 & 1'h1;
  assign act_5965 = v_5966 | v_6231;
  assign v_5966 = v_5967 & 1'h1;
  assign v_5967 = v_5968 & v_6238;
  assign v_5968 = ~v_5969;
  assign v_5970 = v_5971 | v_6225;
  assign v_5971 = act_5972 & 1'h1;
  assign act_5972 = v_5973 | v_6094;
  assign v_5973 = v_5974 & 1'h1;
  assign v_5974 = v_5975 & v_6101;
  assign v_5975 = ~v_5976;
  assign v_5977 = v_5978 | v_6088;
  assign v_5978 = act_5979 & 1'h1;
  assign act_5979 = v_5980 | v_6029;
  assign v_5980 = v_5981 & 1'h1;
  assign v_5981 = v_5982 & v_6036;
  assign v_5982 = ~v_5983;
  assign v_5984 = v_5985 | v_6023;
  assign v_5985 = act_5986 & 1'h1;
  assign act_5986 = v_5987 | v_6000;
  assign v_5987 = v_5988 & 1'h1;
  assign v_5988 = v_5989 & v_6007;
  assign v_5989 = ~v_5990;
  assign v_5991 = v_5992 | v_5994;
  assign v_5992 = act_5993 & 1'h1;
  assign act_5993 = v_456 | v_450;
  assign v_5994 = v_5995 & 1'h1;
  assign v_5995 = v_5996 & v_5997;
  assign v_5996 = ~act_5993;
  assign v_5997 = v_5998 | v_6003;
  assign v_5998 = v_5999 | v_6001;
  assign v_5999 = mux_5999(v_6000);
  assign v_6000 = v_5990 & 1'h1;
  assign v_6001 = mux_6001(v_6002);
  assign v_6002 = ~v_6000;
  assign v_6003 = ~v_5990;
  assign v_6004 = v_6005 | v_6006;
  assign v_6005 = mux_6005(v_5992);
  assign v_6006 = mux_6006(v_5994);
  assign v_6008 = v_6009 | v_6011;
  assign v_6009 = act_6010 & 1'h1;
  assign act_6010 = v_470 | v_464;
  assign v_6011 = v_6012 & 1'h1;
  assign v_6012 = v_6013 & v_6014;
  assign v_6013 = ~act_6010;
  assign v_6014 = v_6015 | v_6019;
  assign v_6015 = v_6016 | v_6017;
  assign v_6016 = mux_6016(v_5987);
  assign v_6017 = mux_6017(v_6018);
  assign v_6018 = ~v_5987;
  assign v_6019 = ~v_6007;
  assign v_6020 = v_6021 | v_6022;
  assign v_6021 = mux_6021(v_6009);
  assign v_6022 = mux_6022(v_6011);
  assign v_6023 = v_6024 & 1'h1;
  assign v_6024 = v_6025 & v_6026;
  assign v_6025 = ~act_5986;
  assign v_6026 = v_6027 | v_6032;
  assign v_6027 = v_6028 | v_6030;
  assign v_6028 = mux_6028(v_6029);
  assign v_6029 = v_5983 & 1'h1;
  assign v_6030 = mux_6030(v_6031);
  assign v_6031 = ~v_6029;
  assign v_6032 = ~v_5983;
  assign v_6033 = v_6034 | v_6035;
  assign v_6034 = mux_6034(v_5985);
  assign v_6035 = mux_6035(v_6023);
  assign v_6037 = v_6038 | v_6076;
  assign v_6038 = act_6039 & 1'h1;
  assign act_6039 = v_6040 | v_6053;
  assign v_6040 = v_6041 & 1'h1;
  assign v_6041 = v_6042 & v_6060;
  assign v_6042 = ~v_6043;
  assign v_6044 = v_6045 | v_6047;
  assign v_6045 = act_6046 & 1'h1;
  assign act_6046 = v_484 | v_478;
  assign v_6047 = v_6048 & 1'h1;
  assign v_6048 = v_6049 & v_6050;
  assign v_6049 = ~act_6046;
  assign v_6050 = v_6051 | v_6056;
  assign v_6051 = v_6052 | v_6054;
  assign v_6052 = mux_6052(v_6053);
  assign v_6053 = v_6043 & 1'h1;
  assign v_6054 = mux_6054(v_6055);
  assign v_6055 = ~v_6053;
  assign v_6056 = ~v_6043;
  assign v_6057 = v_6058 | v_6059;
  assign v_6058 = mux_6058(v_6045);
  assign v_6059 = mux_6059(v_6047);
  assign v_6061 = v_6062 | v_6064;
  assign v_6062 = act_6063 & 1'h1;
  assign act_6063 = v_498 | v_492;
  assign v_6064 = v_6065 & 1'h1;
  assign v_6065 = v_6066 & v_6067;
  assign v_6066 = ~act_6063;
  assign v_6067 = v_6068 | v_6072;
  assign v_6068 = v_6069 | v_6070;
  assign v_6069 = mux_6069(v_6040);
  assign v_6070 = mux_6070(v_6071);
  assign v_6071 = ~v_6040;
  assign v_6072 = ~v_6060;
  assign v_6073 = v_6074 | v_6075;
  assign v_6074 = mux_6074(v_6062);
  assign v_6075 = mux_6075(v_6064);
  assign v_6076 = v_6077 & 1'h1;
  assign v_6077 = v_6078 & v_6079;
  assign v_6078 = ~act_6039;
  assign v_6079 = v_6080 | v_6084;
  assign v_6080 = v_6081 | v_6082;
  assign v_6081 = mux_6081(v_5980);
  assign v_6082 = mux_6082(v_6083);
  assign v_6083 = ~v_5980;
  assign v_6084 = ~v_6036;
  assign v_6085 = v_6086 | v_6087;
  assign v_6086 = mux_6086(v_6038);
  assign v_6087 = mux_6087(v_6076);
  assign v_6088 = v_6089 & 1'h1;
  assign v_6089 = v_6090 & v_6091;
  assign v_6090 = ~act_5979;
  assign v_6091 = v_6092 | v_6097;
  assign v_6092 = v_6093 | v_6095;
  assign v_6093 = mux_6093(v_6094);
  assign v_6094 = v_5976 & 1'h1;
  assign v_6095 = mux_6095(v_6096);
  assign v_6096 = ~v_6094;
  assign v_6097 = ~v_5976;
  assign v_6098 = v_6099 | v_6100;
  assign v_6099 = mux_6099(v_5978);
  assign v_6100 = mux_6100(v_6088);
  assign v_6102 = v_6103 | v_6213;
  assign v_6103 = act_6104 & 1'h1;
  assign act_6104 = v_6105 | v_6154;
  assign v_6105 = v_6106 & 1'h1;
  assign v_6106 = v_6107 & v_6161;
  assign v_6107 = ~v_6108;
  assign v_6109 = v_6110 | v_6148;
  assign v_6110 = act_6111 & 1'h1;
  assign act_6111 = v_6112 | v_6125;
  assign v_6112 = v_6113 & 1'h1;
  assign v_6113 = v_6114 & v_6132;
  assign v_6114 = ~v_6115;
  assign v_6116 = v_6117 | v_6119;
  assign v_6117 = act_6118 & 1'h1;
  assign act_6118 = v_512 | v_506;
  assign v_6119 = v_6120 & 1'h1;
  assign v_6120 = v_6121 & v_6122;
  assign v_6121 = ~act_6118;
  assign v_6122 = v_6123 | v_6128;
  assign v_6123 = v_6124 | v_6126;
  assign v_6124 = mux_6124(v_6125);
  assign v_6125 = v_6115 & 1'h1;
  assign v_6126 = mux_6126(v_6127);
  assign v_6127 = ~v_6125;
  assign v_6128 = ~v_6115;
  assign v_6129 = v_6130 | v_6131;
  assign v_6130 = mux_6130(v_6117);
  assign v_6131 = mux_6131(v_6119);
  assign v_6133 = v_6134 | v_6136;
  assign v_6134 = act_6135 & 1'h1;
  assign act_6135 = v_526 | v_520;
  assign v_6136 = v_6137 & 1'h1;
  assign v_6137 = v_6138 & v_6139;
  assign v_6138 = ~act_6135;
  assign v_6139 = v_6140 | v_6144;
  assign v_6140 = v_6141 | v_6142;
  assign v_6141 = mux_6141(v_6112);
  assign v_6142 = mux_6142(v_6143);
  assign v_6143 = ~v_6112;
  assign v_6144 = ~v_6132;
  assign v_6145 = v_6146 | v_6147;
  assign v_6146 = mux_6146(v_6134);
  assign v_6147 = mux_6147(v_6136);
  assign v_6148 = v_6149 & 1'h1;
  assign v_6149 = v_6150 & v_6151;
  assign v_6150 = ~act_6111;
  assign v_6151 = v_6152 | v_6157;
  assign v_6152 = v_6153 | v_6155;
  assign v_6153 = mux_6153(v_6154);
  assign v_6154 = v_6108 & 1'h1;
  assign v_6155 = mux_6155(v_6156);
  assign v_6156 = ~v_6154;
  assign v_6157 = ~v_6108;
  assign v_6158 = v_6159 | v_6160;
  assign v_6159 = mux_6159(v_6110);
  assign v_6160 = mux_6160(v_6148);
  assign v_6162 = v_6163 | v_6201;
  assign v_6163 = act_6164 & 1'h1;
  assign act_6164 = v_6165 | v_6178;
  assign v_6165 = v_6166 & 1'h1;
  assign v_6166 = v_6167 & v_6185;
  assign v_6167 = ~v_6168;
  assign v_6169 = v_6170 | v_6172;
  assign v_6170 = act_6171 & 1'h1;
  assign act_6171 = v_540 | v_534;
  assign v_6172 = v_6173 & 1'h1;
  assign v_6173 = v_6174 & v_6175;
  assign v_6174 = ~act_6171;
  assign v_6175 = v_6176 | v_6181;
  assign v_6176 = v_6177 | v_6179;
  assign v_6177 = mux_6177(v_6178);
  assign v_6178 = v_6168 & 1'h1;
  assign v_6179 = mux_6179(v_6180);
  assign v_6180 = ~v_6178;
  assign v_6181 = ~v_6168;
  assign v_6182 = v_6183 | v_6184;
  assign v_6183 = mux_6183(v_6170);
  assign v_6184 = mux_6184(v_6172);
  assign v_6186 = v_6187 | v_6189;
  assign v_6187 = act_6188 & 1'h1;
  assign act_6188 = v_554 | v_548;
  assign v_6189 = v_6190 & 1'h1;
  assign v_6190 = v_6191 & v_6192;
  assign v_6191 = ~act_6188;
  assign v_6192 = v_6193 | v_6197;
  assign v_6193 = v_6194 | v_6195;
  assign v_6194 = mux_6194(v_6165);
  assign v_6195 = mux_6195(v_6196);
  assign v_6196 = ~v_6165;
  assign v_6197 = ~v_6185;
  assign v_6198 = v_6199 | v_6200;
  assign v_6199 = mux_6199(v_6187);
  assign v_6200 = mux_6200(v_6189);
  assign v_6201 = v_6202 & 1'h1;
  assign v_6202 = v_6203 & v_6204;
  assign v_6203 = ~act_6164;
  assign v_6204 = v_6205 | v_6209;
  assign v_6205 = v_6206 | v_6207;
  assign v_6206 = mux_6206(v_6105);
  assign v_6207 = mux_6207(v_6208);
  assign v_6208 = ~v_6105;
  assign v_6209 = ~v_6161;
  assign v_6210 = v_6211 | v_6212;
  assign v_6211 = mux_6211(v_6163);
  assign v_6212 = mux_6212(v_6201);
  assign v_6213 = v_6214 & 1'h1;
  assign v_6214 = v_6215 & v_6216;
  assign v_6215 = ~act_6104;
  assign v_6216 = v_6217 | v_6221;
  assign v_6217 = v_6218 | v_6219;
  assign v_6218 = mux_6218(v_5973);
  assign v_6219 = mux_6219(v_6220);
  assign v_6220 = ~v_5973;
  assign v_6221 = ~v_6101;
  assign v_6222 = v_6223 | v_6224;
  assign v_6223 = mux_6223(v_6103);
  assign v_6224 = mux_6224(v_6213);
  assign v_6225 = v_6226 & 1'h1;
  assign v_6226 = v_6227 & v_6228;
  assign v_6227 = ~act_5972;
  assign v_6228 = v_6229 | v_6234;
  assign v_6229 = v_6230 | v_6232;
  assign v_6230 = mux_6230(v_6231);
  assign v_6231 = v_5969 & 1'h1;
  assign v_6232 = mux_6232(v_6233);
  assign v_6233 = ~v_6231;
  assign v_6234 = ~v_5969;
  assign v_6235 = v_6236 | v_6237;
  assign v_6236 = mux_6236(v_5971);
  assign v_6237 = mux_6237(v_6225);
  assign v_6239 = v_6240 | v_6494;
  assign v_6240 = act_6241 & 1'h1;
  assign act_6241 = v_6242 | v_6363;
  assign v_6242 = v_6243 & 1'h1;
  assign v_6243 = v_6244 & v_6370;
  assign v_6244 = ~v_6245;
  assign v_6246 = v_6247 | v_6357;
  assign v_6247 = act_6248 & 1'h1;
  assign act_6248 = v_6249 | v_6298;
  assign v_6249 = v_6250 & 1'h1;
  assign v_6250 = v_6251 & v_6305;
  assign v_6251 = ~v_6252;
  assign v_6253 = v_6254 | v_6292;
  assign v_6254 = act_6255 & 1'h1;
  assign act_6255 = v_6256 | v_6269;
  assign v_6256 = v_6257 & 1'h1;
  assign v_6257 = v_6258 & v_6276;
  assign v_6258 = ~v_6259;
  assign v_6260 = v_6261 | v_6263;
  assign v_6261 = act_6262 & 1'h1;
  assign act_6262 = v_568 | v_562;
  assign v_6263 = v_6264 & 1'h1;
  assign v_6264 = v_6265 & v_6266;
  assign v_6265 = ~act_6262;
  assign v_6266 = v_6267 | v_6272;
  assign v_6267 = v_6268 | v_6270;
  assign v_6268 = mux_6268(v_6269);
  assign v_6269 = v_6259 & 1'h1;
  assign v_6270 = mux_6270(v_6271);
  assign v_6271 = ~v_6269;
  assign v_6272 = ~v_6259;
  assign v_6273 = v_6274 | v_6275;
  assign v_6274 = mux_6274(v_6261);
  assign v_6275 = mux_6275(v_6263);
  assign v_6277 = v_6278 | v_6280;
  assign v_6278 = act_6279 & 1'h1;
  assign act_6279 = v_582 | v_576;
  assign v_6280 = v_6281 & 1'h1;
  assign v_6281 = v_6282 & v_6283;
  assign v_6282 = ~act_6279;
  assign v_6283 = v_6284 | v_6288;
  assign v_6284 = v_6285 | v_6286;
  assign v_6285 = mux_6285(v_6256);
  assign v_6286 = mux_6286(v_6287);
  assign v_6287 = ~v_6256;
  assign v_6288 = ~v_6276;
  assign v_6289 = v_6290 | v_6291;
  assign v_6290 = mux_6290(v_6278);
  assign v_6291 = mux_6291(v_6280);
  assign v_6292 = v_6293 & 1'h1;
  assign v_6293 = v_6294 & v_6295;
  assign v_6294 = ~act_6255;
  assign v_6295 = v_6296 | v_6301;
  assign v_6296 = v_6297 | v_6299;
  assign v_6297 = mux_6297(v_6298);
  assign v_6298 = v_6252 & 1'h1;
  assign v_6299 = mux_6299(v_6300);
  assign v_6300 = ~v_6298;
  assign v_6301 = ~v_6252;
  assign v_6302 = v_6303 | v_6304;
  assign v_6303 = mux_6303(v_6254);
  assign v_6304 = mux_6304(v_6292);
  assign v_6306 = v_6307 | v_6345;
  assign v_6307 = act_6308 & 1'h1;
  assign act_6308 = v_6309 | v_6322;
  assign v_6309 = v_6310 & 1'h1;
  assign v_6310 = v_6311 & v_6329;
  assign v_6311 = ~v_6312;
  assign v_6313 = v_6314 | v_6316;
  assign v_6314 = act_6315 & 1'h1;
  assign act_6315 = v_596 | v_590;
  assign v_6316 = v_6317 & 1'h1;
  assign v_6317 = v_6318 & v_6319;
  assign v_6318 = ~act_6315;
  assign v_6319 = v_6320 | v_6325;
  assign v_6320 = v_6321 | v_6323;
  assign v_6321 = mux_6321(v_6322);
  assign v_6322 = v_6312 & 1'h1;
  assign v_6323 = mux_6323(v_6324);
  assign v_6324 = ~v_6322;
  assign v_6325 = ~v_6312;
  assign v_6326 = v_6327 | v_6328;
  assign v_6327 = mux_6327(v_6314);
  assign v_6328 = mux_6328(v_6316);
  assign v_6330 = v_6331 | v_6333;
  assign v_6331 = act_6332 & 1'h1;
  assign act_6332 = v_610 | v_604;
  assign v_6333 = v_6334 & 1'h1;
  assign v_6334 = v_6335 & v_6336;
  assign v_6335 = ~act_6332;
  assign v_6336 = v_6337 | v_6341;
  assign v_6337 = v_6338 | v_6339;
  assign v_6338 = mux_6338(v_6309);
  assign v_6339 = mux_6339(v_6340);
  assign v_6340 = ~v_6309;
  assign v_6341 = ~v_6329;
  assign v_6342 = v_6343 | v_6344;
  assign v_6343 = mux_6343(v_6331);
  assign v_6344 = mux_6344(v_6333);
  assign v_6345 = v_6346 & 1'h1;
  assign v_6346 = v_6347 & v_6348;
  assign v_6347 = ~act_6308;
  assign v_6348 = v_6349 | v_6353;
  assign v_6349 = v_6350 | v_6351;
  assign v_6350 = mux_6350(v_6249);
  assign v_6351 = mux_6351(v_6352);
  assign v_6352 = ~v_6249;
  assign v_6353 = ~v_6305;
  assign v_6354 = v_6355 | v_6356;
  assign v_6355 = mux_6355(v_6307);
  assign v_6356 = mux_6356(v_6345);
  assign v_6357 = v_6358 & 1'h1;
  assign v_6358 = v_6359 & v_6360;
  assign v_6359 = ~act_6248;
  assign v_6360 = v_6361 | v_6366;
  assign v_6361 = v_6362 | v_6364;
  assign v_6362 = mux_6362(v_6363);
  assign v_6363 = v_6245 & 1'h1;
  assign v_6364 = mux_6364(v_6365);
  assign v_6365 = ~v_6363;
  assign v_6366 = ~v_6245;
  assign v_6367 = v_6368 | v_6369;
  assign v_6368 = mux_6368(v_6247);
  assign v_6369 = mux_6369(v_6357);
  assign v_6371 = v_6372 | v_6482;
  assign v_6372 = act_6373 & 1'h1;
  assign act_6373 = v_6374 | v_6423;
  assign v_6374 = v_6375 & 1'h1;
  assign v_6375 = v_6376 & v_6430;
  assign v_6376 = ~v_6377;
  assign v_6378 = v_6379 | v_6417;
  assign v_6379 = act_6380 & 1'h1;
  assign act_6380 = v_6381 | v_6394;
  assign v_6381 = v_6382 & 1'h1;
  assign v_6382 = v_6383 & v_6401;
  assign v_6383 = ~v_6384;
  assign v_6385 = v_6386 | v_6388;
  assign v_6386 = act_6387 & 1'h1;
  assign act_6387 = v_624 | v_618;
  assign v_6388 = v_6389 & 1'h1;
  assign v_6389 = v_6390 & v_6391;
  assign v_6390 = ~act_6387;
  assign v_6391 = v_6392 | v_6397;
  assign v_6392 = v_6393 | v_6395;
  assign v_6393 = mux_6393(v_6394);
  assign v_6394 = v_6384 & 1'h1;
  assign v_6395 = mux_6395(v_6396);
  assign v_6396 = ~v_6394;
  assign v_6397 = ~v_6384;
  assign v_6398 = v_6399 | v_6400;
  assign v_6399 = mux_6399(v_6386);
  assign v_6400 = mux_6400(v_6388);
  assign v_6402 = v_6403 | v_6405;
  assign v_6403 = act_6404 & 1'h1;
  assign act_6404 = v_638 | v_632;
  assign v_6405 = v_6406 & 1'h1;
  assign v_6406 = v_6407 & v_6408;
  assign v_6407 = ~act_6404;
  assign v_6408 = v_6409 | v_6413;
  assign v_6409 = v_6410 | v_6411;
  assign v_6410 = mux_6410(v_6381);
  assign v_6411 = mux_6411(v_6412);
  assign v_6412 = ~v_6381;
  assign v_6413 = ~v_6401;
  assign v_6414 = v_6415 | v_6416;
  assign v_6415 = mux_6415(v_6403);
  assign v_6416 = mux_6416(v_6405);
  assign v_6417 = v_6418 & 1'h1;
  assign v_6418 = v_6419 & v_6420;
  assign v_6419 = ~act_6380;
  assign v_6420 = v_6421 | v_6426;
  assign v_6421 = v_6422 | v_6424;
  assign v_6422 = mux_6422(v_6423);
  assign v_6423 = v_6377 & 1'h1;
  assign v_6424 = mux_6424(v_6425);
  assign v_6425 = ~v_6423;
  assign v_6426 = ~v_6377;
  assign v_6427 = v_6428 | v_6429;
  assign v_6428 = mux_6428(v_6379);
  assign v_6429 = mux_6429(v_6417);
  assign v_6431 = v_6432 | v_6470;
  assign v_6432 = act_6433 & 1'h1;
  assign act_6433 = v_6434 | v_6447;
  assign v_6434 = v_6435 & 1'h1;
  assign v_6435 = v_6436 & v_6454;
  assign v_6436 = ~v_6437;
  assign v_6438 = v_6439 | v_6441;
  assign v_6439 = act_6440 & 1'h1;
  assign act_6440 = v_652 | v_646;
  assign v_6441 = v_6442 & 1'h1;
  assign v_6442 = v_6443 & v_6444;
  assign v_6443 = ~act_6440;
  assign v_6444 = v_6445 | v_6450;
  assign v_6445 = v_6446 | v_6448;
  assign v_6446 = mux_6446(v_6447);
  assign v_6447 = v_6437 & 1'h1;
  assign v_6448 = mux_6448(v_6449);
  assign v_6449 = ~v_6447;
  assign v_6450 = ~v_6437;
  assign v_6451 = v_6452 | v_6453;
  assign v_6452 = mux_6452(v_6439);
  assign v_6453 = mux_6453(v_6441);
  assign v_6455 = v_6456 | v_6458;
  assign v_6456 = act_6457 & 1'h1;
  assign act_6457 = v_666 | v_660;
  assign v_6458 = v_6459 & 1'h1;
  assign v_6459 = v_6460 & v_6461;
  assign v_6460 = ~act_6457;
  assign v_6461 = v_6462 | v_6466;
  assign v_6462 = v_6463 | v_6464;
  assign v_6463 = mux_6463(v_6434);
  assign v_6464 = mux_6464(v_6465);
  assign v_6465 = ~v_6434;
  assign v_6466 = ~v_6454;
  assign v_6467 = v_6468 | v_6469;
  assign v_6468 = mux_6468(v_6456);
  assign v_6469 = mux_6469(v_6458);
  assign v_6470 = v_6471 & 1'h1;
  assign v_6471 = v_6472 & v_6473;
  assign v_6472 = ~act_6433;
  assign v_6473 = v_6474 | v_6478;
  assign v_6474 = v_6475 | v_6476;
  assign v_6475 = mux_6475(v_6374);
  assign v_6476 = mux_6476(v_6477);
  assign v_6477 = ~v_6374;
  assign v_6478 = ~v_6430;
  assign v_6479 = v_6480 | v_6481;
  assign v_6480 = mux_6480(v_6432);
  assign v_6481 = mux_6481(v_6470);
  assign v_6482 = v_6483 & 1'h1;
  assign v_6483 = v_6484 & v_6485;
  assign v_6484 = ~act_6373;
  assign v_6485 = v_6486 | v_6490;
  assign v_6486 = v_6487 | v_6488;
  assign v_6487 = mux_6487(v_6242);
  assign v_6488 = mux_6488(v_6489);
  assign v_6489 = ~v_6242;
  assign v_6490 = ~v_6370;
  assign v_6491 = v_6492 | v_6493;
  assign v_6492 = mux_6492(v_6372);
  assign v_6493 = mux_6493(v_6482);
  assign v_6494 = v_6495 & 1'h1;
  assign v_6495 = v_6496 & v_6497;
  assign v_6496 = ~act_6241;
  assign v_6497 = v_6498 | v_6502;
  assign v_6498 = v_6499 | v_6500;
  assign v_6499 = mux_6499(v_5966);
  assign v_6500 = mux_6500(v_6501);
  assign v_6501 = ~v_5966;
  assign v_6502 = ~v_6238;
  assign v_6503 = v_6504 | v_6505;
  assign v_6504 = mux_6504(v_6240);
  assign v_6505 = mux_6505(v_6494);
  assign v_6506 = v_6507 & 1'h1;
  assign v_6507 = v_6508 & v_6509;
  assign v_6508 = ~act_5965;
  assign v_6509 = v_6510 | v_6514;
  assign v_6510 = v_6511 | v_6512;
  assign v_6511 = mux_6511(v_5402);
  assign v_6512 = mux_6512(v_6513);
  assign v_6513 = ~v_5402;
  assign v_6514 = ~v_5962;
  assign v_6515 = v_6516 | v_6517;
  assign v_6516 = mux_6516(v_5964);
  assign v_6517 = mux_6517(v_6506);
  assign v_6518 = v_6519 & 1'h1;
  assign v_6519 = v_6520 & v_6521;
  assign v_6520 = ~act_5401;
  assign v_6521 = v_6522 | v_6527;
  assign v_6522 = v_6523 | v_6525;
  assign v_6523 = mux_6523(v_6524);
  assign v_6524 = v_5398 & 1'h1;
  assign v_6525 = mux_6525(v_6526);
  assign v_6526 = ~v_6524;
  assign v_6527 = ~v_5398;
  assign v_6528 = v_6529 | v_6530;
  assign v_6529 = mux_6529(v_5400);
  assign v_6530 = mux_6530(v_6518);
  assign v_6532 = v_6533 | v_7651;
  assign v_6533 = act_6534 & 1'h1;
  assign act_6534 = v_6535 | v_7088;
  assign v_6535 = v_6536 & 1'h1;
  assign v_6536 = v_6537 & v_7095;
  assign v_6537 = ~v_6538;
  assign v_6539 = v_6540 | v_7082;
  assign v_6540 = act_6541 & 1'h1;
  assign act_6541 = v_6542 | v_6807;
  assign v_6542 = v_6543 & 1'h1;
  assign v_6543 = v_6544 & v_6814;
  assign v_6544 = ~v_6545;
  assign v_6546 = v_6547 | v_6801;
  assign v_6547 = act_6548 & 1'h1;
  assign act_6548 = v_6549 | v_6670;
  assign v_6549 = v_6550 & 1'h1;
  assign v_6550 = v_6551 & v_6677;
  assign v_6551 = ~v_6552;
  assign v_6553 = v_6554 | v_6664;
  assign v_6554 = act_6555 & 1'h1;
  assign act_6555 = v_6556 | v_6605;
  assign v_6556 = v_6557 & 1'h1;
  assign v_6557 = v_6558 & v_6612;
  assign v_6558 = ~v_6559;
  assign v_6560 = v_6561 | v_6599;
  assign v_6561 = act_6562 & 1'h1;
  assign act_6562 = v_6563 | v_6576;
  assign v_6563 = v_6564 & 1'h1;
  assign v_6564 = v_6565 & v_6583;
  assign v_6565 = ~v_6566;
  assign v_6567 = v_6568 | v_6570;
  assign v_6568 = act_6569 & 1'h1;
  assign act_6569 = v_680 | v_674;
  assign v_6570 = v_6571 & 1'h1;
  assign v_6571 = v_6572 & v_6573;
  assign v_6572 = ~act_6569;
  assign v_6573 = v_6574 | v_6579;
  assign v_6574 = v_6575 | v_6577;
  assign v_6575 = mux_6575(v_6576);
  assign v_6576 = v_6566 & 1'h1;
  assign v_6577 = mux_6577(v_6578);
  assign v_6578 = ~v_6576;
  assign v_6579 = ~v_6566;
  assign v_6580 = v_6581 | v_6582;
  assign v_6581 = mux_6581(v_6568);
  assign v_6582 = mux_6582(v_6570);
  assign v_6584 = v_6585 | v_6587;
  assign v_6585 = act_6586 & 1'h1;
  assign act_6586 = v_694 | v_688;
  assign v_6587 = v_6588 & 1'h1;
  assign v_6588 = v_6589 & v_6590;
  assign v_6589 = ~act_6586;
  assign v_6590 = v_6591 | v_6595;
  assign v_6591 = v_6592 | v_6593;
  assign v_6592 = mux_6592(v_6563);
  assign v_6593 = mux_6593(v_6594);
  assign v_6594 = ~v_6563;
  assign v_6595 = ~v_6583;
  assign v_6596 = v_6597 | v_6598;
  assign v_6597 = mux_6597(v_6585);
  assign v_6598 = mux_6598(v_6587);
  assign v_6599 = v_6600 & 1'h1;
  assign v_6600 = v_6601 & v_6602;
  assign v_6601 = ~act_6562;
  assign v_6602 = v_6603 | v_6608;
  assign v_6603 = v_6604 | v_6606;
  assign v_6604 = mux_6604(v_6605);
  assign v_6605 = v_6559 & 1'h1;
  assign v_6606 = mux_6606(v_6607);
  assign v_6607 = ~v_6605;
  assign v_6608 = ~v_6559;
  assign v_6609 = v_6610 | v_6611;
  assign v_6610 = mux_6610(v_6561);
  assign v_6611 = mux_6611(v_6599);
  assign v_6613 = v_6614 | v_6652;
  assign v_6614 = act_6615 & 1'h1;
  assign act_6615 = v_6616 | v_6629;
  assign v_6616 = v_6617 & 1'h1;
  assign v_6617 = v_6618 & v_6636;
  assign v_6618 = ~v_6619;
  assign v_6620 = v_6621 | v_6623;
  assign v_6621 = act_6622 & 1'h1;
  assign act_6622 = v_708 | v_702;
  assign v_6623 = v_6624 & 1'h1;
  assign v_6624 = v_6625 & v_6626;
  assign v_6625 = ~act_6622;
  assign v_6626 = v_6627 | v_6632;
  assign v_6627 = v_6628 | v_6630;
  assign v_6628 = mux_6628(v_6629);
  assign v_6629 = v_6619 & 1'h1;
  assign v_6630 = mux_6630(v_6631);
  assign v_6631 = ~v_6629;
  assign v_6632 = ~v_6619;
  assign v_6633 = v_6634 | v_6635;
  assign v_6634 = mux_6634(v_6621);
  assign v_6635 = mux_6635(v_6623);
  assign v_6637 = v_6638 | v_6640;
  assign v_6638 = act_6639 & 1'h1;
  assign act_6639 = v_722 | v_716;
  assign v_6640 = v_6641 & 1'h1;
  assign v_6641 = v_6642 & v_6643;
  assign v_6642 = ~act_6639;
  assign v_6643 = v_6644 | v_6648;
  assign v_6644 = v_6645 | v_6646;
  assign v_6645 = mux_6645(v_6616);
  assign v_6646 = mux_6646(v_6647);
  assign v_6647 = ~v_6616;
  assign v_6648 = ~v_6636;
  assign v_6649 = v_6650 | v_6651;
  assign v_6650 = mux_6650(v_6638);
  assign v_6651 = mux_6651(v_6640);
  assign v_6652 = v_6653 & 1'h1;
  assign v_6653 = v_6654 & v_6655;
  assign v_6654 = ~act_6615;
  assign v_6655 = v_6656 | v_6660;
  assign v_6656 = v_6657 | v_6658;
  assign v_6657 = mux_6657(v_6556);
  assign v_6658 = mux_6658(v_6659);
  assign v_6659 = ~v_6556;
  assign v_6660 = ~v_6612;
  assign v_6661 = v_6662 | v_6663;
  assign v_6662 = mux_6662(v_6614);
  assign v_6663 = mux_6663(v_6652);
  assign v_6664 = v_6665 & 1'h1;
  assign v_6665 = v_6666 & v_6667;
  assign v_6666 = ~act_6555;
  assign v_6667 = v_6668 | v_6673;
  assign v_6668 = v_6669 | v_6671;
  assign v_6669 = mux_6669(v_6670);
  assign v_6670 = v_6552 & 1'h1;
  assign v_6671 = mux_6671(v_6672);
  assign v_6672 = ~v_6670;
  assign v_6673 = ~v_6552;
  assign v_6674 = v_6675 | v_6676;
  assign v_6675 = mux_6675(v_6554);
  assign v_6676 = mux_6676(v_6664);
  assign v_6678 = v_6679 | v_6789;
  assign v_6679 = act_6680 & 1'h1;
  assign act_6680 = v_6681 | v_6730;
  assign v_6681 = v_6682 & 1'h1;
  assign v_6682 = v_6683 & v_6737;
  assign v_6683 = ~v_6684;
  assign v_6685 = v_6686 | v_6724;
  assign v_6686 = act_6687 & 1'h1;
  assign act_6687 = v_6688 | v_6701;
  assign v_6688 = v_6689 & 1'h1;
  assign v_6689 = v_6690 & v_6708;
  assign v_6690 = ~v_6691;
  assign v_6692 = v_6693 | v_6695;
  assign v_6693 = act_6694 & 1'h1;
  assign act_6694 = v_736 | v_730;
  assign v_6695 = v_6696 & 1'h1;
  assign v_6696 = v_6697 & v_6698;
  assign v_6697 = ~act_6694;
  assign v_6698 = v_6699 | v_6704;
  assign v_6699 = v_6700 | v_6702;
  assign v_6700 = mux_6700(v_6701);
  assign v_6701 = v_6691 & 1'h1;
  assign v_6702 = mux_6702(v_6703);
  assign v_6703 = ~v_6701;
  assign v_6704 = ~v_6691;
  assign v_6705 = v_6706 | v_6707;
  assign v_6706 = mux_6706(v_6693);
  assign v_6707 = mux_6707(v_6695);
  assign v_6709 = v_6710 | v_6712;
  assign v_6710 = act_6711 & 1'h1;
  assign act_6711 = v_750 | v_744;
  assign v_6712 = v_6713 & 1'h1;
  assign v_6713 = v_6714 & v_6715;
  assign v_6714 = ~act_6711;
  assign v_6715 = v_6716 | v_6720;
  assign v_6716 = v_6717 | v_6718;
  assign v_6717 = mux_6717(v_6688);
  assign v_6718 = mux_6718(v_6719);
  assign v_6719 = ~v_6688;
  assign v_6720 = ~v_6708;
  assign v_6721 = v_6722 | v_6723;
  assign v_6722 = mux_6722(v_6710);
  assign v_6723 = mux_6723(v_6712);
  assign v_6724 = v_6725 & 1'h1;
  assign v_6725 = v_6726 & v_6727;
  assign v_6726 = ~act_6687;
  assign v_6727 = v_6728 | v_6733;
  assign v_6728 = v_6729 | v_6731;
  assign v_6729 = mux_6729(v_6730);
  assign v_6730 = v_6684 & 1'h1;
  assign v_6731 = mux_6731(v_6732);
  assign v_6732 = ~v_6730;
  assign v_6733 = ~v_6684;
  assign v_6734 = v_6735 | v_6736;
  assign v_6735 = mux_6735(v_6686);
  assign v_6736 = mux_6736(v_6724);
  assign v_6738 = v_6739 | v_6777;
  assign v_6739 = act_6740 & 1'h1;
  assign act_6740 = v_6741 | v_6754;
  assign v_6741 = v_6742 & 1'h1;
  assign v_6742 = v_6743 & v_6761;
  assign v_6743 = ~v_6744;
  assign v_6745 = v_6746 | v_6748;
  assign v_6746 = act_6747 & 1'h1;
  assign act_6747 = v_764 | v_758;
  assign v_6748 = v_6749 & 1'h1;
  assign v_6749 = v_6750 & v_6751;
  assign v_6750 = ~act_6747;
  assign v_6751 = v_6752 | v_6757;
  assign v_6752 = v_6753 | v_6755;
  assign v_6753 = mux_6753(v_6754);
  assign v_6754 = v_6744 & 1'h1;
  assign v_6755 = mux_6755(v_6756);
  assign v_6756 = ~v_6754;
  assign v_6757 = ~v_6744;
  assign v_6758 = v_6759 | v_6760;
  assign v_6759 = mux_6759(v_6746);
  assign v_6760 = mux_6760(v_6748);
  assign v_6762 = v_6763 | v_6765;
  assign v_6763 = act_6764 & 1'h1;
  assign act_6764 = v_778 | v_772;
  assign v_6765 = v_6766 & 1'h1;
  assign v_6766 = v_6767 & v_6768;
  assign v_6767 = ~act_6764;
  assign v_6768 = v_6769 | v_6773;
  assign v_6769 = v_6770 | v_6771;
  assign v_6770 = mux_6770(v_6741);
  assign v_6771 = mux_6771(v_6772);
  assign v_6772 = ~v_6741;
  assign v_6773 = ~v_6761;
  assign v_6774 = v_6775 | v_6776;
  assign v_6775 = mux_6775(v_6763);
  assign v_6776 = mux_6776(v_6765);
  assign v_6777 = v_6778 & 1'h1;
  assign v_6778 = v_6779 & v_6780;
  assign v_6779 = ~act_6740;
  assign v_6780 = v_6781 | v_6785;
  assign v_6781 = v_6782 | v_6783;
  assign v_6782 = mux_6782(v_6681);
  assign v_6783 = mux_6783(v_6784);
  assign v_6784 = ~v_6681;
  assign v_6785 = ~v_6737;
  assign v_6786 = v_6787 | v_6788;
  assign v_6787 = mux_6787(v_6739);
  assign v_6788 = mux_6788(v_6777);
  assign v_6789 = v_6790 & 1'h1;
  assign v_6790 = v_6791 & v_6792;
  assign v_6791 = ~act_6680;
  assign v_6792 = v_6793 | v_6797;
  assign v_6793 = v_6794 | v_6795;
  assign v_6794 = mux_6794(v_6549);
  assign v_6795 = mux_6795(v_6796);
  assign v_6796 = ~v_6549;
  assign v_6797 = ~v_6677;
  assign v_6798 = v_6799 | v_6800;
  assign v_6799 = mux_6799(v_6679);
  assign v_6800 = mux_6800(v_6789);
  assign v_6801 = v_6802 & 1'h1;
  assign v_6802 = v_6803 & v_6804;
  assign v_6803 = ~act_6548;
  assign v_6804 = v_6805 | v_6810;
  assign v_6805 = v_6806 | v_6808;
  assign v_6806 = mux_6806(v_6807);
  assign v_6807 = v_6545 & 1'h1;
  assign v_6808 = mux_6808(v_6809);
  assign v_6809 = ~v_6807;
  assign v_6810 = ~v_6545;
  assign v_6811 = v_6812 | v_6813;
  assign v_6812 = mux_6812(v_6547);
  assign v_6813 = mux_6813(v_6801);
  assign v_6815 = v_6816 | v_7070;
  assign v_6816 = act_6817 & 1'h1;
  assign act_6817 = v_6818 | v_6939;
  assign v_6818 = v_6819 & 1'h1;
  assign v_6819 = v_6820 & v_6946;
  assign v_6820 = ~v_6821;
  assign v_6822 = v_6823 | v_6933;
  assign v_6823 = act_6824 & 1'h1;
  assign act_6824 = v_6825 | v_6874;
  assign v_6825 = v_6826 & 1'h1;
  assign v_6826 = v_6827 & v_6881;
  assign v_6827 = ~v_6828;
  assign v_6829 = v_6830 | v_6868;
  assign v_6830 = act_6831 & 1'h1;
  assign act_6831 = v_6832 | v_6845;
  assign v_6832 = v_6833 & 1'h1;
  assign v_6833 = v_6834 & v_6852;
  assign v_6834 = ~v_6835;
  assign v_6836 = v_6837 | v_6839;
  assign v_6837 = act_6838 & 1'h1;
  assign act_6838 = v_792 | v_786;
  assign v_6839 = v_6840 & 1'h1;
  assign v_6840 = v_6841 & v_6842;
  assign v_6841 = ~act_6838;
  assign v_6842 = v_6843 | v_6848;
  assign v_6843 = v_6844 | v_6846;
  assign v_6844 = mux_6844(v_6845);
  assign v_6845 = v_6835 & 1'h1;
  assign v_6846 = mux_6846(v_6847);
  assign v_6847 = ~v_6845;
  assign v_6848 = ~v_6835;
  assign v_6849 = v_6850 | v_6851;
  assign v_6850 = mux_6850(v_6837);
  assign v_6851 = mux_6851(v_6839);
  assign v_6853 = v_6854 | v_6856;
  assign v_6854 = act_6855 & 1'h1;
  assign act_6855 = v_806 | v_800;
  assign v_6856 = v_6857 & 1'h1;
  assign v_6857 = v_6858 & v_6859;
  assign v_6858 = ~act_6855;
  assign v_6859 = v_6860 | v_6864;
  assign v_6860 = v_6861 | v_6862;
  assign v_6861 = mux_6861(v_6832);
  assign v_6862 = mux_6862(v_6863);
  assign v_6863 = ~v_6832;
  assign v_6864 = ~v_6852;
  assign v_6865 = v_6866 | v_6867;
  assign v_6866 = mux_6866(v_6854);
  assign v_6867 = mux_6867(v_6856);
  assign v_6868 = v_6869 & 1'h1;
  assign v_6869 = v_6870 & v_6871;
  assign v_6870 = ~act_6831;
  assign v_6871 = v_6872 | v_6877;
  assign v_6872 = v_6873 | v_6875;
  assign v_6873 = mux_6873(v_6874);
  assign v_6874 = v_6828 & 1'h1;
  assign v_6875 = mux_6875(v_6876);
  assign v_6876 = ~v_6874;
  assign v_6877 = ~v_6828;
  assign v_6878 = v_6879 | v_6880;
  assign v_6879 = mux_6879(v_6830);
  assign v_6880 = mux_6880(v_6868);
  assign v_6882 = v_6883 | v_6921;
  assign v_6883 = act_6884 & 1'h1;
  assign act_6884 = v_6885 | v_6898;
  assign v_6885 = v_6886 & 1'h1;
  assign v_6886 = v_6887 & v_6905;
  assign v_6887 = ~v_6888;
  assign v_6889 = v_6890 | v_6892;
  assign v_6890 = act_6891 & 1'h1;
  assign act_6891 = v_820 | v_814;
  assign v_6892 = v_6893 & 1'h1;
  assign v_6893 = v_6894 & v_6895;
  assign v_6894 = ~act_6891;
  assign v_6895 = v_6896 | v_6901;
  assign v_6896 = v_6897 | v_6899;
  assign v_6897 = mux_6897(v_6898);
  assign v_6898 = v_6888 & 1'h1;
  assign v_6899 = mux_6899(v_6900);
  assign v_6900 = ~v_6898;
  assign v_6901 = ~v_6888;
  assign v_6902 = v_6903 | v_6904;
  assign v_6903 = mux_6903(v_6890);
  assign v_6904 = mux_6904(v_6892);
  assign v_6906 = v_6907 | v_6909;
  assign v_6907 = act_6908 & 1'h1;
  assign act_6908 = v_834 | v_828;
  assign v_6909 = v_6910 & 1'h1;
  assign v_6910 = v_6911 & v_6912;
  assign v_6911 = ~act_6908;
  assign v_6912 = v_6913 | v_6917;
  assign v_6913 = v_6914 | v_6915;
  assign v_6914 = mux_6914(v_6885);
  assign v_6915 = mux_6915(v_6916);
  assign v_6916 = ~v_6885;
  assign v_6917 = ~v_6905;
  assign v_6918 = v_6919 | v_6920;
  assign v_6919 = mux_6919(v_6907);
  assign v_6920 = mux_6920(v_6909);
  assign v_6921 = v_6922 & 1'h1;
  assign v_6922 = v_6923 & v_6924;
  assign v_6923 = ~act_6884;
  assign v_6924 = v_6925 | v_6929;
  assign v_6925 = v_6926 | v_6927;
  assign v_6926 = mux_6926(v_6825);
  assign v_6927 = mux_6927(v_6928);
  assign v_6928 = ~v_6825;
  assign v_6929 = ~v_6881;
  assign v_6930 = v_6931 | v_6932;
  assign v_6931 = mux_6931(v_6883);
  assign v_6932 = mux_6932(v_6921);
  assign v_6933 = v_6934 & 1'h1;
  assign v_6934 = v_6935 & v_6936;
  assign v_6935 = ~act_6824;
  assign v_6936 = v_6937 | v_6942;
  assign v_6937 = v_6938 | v_6940;
  assign v_6938 = mux_6938(v_6939);
  assign v_6939 = v_6821 & 1'h1;
  assign v_6940 = mux_6940(v_6941);
  assign v_6941 = ~v_6939;
  assign v_6942 = ~v_6821;
  assign v_6943 = v_6944 | v_6945;
  assign v_6944 = mux_6944(v_6823);
  assign v_6945 = mux_6945(v_6933);
  assign v_6947 = v_6948 | v_7058;
  assign v_6948 = act_6949 & 1'h1;
  assign act_6949 = v_6950 | v_6999;
  assign v_6950 = v_6951 & 1'h1;
  assign v_6951 = v_6952 & v_7006;
  assign v_6952 = ~v_6953;
  assign v_6954 = v_6955 | v_6993;
  assign v_6955 = act_6956 & 1'h1;
  assign act_6956 = v_6957 | v_6970;
  assign v_6957 = v_6958 & 1'h1;
  assign v_6958 = v_6959 & v_6977;
  assign v_6959 = ~v_6960;
  assign v_6961 = v_6962 | v_6964;
  assign v_6962 = act_6963 & 1'h1;
  assign act_6963 = v_848 | v_842;
  assign v_6964 = v_6965 & 1'h1;
  assign v_6965 = v_6966 & v_6967;
  assign v_6966 = ~act_6963;
  assign v_6967 = v_6968 | v_6973;
  assign v_6968 = v_6969 | v_6971;
  assign v_6969 = mux_6969(v_6970);
  assign v_6970 = v_6960 & 1'h1;
  assign v_6971 = mux_6971(v_6972);
  assign v_6972 = ~v_6970;
  assign v_6973 = ~v_6960;
  assign v_6974 = v_6975 | v_6976;
  assign v_6975 = mux_6975(v_6962);
  assign v_6976 = mux_6976(v_6964);
  assign v_6978 = v_6979 | v_6981;
  assign v_6979 = act_6980 & 1'h1;
  assign act_6980 = v_862 | v_856;
  assign v_6981 = v_6982 & 1'h1;
  assign v_6982 = v_6983 & v_6984;
  assign v_6983 = ~act_6980;
  assign v_6984 = v_6985 | v_6989;
  assign v_6985 = v_6986 | v_6987;
  assign v_6986 = mux_6986(v_6957);
  assign v_6987 = mux_6987(v_6988);
  assign v_6988 = ~v_6957;
  assign v_6989 = ~v_6977;
  assign v_6990 = v_6991 | v_6992;
  assign v_6991 = mux_6991(v_6979);
  assign v_6992 = mux_6992(v_6981);
  assign v_6993 = v_6994 & 1'h1;
  assign v_6994 = v_6995 & v_6996;
  assign v_6995 = ~act_6956;
  assign v_6996 = v_6997 | v_7002;
  assign v_6997 = v_6998 | v_7000;
  assign v_6998 = mux_6998(v_6999);
  assign v_6999 = v_6953 & 1'h1;
  assign v_7000 = mux_7000(v_7001);
  assign v_7001 = ~v_6999;
  assign v_7002 = ~v_6953;
  assign v_7003 = v_7004 | v_7005;
  assign v_7004 = mux_7004(v_6955);
  assign v_7005 = mux_7005(v_6993);
  assign v_7007 = v_7008 | v_7046;
  assign v_7008 = act_7009 & 1'h1;
  assign act_7009 = v_7010 | v_7023;
  assign v_7010 = v_7011 & 1'h1;
  assign v_7011 = v_7012 & v_7030;
  assign v_7012 = ~v_7013;
  assign v_7014 = v_7015 | v_7017;
  assign v_7015 = act_7016 & 1'h1;
  assign act_7016 = v_876 | v_870;
  assign v_7017 = v_7018 & 1'h1;
  assign v_7018 = v_7019 & v_7020;
  assign v_7019 = ~act_7016;
  assign v_7020 = v_7021 | v_7026;
  assign v_7021 = v_7022 | v_7024;
  assign v_7022 = mux_7022(v_7023);
  assign v_7023 = v_7013 & 1'h1;
  assign v_7024 = mux_7024(v_7025);
  assign v_7025 = ~v_7023;
  assign v_7026 = ~v_7013;
  assign v_7027 = v_7028 | v_7029;
  assign v_7028 = mux_7028(v_7015);
  assign v_7029 = mux_7029(v_7017);
  assign v_7031 = v_7032 | v_7034;
  assign v_7032 = act_7033 & 1'h1;
  assign act_7033 = v_890 | v_884;
  assign v_7034 = v_7035 & 1'h1;
  assign v_7035 = v_7036 & v_7037;
  assign v_7036 = ~act_7033;
  assign v_7037 = v_7038 | v_7042;
  assign v_7038 = v_7039 | v_7040;
  assign v_7039 = mux_7039(v_7010);
  assign v_7040 = mux_7040(v_7041);
  assign v_7041 = ~v_7010;
  assign v_7042 = ~v_7030;
  assign v_7043 = v_7044 | v_7045;
  assign v_7044 = mux_7044(v_7032);
  assign v_7045 = mux_7045(v_7034);
  assign v_7046 = v_7047 & 1'h1;
  assign v_7047 = v_7048 & v_7049;
  assign v_7048 = ~act_7009;
  assign v_7049 = v_7050 | v_7054;
  assign v_7050 = v_7051 | v_7052;
  assign v_7051 = mux_7051(v_6950);
  assign v_7052 = mux_7052(v_7053);
  assign v_7053 = ~v_6950;
  assign v_7054 = ~v_7006;
  assign v_7055 = v_7056 | v_7057;
  assign v_7056 = mux_7056(v_7008);
  assign v_7057 = mux_7057(v_7046);
  assign v_7058 = v_7059 & 1'h1;
  assign v_7059 = v_7060 & v_7061;
  assign v_7060 = ~act_6949;
  assign v_7061 = v_7062 | v_7066;
  assign v_7062 = v_7063 | v_7064;
  assign v_7063 = mux_7063(v_6818);
  assign v_7064 = mux_7064(v_7065);
  assign v_7065 = ~v_6818;
  assign v_7066 = ~v_6946;
  assign v_7067 = v_7068 | v_7069;
  assign v_7068 = mux_7068(v_6948);
  assign v_7069 = mux_7069(v_7058);
  assign v_7070 = v_7071 & 1'h1;
  assign v_7071 = v_7072 & v_7073;
  assign v_7072 = ~act_6817;
  assign v_7073 = v_7074 | v_7078;
  assign v_7074 = v_7075 | v_7076;
  assign v_7075 = mux_7075(v_6542);
  assign v_7076 = mux_7076(v_7077);
  assign v_7077 = ~v_6542;
  assign v_7078 = ~v_6814;
  assign v_7079 = v_7080 | v_7081;
  assign v_7080 = mux_7080(v_6816);
  assign v_7081 = mux_7081(v_7070);
  assign v_7082 = v_7083 & 1'h1;
  assign v_7083 = v_7084 & v_7085;
  assign v_7084 = ~act_6541;
  assign v_7085 = v_7086 | v_7091;
  assign v_7086 = v_7087 | v_7089;
  assign v_7087 = mux_7087(v_7088);
  assign v_7088 = v_6538 & 1'h1;
  assign v_7089 = mux_7089(v_7090);
  assign v_7090 = ~v_7088;
  assign v_7091 = ~v_6538;
  assign v_7092 = v_7093 | v_7094;
  assign v_7093 = mux_7093(v_6540);
  assign v_7094 = mux_7094(v_7082);
  assign v_7096 = v_7097 | v_7639;
  assign v_7097 = act_7098 & 1'h1;
  assign act_7098 = v_7099 | v_7364;
  assign v_7099 = v_7100 & 1'h1;
  assign v_7100 = v_7101 & v_7371;
  assign v_7101 = ~v_7102;
  assign v_7103 = v_7104 | v_7358;
  assign v_7104 = act_7105 & 1'h1;
  assign act_7105 = v_7106 | v_7227;
  assign v_7106 = v_7107 & 1'h1;
  assign v_7107 = v_7108 & v_7234;
  assign v_7108 = ~v_7109;
  assign v_7110 = v_7111 | v_7221;
  assign v_7111 = act_7112 & 1'h1;
  assign act_7112 = v_7113 | v_7162;
  assign v_7113 = v_7114 & 1'h1;
  assign v_7114 = v_7115 & v_7169;
  assign v_7115 = ~v_7116;
  assign v_7117 = v_7118 | v_7156;
  assign v_7118 = act_7119 & 1'h1;
  assign act_7119 = v_7120 | v_7133;
  assign v_7120 = v_7121 & 1'h1;
  assign v_7121 = v_7122 & v_7140;
  assign v_7122 = ~v_7123;
  assign v_7124 = v_7125 | v_7127;
  assign v_7125 = act_7126 & 1'h1;
  assign act_7126 = v_904 | v_898;
  assign v_7127 = v_7128 & 1'h1;
  assign v_7128 = v_7129 & v_7130;
  assign v_7129 = ~act_7126;
  assign v_7130 = v_7131 | v_7136;
  assign v_7131 = v_7132 | v_7134;
  assign v_7132 = mux_7132(v_7133);
  assign v_7133 = v_7123 & 1'h1;
  assign v_7134 = mux_7134(v_7135);
  assign v_7135 = ~v_7133;
  assign v_7136 = ~v_7123;
  assign v_7137 = v_7138 | v_7139;
  assign v_7138 = mux_7138(v_7125);
  assign v_7139 = mux_7139(v_7127);
  assign v_7141 = v_7142 | v_7144;
  assign v_7142 = act_7143 & 1'h1;
  assign act_7143 = v_918 | v_912;
  assign v_7144 = v_7145 & 1'h1;
  assign v_7145 = v_7146 & v_7147;
  assign v_7146 = ~act_7143;
  assign v_7147 = v_7148 | v_7152;
  assign v_7148 = v_7149 | v_7150;
  assign v_7149 = mux_7149(v_7120);
  assign v_7150 = mux_7150(v_7151);
  assign v_7151 = ~v_7120;
  assign v_7152 = ~v_7140;
  assign v_7153 = v_7154 | v_7155;
  assign v_7154 = mux_7154(v_7142);
  assign v_7155 = mux_7155(v_7144);
  assign v_7156 = v_7157 & 1'h1;
  assign v_7157 = v_7158 & v_7159;
  assign v_7158 = ~act_7119;
  assign v_7159 = v_7160 | v_7165;
  assign v_7160 = v_7161 | v_7163;
  assign v_7161 = mux_7161(v_7162);
  assign v_7162 = v_7116 & 1'h1;
  assign v_7163 = mux_7163(v_7164);
  assign v_7164 = ~v_7162;
  assign v_7165 = ~v_7116;
  assign v_7166 = v_7167 | v_7168;
  assign v_7167 = mux_7167(v_7118);
  assign v_7168 = mux_7168(v_7156);
  assign v_7170 = v_7171 | v_7209;
  assign v_7171 = act_7172 & 1'h1;
  assign act_7172 = v_7173 | v_7186;
  assign v_7173 = v_7174 & 1'h1;
  assign v_7174 = v_7175 & v_7193;
  assign v_7175 = ~v_7176;
  assign v_7177 = v_7178 | v_7180;
  assign v_7178 = act_7179 & 1'h1;
  assign act_7179 = v_932 | v_926;
  assign v_7180 = v_7181 & 1'h1;
  assign v_7181 = v_7182 & v_7183;
  assign v_7182 = ~act_7179;
  assign v_7183 = v_7184 | v_7189;
  assign v_7184 = v_7185 | v_7187;
  assign v_7185 = mux_7185(v_7186);
  assign v_7186 = v_7176 & 1'h1;
  assign v_7187 = mux_7187(v_7188);
  assign v_7188 = ~v_7186;
  assign v_7189 = ~v_7176;
  assign v_7190 = v_7191 | v_7192;
  assign v_7191 = mux_7191(v_7178);
  assign v_7192 = mux_7192(v_7180);
  assign v_7194 = v_7195 | v_7197;
  assign v_7195 = act_7196 & 1'h1;
  assign act_7196 = v_946 | v_940;
  assign v_7197 = v_7198 & 1'h1;
  assign v_7198 = v_7199 & v_7200;
  assign v_7199 = ~act_7196;
  assign v_7200 = v_7201 | v_7205;
  assign v_7201 = v_7202 | v_7203;
  assign v_7202 = mux_7202(v_7173);
  assign v_7203 = mux_7203(v_7204);
  assign v_7204 = ~v_7173;
  assign v_7205 = ~v_7193;
  assign v_7206 = v_7207 | v_7208;
  assign v_7207 = mux_7207(v_7195);
  assign v_7208 = mux_7208(v_7197);
  assign v_7209 = v_7210 & 1'h1;
  assign v_7210 = v_7211 & v_7212;
  assign v_7211 = ~act_7172;
  assign v_7212 = v_7213 | v_7217;
  assign v_7213 = v_7214 | v_7215;
  assign v_7214 = mux_7214(v_7113);
  assign v_7215 = mux_7215(v_7216);
  assign v_7216 = ~v_7113;
  assign v_7217 = ~v_7169;
  assign v_7218 = v_7219 | v_7220;
  assign v_7219 = mux_7219(v_7171);
  assign v_7220 = mux_7220(v_7209);
  assign v_7221 = v_7222 & 1'h1;
  assign v_7222 = v_7223 & v_7224;
  assign v_7223 = ~act_7112;
  assign v_7224 = v_7225 | v_7230;
  assign v_7225 = v_7226 | v_7228;
  assign v_7226 = mux_7226(v_7227);
  assign v_7227 = v_7109 & 1'h1;
  assign v_7228 = mux_7228(v_7229);
  assign v_7229 = ~v_7227;
  assign v_7230 = ~v_7109;
  assign v_7231 = v_7232 | v_7233;
  assign v_7232 = mux_7232(v_7111);
  assign v_7233 = mux_7233(v_7221);
  assign v_7235 = v_7236 | v_7346;
  assign v_7236 = act_7237 & 1'h1;
  assign act_7237 = v_7238 | v_7287;
  assign v_7238 = v_7239 & 1'h1;
  assign v_7239 = v_7240 & v_7294;
  assign v_7240 = ~v_7241;
  assign v_7242 = v_7243 | v_7281;
  assign v_7243 = act_7244 & 1'h1;
  assign act_7244 = v_7245 | v_7258;
  assign v_7245 = v_7246 & 1'h1;
  assign v_7246 = v_7247 & v_7265;
  assign v_7247 = ~v_7248;
  assign v_7249 = v_7250 | v_7252;
  assign v_7250 = act_7251 & 1'h1;
  assign act_7251 = v_960 | v_954;
  assign v_7252 = v_7253 & 1'h1;
  assign v_7253 = v_7254 & v_7255;
  assign v_7254 = ~act_7251;
  assign v_7255 = v_7256 | v_7261;
  assign v_7256 = v_7257 | v_7259;
  assign v_7257 = mux_7257(v_7258);
  assign v_7258 = v_7248 & 1'h1;
  assign v_7259 = mux_7259(v_7260);
  assign v_7260 = ~v_7258;
  assign v_7261 = ~v_7248;
  assign v_7262 = v_7263 | v_7264;
  assign v_7263 = mux_7263(v_7250);
  assign v_7264 = mux_7264(v_7252);
  assign v_7266 = v_7267 | v_7269;
  assign v_7267 = act_7268 & 1'h1;
  assign act_7268 = v_974 | v_968;
  assign v_7269 = v_7270 & 1'h1;
  assign v_7270 = v_7271 & v_7272;
  assign v_7271 = ~act_7268;
  assign v_7272 = v_7273 | v_7277;
  assign v_7273 = v_7274 | v_7275;
  assign v_7274 = mux_7274(v_7245);
  assign v_7275 = mux_7275(v_7276);
  assign v_7276 = ~v_7245;
  assign v_7277 = ~v_7265;
  assign v_7278 = v_7279 | v_7280;
  assign v_7279 = mux_7279(v_7267);
  assign v_7280 = mux_7280(v_7269);
  assign v_7281 = v_7282 & 1'h1;
  assign v_7282 = v_7283 & v_7284;
  assign v_7283 = ~act_7244;
  assign v_7284 = v_7285 | v_7290;
  assign v_7285 = v_7286 | v_7288;
  assign v_7286 = mux_7286(v_7287);
  assign v_7287 = v_7241 & 1'h1;
  assign v_7288 = mux_7288(v_7289);
  assign v_7289 = ~v_7287;
  assign v_7290 = ~v_7241;
  assign v_7291 = v_7292 | v_7293;
  assign v_7292 = mux_7292(v_7243);
  assign v_7293 = mux_7293(v_7281);
  assign v_7295 = v_7296 | v_7334;
  assign v_7296 = act_7297 & 1'h1;
  assign act_7297 = v_7298 | v_7311;
  assign v_7298 = v_7299 & 1'h1;
  assign v_7299 = v_7300 & v_7318;
  assign v_7300 = ~v_7301;
  assign v_7302 = v_7303 | v_7305;
  assign v_7303 = act_7304 & 1'h1;
  assign act_7304 = v_988 | v_982;
  assign v_7305 = v_7306 & 1'h1;
  assign v_7306 = v_7307 & v_7308;
  assign v_7307 = ~act_7304;
  assign v_7308 = v_7309 | v_7314;
  assign v_7309 = v_7310 | v_7312;
  assign v_7310 = mux_7310(v_7311);
  assign v_7311 = v_7301 & 1'h1;
  assign v_7312 = mux_7312(v_7313);
  assign v_7313 = ~v_7311;
  assign v_7314 = ~v_7301;
  assign v_7315 = v_7316 | v_7317;
  assign v_7316 = mux_7316(v_7303);
  assign v_7317 = mux_7317(v_7305);
  assign v_7319 = v_7320 | v_7322;
  assign v_7320 = act_7321 & 1'h1;
  assign act_7321 = v_1002 | v_996;
  assign v_7322 = v_7323 & 1'h1;
  assign v_7323 = v_7324 & v_7325;
  assign v_7324 = ~act_7321;
  assign v_7325 = v_7326 | v_7330;
  assign v_7326 = v_7327 | v_7328;
  assign v_7327 = mux_7327(v_7298);
  assign v_7328 = mux_7328(v_7329);
  assign v_7329 = ~v_7298;
  assign v_7330 = ~v_7318;
  assign v_7331 = v_7332 | v_7333;
  assign v_7332 = mux_7332(v_7320);
  assign v_7333 = mux_7333(v_7322);
  assign v_7334 = v_7335 & 1'h1;
  assign v_7335 = v_7336 & v_7337;
  assign v_7336 = ~act_7297;
  assign v_7337 = v_7338 | v_7342;
  assign v_7338 = v_7339 | v_7340;
  assign v_7339 = mux_7339(v_7238);
  assign v_7340 = mux_7340(v_7341);
  assign v_7341 = ~v_7238;
  assign v_7342 = ~v_7294;
  assign v_7343 = v_7344 | v_7345;
  assign v_7344 = mux_7344(v_7296);
  assign v_7345 = mux_7345(v_7334);
  assign v_7346 = v_7347 & 1'h1;
  assign v_7347 = v_7348 & v_7349;
  assign v_7348 = ~act_7237;
  assign v_7349 = v_7350 | v_7354;
  assign v_7350 = v_7351 | v_7352;
  assign v_7351 = mux_7351(v_7106);
  assign v_7352 = mux_7352(v_7353);
  assign v_7353 = ~v_7106;
  assign v_7354 = ~v_7234;
  assign v_7355 = v_7356 | v_7357;
  assign v_7356 = mux_7356(v_7236);
  assign v_7357 = mux_7357(v_7346);
  assign v_7358 = v_7359 & 1'h1;
  assign v_7359 = v_7360 & v_7361;
  assign v_7360 = ~act_7105;
  assign v_7361 = v_7362 | v_7367;
  assign v_7362 = v_7363 | v_7365;
  assign v_7363 = mux_7363(v_7364);
  assign v_7364 = v_7102 & 1'h1;
  assign v_7365 = mux_7365(v_7366);
  assign v_7366 = ~v_7364;
  assign v_7367 = ~v_7102;
  assign v_7368 = v_7369 | v_7370;
  assign v_7369 = mux_7369(v_7104);
  assign v_7370 = mux_7370(v_7358);
  assign v_7372 = v_7373 | v_7627;
  assign v_7373 = act_7374 & 1'h1;
  assign act_7374 = v_7375 | v_7496;
  assign v_7375 = v_7376 & 1'h1;
  assign v_7376 = v_7377 & v_7503;
  assign v_7377 = ~v_7378;
  assign v_7379 = v_7380 | v_7490;
  assign v_7380 = act_7381 & 1'h1;
  assign act_7381 = v_7382 | v_7431;
  assign v_7382 = v_7383 & 1'h1;
  assign v_7383 = v_7384 & v_7438;
  assign v_7384 = ~v_7385;
  assign v_7386 = v_7387 | v_7425;
  assign v_7387 = act_7388 & 1'h1;
  assign act_7388 = v_7389 | v_7402;
  assign v_7389 = v_7390 & 1'h1;
  assign v_7390 = v_7391 & v_7409;
  assign v_7391 = ~v_7392;
  assign v_7393 = v_7394 | v_7396;
  assign v_7394 = act_7395 & 1'h1;
  assign act_7395 = v_1016 | v_1010;
  assign v_7396 = v_7397 & 1'h1;
  assign v_7397 = v_7398 & v_7399;
  assign v_7398 = ~act_7395;
  assign v_7399 = v_7400 | v_7405;
  assign v_7400 = v_7401 | v_7403;
  assign v_7401 = mux_7401(v_7402);
  assign v_7402 = v_7392 & 1'h1;
  assign v_7403 = mux_7403(v_7404);
  assign v_7404 = ~v_7402;
  assign v_7405 = ~v_7392;
  assign v_7406 = v_7407 | v_7408;
  assign v_7407 = mux_7407(v_7394);
  assign v_7408 = mux_7408(v_7396);
  assign v_7410 = v_7411 | v_7413;
  assign v_7411 = act_7412 & 1'h1;
  assign act_7412 = v_1030 | v_1024;
  assign v_7413 = v_7414 & 1'h1;
  assign v_7414 = v_7415 & v_7416;
  assign v_7415 = ~act_7412;
  assign v_7416 = v_7417 | v_7421;
  assign v_7417 = v_7418 | v_7419;
  assign v_7418 = mux_7418(v_7389);
  assign v_7419 = mux_7419(v_7420);
  assign v_7420 = ~v_7389;
  assign v_7421 = ~v_7409;
  assign v_7422 = v_7423 | v_7424;
  assign v_7423 = mux_7423(v_7411);
  assign v_7424 = mux_7424(v_7413);
  assign v_7425 = v_7426 & 1'h1;
  assign v_7426 = v_7427 & v_7428;
  assign v_7427 = ~act_7388;
  assign v_7428 = v_7429 | v_7434;
  assign v_7429 = v_7430 | v_7432;
  assign v_7430 = mux_7430(v_7431);
  assign v_7431 = v_7385 & 1'h1;
  assign v_7432 = mux_7432(v_7433);
  assign v_7433 = ~v_7431;
  assign v_7434 = ~v_7385;
  assign v_7435 = v_7436 | v_7437;
  assign v_7436 = mux_7436(v_7387);
  assign v_7437 = mux_7437(v_7425);
  assign v_7439 = v_7440 | v_7478;
  assign v_7440 = act_7441 & 1'h1;
  assign act_7441 = v_7442 | v_7455;
  assign v_7442 = v_7443 & 1'h1;
  assign v_7443 = v_7444 & v_7462;
  assign v_7444 = ~v_7445;
  assign v_7446 = v_7447 | v_7449;
  assign v_7447 = act_7448 & 1'h1;
  assign act_7448 = v_1044 | v_1038;
  assign v_7449 = v_7450 & 1'h1;
  assign v_7450 = v_7451 & v_7452;
  assign v_7451 = ~act_7448;
  assign v_7452 = v_7453 | v_7458;
  assign v_7453 = v_7454 | v_7456;
  assign v_7454 = mux_7454(v_7455);
  assign v_7455 = v_7445 & 1'h1;
  assign v_7456 = mux_7456(v_7457);
  assign v_7457 = ~v_7455;
  assign v_7458 = ~v_7445;
  assign v_7459 = v_7460 | v_7461;
  assign v_7460 = mux_7460(v_7447);
  assign v_7461 = mux_7461(v_7449);
  assign v_7463 = v_7464 | v_7466;
  assign v_7464 = act_7465 & 1'h1;
  assign act_7465 = v_1058 | v_1052;
  assign v_7466 = v_7467 & 1'h1;
  assign v_7467 = v_7468 & v_7469;
  assign v_7468 = ~act_7465;
  assign v_7469 = v_7470 | v_7474;
  assign v_7470 = v_7471 | v_7472;
  assign v_7471 = mux_7471(v_7442);
  assign v_7472 = mux_7472(v_7473);
  assign v_7473 = ~v_7442;
  assign v_7474 = ~v_7462;
  assign v_7475 = v_7476 | v_7477;
  assign v_7476 = mux_7476(v_7464);
  assign v_7477 = mux_7477(v_7466);
  assign v_7478 = v_7479 & 1'h1;
  assign v_7479 = v_7480 & v_7481;
  assign v_7480 = ~act_7441;
  assign v_7481 = v_7482 | v_7486;
  assign v_7482 = v_7483 | v_7484;
  assign v_7483 = mux_7483(v_7382);
  assign v_7484 = mux_7484(v_7485);
  assign v_7485 = ~v_7382;
  assign v_7486 = ~v_7438;
  assign v_7487 = v_7488 | v_7489;
  assign v_7488 = mux_7488(v_7440);
  assign v_7489 = mux_7489(v_7478);
  assign v_7490 = v_7491 & 1'h1;
  assign v_7491 = v_7492 & v_7493;
  assign v_7492 = ~act_7381;
  assign v_7493 = v_7494 | v_7499;
  assign v_7494 = v_7495 | v_7497;
  assign v_7495 = mux_7495(v_7496);
  assign v_7496 = v_7378 & 1'h1;
  assign v_7497 = mux_7497(v_7498);
  assign v_7498 = ~v_7496;
  assign v_7499 = ~v_7378;
  assign v_7500 = v_7501 | v_7502;
  assign v_7501 = mux_7501(v_7380);
  assign v_7502 = mux_7502(v_7490);
  assign v_7504 = v_7505 | v_7615;
  assign v_7505 = act_7506 & 1'h1;
  assign act_7506 = v_7507 | v_7556;
  assign v_7507 = v_7508 & 1'h1;
  assign v_7508 = v_7509 & v_7563;
  assign v_7509 = ~v_7510;
  assign v_7511 = v_7512 | v_7550;
  assign v_7512 = act_7513 & 1'h1;
  assign act_7513 = v_7514 | v_7527;
  assign v_7514 = v_7515 & 1'h1;
  assign v_7515 = v_7516 & v_7534;
  assign v_7516 = ~v_7517;
  assign v_7518 = v_7519 | v_7521;
  assign v_7519 = act_7520 & 1'h1;
  assign act_7520 = v_1072 | v_1066;
  assign v_7521 = v_7522 & 1'h1;
  assign v_7522 = v_7523 & v_7524;
  assign v_7523 = ~act_7520;
  assign v_7524 = v_7525 | v_7530;
  assign v_7525 = v_7526 | v_7528;
  assign v_7526 = mux_7526(v_7527);
  assign v_7527 = v_7517 & 1'h1;
  assign v_7528 = mux_7528(v_7529);
  assign v_7529 = ~v_7527;
  assign v_7530 = ~v_7517;
  assign v_7531 = v_7532 | v_7533;
  assign v_7532 = mux_7532(v_7519);
  assign v_7533 = mux_7533(v_7521);
  assign v_7535 = v_7536 | v_7538;
  assign v_7536 = act_7537 & 1'h1;
  assign act_7537 = v_1086 | v_1080;
  assign v_7538 = v_7539 & 1'h1;
  assign v_7539 = v_7540 & v_7541;
  assign v_7540 = ~act_7537;
  assign v_7541 = v_7542 | v_7546;
  assign v_7542 = v_7543 | v_7544;
  assign v_7543 = mux_7543(v_7514);
  assign v_7544 = mux_7544(v_7545);
  assign v_7545 = ~v_7514;
  assign v_7546 = ~v_7534;
  assign v_7547 = v_7548 | v_7549;
  assign v_7548 = mux_7548(v_7536);
  assign v_7549 = mux_7549(v_7538);
  assign v_7550 = v_7551 & 1'h1;
  assign v_7551 = v_7552 & v_7553;
  assign v_7552 = ~act_7513;
  assign v_7553 = v_7554 | v_7559;
  assign v_7554 = v_7555 | v_7557;
  assign v_7555 = mux_7555(v_7556);
  assign v_7556 = v_7510 & 1'h1;
  assign v_7557 = mux_7557(v_7558);
  assign v_7558 = ~v_7556;
  assign v_7559 = ~v_7510;
  assign v_7560 = v_7561 | v_7562;
  assign v_7561 = mux_7561(v_7512);
  assign v_7562 = mux_7562(v_7550);
  assign v_7564 = v_7565 | v_7603;
  assign v_7565 = act_7566 & 1'h1;
  assign act_7566 = v_7567 | v_7580;
  assign v_7567 = v_7568 & 1'h1;
  assign v_7568 = v_7569 & v_7587;
  assign v_7569 = ~v_7570;
  assign v_7571 = v_7572 | v_7574;
  assign v_7572 = act_7573 & 1'h1;
  assign act_7573 = v_1100 | v_1094;
  assign v_7574 = v_7575 & 1'h1;
  assign v_7575 = v_7576 & v_7577;
  assign v_7576 = ~act_7573;
  assign v_7577 = v_7578 | v_7583;
  assign v_7578 = v_7579 | v_7581;
  assign v_7579 = mux_7579(v_7580);
  assign v_7580 = v_7570 & 1'h1;
  assign v_7581 = mux_7581(v_7582);
  assign v_7582 = ~v_7580;
  assign v_7583 = ~v_7570;
  assign v_7584 = v_7585 | v_7586;
  assign v_7585 = mux_7585(v_7572);
  assign v_7586 = mux_7586(v_7574);
  assign v_7588 = v_7589 | v_7591;
  assign v_7589 = act_7590 & 1'h1;
  assign act_7590 = v_1114 | v_1108;
  assign v_7591 = v_7592 & 1'h1;
  assign v_7592 = v_7593 & v_7594;
  assign v_7593 = ~act_7590;
  assign v_7594 = v_7595 | v_7599;
  assign v_7595 = v_7596 | v_7597;
  assign v_7596 = mux_7596(v_7567);
  assign v_7597 = mux_7597(v_7598);
  assign v_7598 = ~v_7567;
  assign v_7599 = ~v_7587;
  assign v_7600 = v_7601 | v_7602;
  assign v_7601 = mux_7601(v_7589);
  assign v_7602 = mux_7602(v_7591);
  assign v_7603 = v_7604 & 1'h1;
  assign v_7604 = v_7605 & v_7606;
  assign v_7605 = ~act_7566;
  assign v_7606 = v_7607 | v_7611;
  assign v_7607 = v_7608 | v_7609;
  assign v_7608 = mux_7608(v_7507);
  assign v_7609 = mux_7609(v_7610);
  assign v_7610 = ~v_7507;
  assign v_7611 = ~v_7563;
  assign v_7612 = v_7613 | v_7614;
  assign v_7613 = mux_7613(v_7565);
  assign v_7614 = mux_7614(v_7603);
  assign v_7615 = v_7616 & 1'h1;
  assign v_7616 = v_7617 & v_7618;
  assign v_7617 = ~act_7506;
  assign v_7618 = v_7619 | v_7623;
  assign v_7619 = v_7620 | v_7621;
  assign v_7620 = mux_7620(v_7375);
  assign v_7621 = mux_7621(v_7622);
  assign v_7622 = ~v_7375;
  assign v_7623 = ~v_7503;
  assign v_7624 = v_7625 | v_7626;
  assign v_7625 = mux_7625(v_7505);
  assign v_7626 = mux_7626(v_7615);
  assign v_7627 = v_7628 & 1'h1;
  assign v_7628 = v_7629 & v_7630;
  assign v_7629 = ~act_7374;
  assign v_7630 = v_7631 | v_7635;
  assign v_7631 = v_7632 | v_7633;
  assign v_7632 = mux_7632(v_7099);
  assign v_7633 = mux_7633(v_7634);
  assign v_7634 = ~v_7099;
  assign v_7635 = ~v_7371;
  assign v_7636 = v_7637 | v_7638;
  assign v_7637 = mux_7637(v_7373);
  assign v_7638 = mux_7638(v_7627);
  assign v_7639 = v_7640 & 1'h1;
  assign v_7640 = v_7641 & v_7642;
  assign v_7641 = ~act_7098;
  assign v_7642 = v_7643 | v_7647;
  assign v_7643 = v_7644 | v_7645;
  assign v_7644 = mux_7644(v_6535);
  assign v_7645 = mux_7645(v_7646);
  assign v_7646 = ~v_6535;
  assign v_7647 = ~v_7095;
  assign v_7648 = v_7649 | v_7650;
  assign v_7649 = mux_7649(v_7097);
  assign v_7650 = mux_7650(v_7639);
  assign v_7651 = v_7652 & 1'h1;
  assign v_7652 = v_7653 & v_7654;
  assign v_7653 = ~act_6534;
  assign v_7654 = v_7655 | v_7659;
  assign v_7655 = v_7656 | v_7657;
  assign v_7656 = mux_7656(v_5395);
  assign v_7657 = mux_7657(v_7658);
  assign v_7658 = ~v_5395;
  assign v_7659 = ~v_6531;
  assign v_7660 = v_7661 | v_7662;
  assign v_7661 = mux_7661(v_6533);
  assign v_7662 = mux_7662(v_7651);
  assign v_7663 = v_7664 & 1'h1;
  assign v_7664 = v_7665 & v_7666;
  assign v_7665 = ~act_5394;
  assign v_7666 = v_7667 | v_7672;
  assign v_7667 = v_7668 | v_7670;
  assign v_7668 = mux_7668(v_7669);
  assign v_7669 = v_5391 & 1'h1;
  assign v_7670 = mux_7670(v_7671);
  assign v_7671 = ~v_7669;
  assign v_7672 = ~v_5391;
  assign v_7673 = v_7674 | v_7675;
  assign v_7674 = mux_7674(v_5393);
  assign v_7675 = mux_7675(v_7663);
  assign v_7677 = v_7678 | v_9948;
  assign v_7678 = act_7679 & 1'h1;
  assign act_7679 = v_7680 | v_8809;
  assign v_7680 = v_7681 & 1'h1;
  assign v_7681 = v_7682 & v_8816;
  assign v_7682 = ~v_7683;
  assign v_7684 = v_7685 | v_8803;
  assign v_7685 = act_7686 & 1'h1;
  assign act_7686 = v_7687 | v_8240;
  assign v_7687 = v_7688 & 1'h1;
  assign v_7688 = v_7689 & v_8247;
  assign v_7689 = ~v_7690;
  assign v_7691 = v_7692 | v_8234;
  assign v_7692 = act_7693 & 1'h1;
  assign act_7693 = v_7694 | v_7959;
  assign v_7694 = v_7695 & 1'h1;
  assign v_7695 = v_7696 & v_7966;
  assign v_7696 = ~v_7697;
  assign v_7698 = v_7699 | v_7953;
  assign v_7699 = act_7700 & 1'h1;
  assign act_7700 = v_7701 | v_7822;
  assign v_7701 = v_7702 & 1'h1;
  assign v_7702 = v_7703 & v_7829;
  assign v_7703 = ~v_7704;
  assign v_7705 = v_7706 | v_7816;
  assign v_7706 = act_7707 & 1'h1;
  assign act_7707 = v_7708 | v_7757;
  assign v_7708 = v_7709 & 1'h1;
  assign v_7709 = v_7710 & v_7764;
  assign v_7710 = ~v_7711;
  assign v_7712 = v_7713 | v_7751;
  assign v_7713 = act_7714 & 1'h1;
  assign act_7714 = v_7715 | v_7728;
  assign v_7715 = v_7716 & 1'h1;
  assign v_7716 = v_7717 & v_7735;
  assign v_7717 = ~v_7718;
  assign v_7719 = v_7720 | v_7722;
  assign v_7720 = act_7721 & 1'h1;
  assign act_7721 = v_1128 | v_1122;
  assign v_7722 = v_7723 & 1'h1;
  assign v_7723 = v_7724 & v_7725;
  assign v_7724 = ~act_7721;
  assign v_7725 = v_7726 | v_7731;
  assign v_7726 = v_7727 | v_7729;
  assign v_7727 = mux_7727(v_7728);
  assign v_7728 = v_7718 & 1'h1;
  assign v_7729 = mux_7729(v_7730);
  assign v_7730 = ~v_7728;
  assign v_7731 = ~v_7718;
  assign v_7732 = v_7733 | v_7734;
  assign v_7733 = mux_7733(v_7720);
  assign v_7734 = mux_7734(v_7722);
  assign v_7736 = v_7737 | v_7739;
  assign v_7737 = act_7738 & 1'h1;
  assign act_7738 = v_1142 | v_1136;
  assign v_7739 = v_7740 & 1'h1;
  assign v_7740 = v_7741 & v_7742;
  assign v_7741 = ~act_7738;
  assign v_7742 = v_7743 | v_7747;
  assign v_7743 = v_7744 | v_7745;
  assign v_7744 = mux_7744(v_7715);
  assign v_7745 = mux_7745(v_7746);
  assign v_7746 = ~v_7715;
  assign v_7747 = ~v_7735;
  assign v_7748 = v_7749 | v_7750;
  assign v_7749 = mux_7749(v_7737);
  assign v_7750 = mux_7750(v_7739);
  assign v_7751 = v_7752 & 1'h1;
  assign v_7752 = v_7753 & v_7754;
  assign v_7753 = ~act_7714;
  assign v_7754 = v_7755 | v_7760;
  assign v_7755 = v_7756 | v_7758;
  assign v_7756 = mux_7756(v_7757);
  assign v_7757 = v_7711 & 1'h1;
  assign v_7758 = mux_7758(v_7759);
  assign v_7759 = ~v_7757;
  assign v_7760 = ~v_7711;
  assign v_7761 = v_7762 | v_7763;
  assign v_7762 = mux_7762(v_7713);
  assign v_7763 = mux_7763(v_7751);
  assign v_7765 = v_7766 | v_7804;
  assign v_7766 = act_7767 & 1'h1;
  assign act_7767 = v_7768 | v_7781;
  assign v_7768 = v_7769 & 1'h1;
  assign v_7769 = v_7770 & v_7788;
  assign v_7770 = ~v_7771;
  assign v_7772 = v_7773 | v_7775;
  assign v_7773 = act_7774 & 1'h1;
  assign act_7774 = v_1156 | v_1150;
  assign v_7775 = v_7776 & 1'h1;
  assign v_7776 = v_7777 & v_7778;
  assign v_7777 = ~act_7774;
  assign v_7778 = v_7779 | v_7784;
  assign v_7779 = v_7780 | v_7782;
  assign v_7780 = mux_7780(v_7781);
  assign v_7781 = v_7771 & 1'h1;
  assign v_7782 = mux_7782(v_7783);
  assign v_7783 = ~v_7781;
  assign v_7784 = ~v_7771;
  assign v_7785 = v_7786 | v_7787;
  assign v_7786 = mux_7786(v_7773);
  assign v_7787 = mux_7787(v_7775);
  assign v_7789 = v_7790 | v_7792;
  assign v_7790 = act_7791 & 1'h1;
  assign act_7791 = v_1170 | v_1164;
  assign v_7792 = v_7793 & 1'h1;
  assign v_7793 = v_7794 & v_7795;
  assign v_7794 = ~act_7791;
  assign v_7795 = v_7796 | v_7800;
  assign v_7796 = v_7797 | v_7798;
  assign v_7797 = mux_7797(v_7768);
  assign v_7798 = mux_7798(v_7799);
  assign v_7799 = ~v_7768;
  assign v_7800 = ~v_7788;
  assign v_7801 = v_7802 | v_7803;
  assign v_7802 = mux_7802(v_7790);
  assign v_7803 = mux_7803(v_7792);
  assign v_7804 = v_7805 & 1'h1;
  assign v_7805 = v_7806 & v_7807;
  assign v_7806 = ~act_7767;
  assign v_7807 = v_7808 | v_7812;
  assign v_7808 = v_7809 | v_7810;
  assign v_7809 = mux_7809(v_7708);
  assign v_7810 = mux_7810(v_7811);
  assign v_7811 = ~v_7708;
  assign v_7812 = ~v_7764;
  assign v_7813 = v_7814 | v_7815;
  assign v_7814 = mux_7814(v_7766);
  assign v_7815 = mux_7815(v_7804);
  assign v_7816 = v_7817 & 1'h1;
  assign v_7817 = v_7818 & v_7819;
  assign v_7818 = ~act_7707;
  assign v_7819 = v_7820 | v_7825;
  assign v_7820 = v_7821 | v_7823;
  assign v_7821 = mux_7821(v_7822);
  assign v_7822 = v_7704 & 1'h1;
  assign v_7823 = mux_7823(v_7824);
  assign v_7824 = ~v_7822;
  assign v_7825 = ~v_7704;
  assign v_7826 = v_7827 | v_7828;
  assign v_7827 = mux_7827(v_7706);
  assign v_7828 = mux_7828(v_7816);
  assign v_7830 = v_7831 | v_7941;
  assign v_7831 = act_7832 & 1'h1;
  assign act_7832 = v_7833 | v_7882;
  assign v_7833 = v_7834 & 1'h1;
  assign v_7834 = v_7835 & v_7889;
  assign v_7835 = ~v_7836;
  assign v_7837 = v_7838 | v_7876;
  assign v_7838 = act_7839 & 1'h1;
  assign act_7839 = v_7840 | v_7853;
  assign v_7840 = v_7841 & 1'h1;
  assign v_7841 = v_7842 & v_7860;
  assign v_7842 = ~v_7843;
  assign v_7844 = v_7845 | v_7847;
  assign v_7845 = act_7846 & 1'h1;
  assign act_7846 = v_1184 | v_1178;
  assign v_7847 = v_7848 & 1'h1;
  assign v_7848 = v_7849 & v_7850;
  assign v_7849 = ~act_7846;
  assign v_7850 = v_7851 | v_7856;
  assign v_7851 = v_7852 | v_7854;
  assign v_7852 = mux_7852(v_7853);
  assign v_7853 = v_7843 & 1'h1;
  assign v_7854 = mux_7854(v_7855);
  assign v_7855 = ~v_7853;
  assign v_7856 = ~v_7843;
  assign v_7857 = v_7858 | v_7859;
  assign v_7858 = mux_7858(v_7845);
  assign v_7859 = mux_7859(v_7847);
  assign v_7861 = v_7862 | v_7864;
  assign v_7862 = act_7863 & 1'h1;
  assign act_7863 = v_1198 | v_1192;
  assign v_7864 = v_7865 & 1'h1;
  assign v_7865 = v_7866 & v_7867;
  assign v_7866 = ~act_7863;
  assign v_7867 = v_7868 | v_7872;
  assign v_7868 = v_7869 | v_7870;
  assign v_7869 = mux_7869(v_7840);
  assign v_7870 = mux_7870(v_7871);
  assign v_7871 = ~v_7840;
  assign v_7872 = ~v_7860;
  assign v_7873 = v_7874 | v_7875;
  assign v_7874 = mux_7874(v_7862);
  assign v_7875 = mux_7875(v_7864);
  assign v_7876 = v_7877 & 1'h1;
  assign v_7877 = v_7878 & v_7879;
  assign v_7878 = ~act_7839;
  assign v_7879 = v_7880 | v_7885;
  assign v_7880 = v_7881 | v_7883;
  assign v_7881 = mux_7881(v_7882);
  assign v_7882 = v_7836 & 1'h1;
  assign v_7883 = mux_7883(v_7884);
  assign v_7884 = ~v_7882;
  assign v_7885 = ~v_7836;
  assign v_7886 = v_7887 | v_7888;
  assign v_7887 = mux_7887(v_7838);
  assign v_7888 = mux_7888(v_7876);
  assign v_7890 = v_7891 | v_7929;
  assign v_7891 = act_7892 & 1'h1;
  assign act_7892 = v_7893 | v_7906;
  assign v_7893 = v_7894 & 1'h1;
  assign v_7894 = v_7895 & v_7913;
  assign v_7895 = ~v_7896;
  assign v_7897 = v_7898 | v_7900;
  assign v_7898 = act_7899 & 1'h1;
  assign act_7899 = v_1212 | v_1206;
  assign v_7900 = v_7901 & 1'h1;
  assign v_7901 = v_7902 & v_7903;
  assign v_7902 = ~act_7899;
  assign v_7903 = v_7904 | v_7909;
  assign v_7904 = v_7905 | v_7907;
  assign v_7905 = mux_7905(v_7906);
  assign v_7906 = v_7896 & 1'h1;
  assign v_7907 = mux_7907(v_7908);
  assign v_7908 = ~v_7906;
  assign v_7909 = ~v_7896;
  assign v_7910 = v_7911 | v_7912;
  assign v_7911 = mux_7911(v_7898);
  assign v_7912 = mux_7912(v_7900);
  assign v_7914 = v_7915 | v_7917;
  assign v_7915 = act_7916 & 1'h1;
  assign act_7916 = v_1226 | v_1220;
  assign v_7917 = v_7918 & 1'h1;
  assign v_7918 = v_7919 & v_7920;
  assign v_7919 = ~act_7916;
  assign v_7920 = v_7921 | v_7925;
  assign v_7921 = v_7922 | v_7923;
  assign v_7922 = mux_7922(v_7893);
  assign v_7923 = mux_7923(v_7924);
  assign v_7924 = ~v_7893;
  assign v_7925 = ~v_7913;
  assign v_7926 = v_7927 | v_7928;
  assign v_7927 = mux_7927(v_7915);
  assign v_7928 = mux_7928(v_7917);
  assign v_7929 = v_7930 & 1'h1;
  assign v_7930 = v_7931 & v_7932;
  assign v_7931 = ~act_7892;
  assign v_7932 = v_7933 | v_7937;
  assign v_7933 = v_7934 | v_7935;
  assign v_7934 = mux_7934(v_7833);
  assign v_7935 = mux_7935(v_7936);
  assign v_7936 = ~v_7833;
  assign v_7937 = ~v_7889;
  assign v_7938 = v_7939 | v_7940;
  assign v_7939 = mux_7939(v_7891);
  assign v_7940 = mux_7940(v_7929);
  assign v_7941 = v_7942 & 1'h1;
  assign v_7942 = v_7943 & v_7944;
  assign v_7943 = ~act_7832;
  assign v_7944 = v_7945 | v_7949;
  assign v_7945 = v_7946 | v_7947;
  assign v_7946 = mux_7946(v_7701);
  assign v_7947 = mux_7947(v_7948);
  assign v_7948 = ~v_7701;
  assign v_7949 = ~v_7829;
  assign v_7950 = v_7951 | v_7952;
  assign v_7951 = mux_7951(v_7831);
  assign v_7952 = mux_7952(v_7941);
  assign v_7953 = v_7954 & 1'h1;
  assign v_7954 = v_7955 & v_7956;
  assign v_7955 = ~act_7700;
  assign v_7956 = v_7957 | v_7962;
  assign v_7957 = v_7958 | v_7960;
  assign v_7958 = mux_7958(v_7959);
  assign v_7959 = v_7697 & 1'h1;
  assign v_7960 = mux_7960(v_7961);
  assign v_7961 = ~v_7959;
  assign v_7962 = ~v_7697;
  assign v_7963 = v_7964 | v_7965;
  assign v_7964 = mux_7964(v_7699);
  assign v_7965 = mux_7965(v_7953);
  assign v_7967 = v_7968 | v_8222;
  assign v_7968 = act_7969 & 1'h1;
  assign act_7969 = v_7970 | v_8091;
  assign v_7970 = v_7971 & 1'h1;
  assign v_7971 = v_7972 & v_8098;
  assign v_7972 = ~v_7973;
  assign v_7974 = v_7975 | v_8085;
  assign v_7975 = act_7976 & 1'h1;
  assign act_7976 = v_7977 | v_8026;
  assign v_7977 = v_7978 & 1'h1;
  assign v_7978 = v_7979 & v_8033;
  assign v_7979 = ~v_7980;
  assign v_7981 = v_7982 | v_8020;
  assign v_7982 = act_7983 & 1'h1;
  assign act_7983 = v_7984 | v_7997;
  assign v_7984 = v_7985 & 1'h1;
  assign v_7985 = v_7986 & v_8004;
  assign v_7986 = ~v_7987;
  assign v_7988 = v_7989 | v_7991;
  assign v_7989 = act_7990 & 1'h1;
  assign act_7990 = v_1240 | v_1234;
  assign v_7991 = v_7992 & 1'h1;
  assign v_7992 = v_7993 & v_7994;
  assign v_7993 = ~act_7990;
  assign v_7994 = v_7995 | v_8000;
  assign v_7995 = v_7996 | v_7998;
  assign v_7996 = mux_7996(v_7997);
  assign v_7997 = v_7987 & 1'h1;
  assign v_7998 = mux_7998(v_7999);
  assign v_7999 = ~v_7997;
  assign v_8000 = ~v_7987;
  assign v_8001 = v_8002 | v_8003;
  assign v_8002 = mux_8002(v_7989);
  assign v_8003 = mux_8003(v_7991);
  assign v_8005 = v_8006 | v_8008;
  assign v_8006 = act_8007 & 1'h1;
  assign act_8007 = v_1254 | v_1248;
  assign v_8008 = v_8009 & 1'h1;
  assign v_8009 = v_8010 & v_8011;
  assign v_8010 = ~act_8007;
  assign v_8011 = v_8012 | v_8016;
  assign v_8012 = v_8013 | v_8014;
  assign v_8013 = mux_8013(v_7984);
  assign v_8014 = mux_8014(v_8015);
  assign v_8015 = ~v_7984;
  assign v_8016 = ~v_8004;
  assign v_8017 = v_8018 | v_8019;
  assign v_8018 = mux_8018(v_8006);
  assign v_8019 = mux_8019(v_8008);
  assign v_8020 = v_8021 & 1'h1;
  assign v_8021 = v_8022 & v_8023;
  assign v_8022 = ~act_7983;
  assign v_8023 = v_8024 | v_8029;
  assign v_8024 = v_8025 | v_8027;
  assign v_8025 = mux_8025(v_8026);
  assign v_8026 = v_7980 & 1'h1;
  assign v_8027 = mux_8027(v_8028);
  assign v_8028 = ~v_8026;
  assign v_8029 = ~v_7980;
  assign v_8030 = v_8031 | v_8032;
  assign v_8031 = mux_8031(v_7982);
  assign v_8032 = mux_8032(v_8020);
  assign v_8034 = v_8035 | v_8073;
  assign v_8035 = act_8036 & 1'h1;
  assign act_8036 = v_8037 | v_8050;
  assign v_8037 = v_8038 & 1'h1;
  assign v_8038 = v_8039 & v_8057;
  assign v_8039 = ~v_8040;
  assign v_8041 = v_8042 | v_8044;
  assign v_8042 = act_8043 & 1'h1;
  assign act_8043 = v_1268 | v_1262;
  assign v_8044 = v_8045 & 1'h1;
  assign v_8045 = v_8046 & v_8047;
  assign v_8046 = ~act_8043;
  assign v_8047 = v_8048 | v_8053;
  assign v_8048 = v_8049 | v_8051;
  assign v_8049 = mux_8049(v_8050);
  assign v_8050 = v_8040 & 1'h1;
  assign v_8051 = mux_8051(v_8052);
  assign v_8052 = ~v_8050;
  assign v_8053 = ~v_8040;
  assign v_8054 = v_8055 | v_8056;
  assign v_8055 = mux_8055(v_8042);
  assign v_8056 = mux_8056(v_8044);
  assign v_8058 = v_8059 | v_8061;
  assign v_8059 = act_8060 & 1'h1;
  assign act_8060 = v_1282 | v_1276;
  assign v_8061 = v_8062 & 1'h1;
  assign v_8062 = v_8063 & v_8064;
  assign v_8063 = ~act_8060;
  assign v_8064 = v_8065 | v_8069;
  assign v_8065 = v_8066 | v_8067;
  assign v_8066 = mux_8066(v_8037);
  assign v_8067 = mux_8067(v_8068);
  assign v_8068 = ~v_8037;
  assign v_8069 = ~v_8057;
  assign v_8070 = v_8071 | v_8072;
  assign v_8071 = mux_8071(v_8059);
  assign v_8072 = mux_8072(v_8061);
  assign v_8073 = v_8074 & 1'h1;
  assign v_8074 = v_8075 & v_8076;
  assign v_8075 = ~act_8036;
  assign v_8076 = v_8077 | v_8081;
  assign v_8077 = v_8078 | v_8079;
  assign v_8078 = mux_8078(v_7977);
  assign v_8079 = mux_8079(v_8080);
  assign v_8080 = ~v_7977;
  assign v_8081 = ~v_8033;
  assign v_8082 = v_8083 | v_8084;
  assign v_8083 = mux_8083(v_8035);
  assign v_8084 = mux_8084(v_8073);
  assign v_8085 = v_8086 & 1'h1;
  assign v_8086 = v_8087 & v_8088;
  assign v_8087 = ~act_7976;
  assign v_8088 = v_8089 | v_8094;
  assign v_8089 = v_8090 | v_8092;
  assign v_8090 = mux_8090(v_8091);
  assign v_8091 = v_7973 & 1'h1;
  assign v_8092 = mux_8092(v_8093);
  assign v_8093 = ~v_8091;
  assign v_8094 = ~v_7973;
  assign v_8095 = v_8096 | v_8097;
  assign v_8096 = mux_8096(v_7975);
  assign v_8097 = mux_8097(v_8085);
  assign v_8099 = v_8100 | v_8210;
  assign v_8100 = act_8101 & 1'h1;
  assign act_8101 = v_8102 | v_8151;
  assign v_8102 = v_8103 & 1'h1;
  assign v_8103 = v_8104 & v_8158;
  assign v_8104 = ~v_8105;
  assign v_8106 = v_8107 | v_8145;
  assign v_8107 = act_8108 & 1'h1;
  assign act_8108 = v_8109 | v_8122;
  assign v_8109 = v_8110 & 1'h1;
  assign v_8110 = v_8111 & v_8129;
  assign v_8111 = ~v_8112;
  assign v_8113 = v_8114 | v_8116;
  assign v_8114 = act_8115 & 1'h1;
  assign act_8115 = v_1296 | v_1290;
  assign v_8116 = v_8117 & 1'h1;
  assign v_8117 = v_8118 & v_8119;
  assign v_8118 = ~act_8115;
  assign v_8119 = v_8120 | v_8125;
  assign v_8120 = v_8121 | v_8123;
  assign v_8121 = mux_8121(v_8122);
  assign v_8122 = v_8112 & 1'h1;
  assign v_8123 = mux_8123(v_8124);
  assign v_8124 = ~v_8122;
  assign v_8125 = ~v_8112;
  assign v_8126 = v_8127 | v_8128;
  assign v_8127 = mux_8127(v_8114);
  assign v_8128 = mux_8128(v_8116);
  assign v_8130 = v_8131 | v_8133;
  assign v_8131 = act_8132 & 1'h1;
  assign act_8132 = v_1310 | v_1304;
  assign v_8133 = v_8134 & 1'h1;
  assign v_8134 = v_8135 & v_8136;
  assign v_8135 = ~act_8132;
  assign v_8136 = v_8137 | v_8141;
  assign v_8137 = v_8138 | v_8139;
  assign v_8138 = mux_8138(v_8109);
  assign v_8139 = mux_8139(v_8140);
  assign v_8140 = ~v_8109;
  assign v_8141 = ~v_8129;
  assign v_8142 = v_8143 | v_8144;
  assign v_8143 = mux_8143(v_8131);
  assign v_8144 = mux_8144(v_8133);
  assign v_8145 = v_8146 & 1'h1;
  assign v_8146 = v_8147 & v_8148;
  assign v_8147 = ~act_8108;
  assign v_8148 = v_8149 | v_8154;
  assign v_8149 = v_8150 | v_8152;
  assign v_8150 = mux_8150(v_8151);
  assign v_8151 = v_8105 & 1'h1;
  assign v_8152 = mux_8152(v_8153);
  assign v_8153 = ~v_8151;
  assign v_8154 = ~v_8105;
  assign v_8155 = v_8156 | v_8157;
  assign v_8156 = mux_8156(v_8107);
  assign v_8157 = mux_8157(v_8145);
  assign v_8159 = v_8160 | v_8198;
  assign v_8160 = act_8161 & 1'h1;
  assign act_8161 = v_8162 | v_8175;
  assign v_8162 = v_8163 & 1'h1;
  assign v_8163 = v_8164 & v_8182;
  assign v_8164 = ~v_8165;
  assign v_8166 = v_8167 | v_8169;
  assign v_8167 = act_8168 & 1'h1;
  assign act_8168 = v_1324 | v_1318;
  assign v_8169 = v_8170 & 1'h1;
  assign v_8170 = v_8171 & v_8172;
  assign v_8171 = ~act_8168;
  assign v_8172 = v_8173 | v_8178;
  assign v_8173 = v_8174 | v_8176;
  assign v_8174 = mux_8174(v_8175);
  assign v_8175 = v_8165 & 1'h1;
  assign v_8176 = mux_8176(v_8177);
  assign v_8177 = ~v_8175;
  assign v_8178 = ~v_8165;
  assign v_8179 = v_8180 | v_8181;
  assign v_8180 = mux_8180(v_8167);
  assign v_8181 = mux_8181(v_8169);
  assign v_8183 = v_8184 | v_8186;
  assign v_8184 = act_8185 & 1'h1;
  assign act_8185 = v_1338 | v_1332;
  assign v_8186 = v_8187 & 1'h1;
  assign v_8187 = v_8188 & v_8189;
  assign v_8188 = ~act_8185;
  assign v_8189 = v_8190 | v_8194;
  assign v_8190 = v_8191 | v_8192;
  assign v_8191 = mux_8191(v_8162);
  assign v_8192 = mux_8192(v_8193);
  assign v_8193 = ~v_8162;
  assign v_8194 = ~v_8182;
  assign v_8195 = v_8196 | v_8197;
  assign v_8196 = mux_8196(v_8184);
  assign v_8197 = mux_8197(v_8186);
  assign v_8198 = v_8199 & 1'h1;
  assign v_8199 = v_8200 & v_8201;
  assign v_8200 = ~act_8161;
  assign v_8201 = v_8202 | v_8206;
  assign v_8202 = v_8203 | v_8204;
  assign v_8203 = mux_8203(v_8102);
  assign v_8204 = mux_8204(v_8205);
  assign v_8205 = ~v_8102;
  assign v_8206 = ~v_8158;
  assign v_8207 = v_8208 | v_8209;
  assign v_8208 = mux_8208(v_8160);
  assign v_8209 = mux_8209(v_8198);
  assign v_8210 = v_8211 & 1'h1;
  assign v_8211 = v_8212 & v_8213;
  assign v_8212 = ~act_8101;
  assign v_8213 = v_8214 | v_8218;
  assign v_8214 = v_8215 | v_8216;
  assign v_8215 = mux_8215(v_7970);
  assign v_8216 = mux_8216(v_8217);
  assign v_8217 = ~v_7970;
  assign v_8218 = ~v_8098;
  assign v_8219 = v_8220 | v_8221;
  assign v_8220 = mux_8220(v_8100);
  assign v_8221 = mux_8221(v_8210);
  assign v_8222 = v_8223 & 1'h1;
  assign v_8223 = v_8224 & v_8225;
  assign v_8224 = ~act_7969;
  assign v_8225 = v_8226 | v_8230;
  assign v_8226 = v_8227 | v_8228;
  assign v_8227 = mux_8227(v_7694);
  assign v_8228 = mux_8228(v_8229);
  assign v_8229 = ~v_7694;
  assign v_8230 = ~v_7966;
  assign v_8231 = v_8232 | v_8233;
  assign v_8232 = mux_8232(v_7968);
  assign v_8233 = mux_8233(v_8222);
  assign v_8234 = v_8235 & 1'h1;
  assign v_8235 = v_8236 & v_8237;
  assign v_8236 = ~act_7693;
  assign v_8237 = v_8238 | v_8243;
  assign v_8238 = v_8239 | v_8241;
  assign v_8239 = mux_8239(v_8240);
  assign v_8240 = v_7690 & 1'h1;
  assign v_8241 = mux_8241(v_8242);
  assign v_8242 = ~v_8240;
  assign v_8243 = ~v_7690;
  assign v_8244 = v_8245 | v_8246;
  assign v_8245 = mux_8245(v_7692);
  assign v_8246 = mux_8246(v_8234);
  assign v_8248 = v_8249 | v_8791;
  assign v_8249 = act_8250 & 1'h1;
  assign act_8250 = v_8251 | v_8516;
  assign v_8251 = v_8252 & 1'h1;
  assign v_8252 = v_8253 & v_8523;
  assign v_8253 = ~v_8254;
  assign v_8255 = v_8256 | v_8510;
  assign v_8256 = act_8257 & 1'h1;
  assign act_8257 = v_8258 | v_8379;
  assign v_8258 = v_8259 & 1'h1;
  assign v_8259 = v_8260 & v_8386;
  assign v_8260 = ~v_8261;
  assign v_8262 = v_8263 | v_8373;
  assign v_8263 = act_8264 & 1'h1;
  assign act_8264 = v_8265 | v_8314;
  assign v_8265 = v_8266 & 1'h1;
  assign v_8266 = v_8267 & v_8321;
  assign v_8267 = ~v_8268;
  assign v_8269 = v_8270 | v_8308;
  assign v_8270 = act_8271 & 1'h1;
  assign act_8271 = v_8272 | v_8285;
  assign v_8272 = v_8273 & 1'h1;
  assign v_8273 = v_8274 & v_8292;
  assign v_8274 = ~v_8275;
  assign v_8276 = v_8277 | v_8279;
  assign v_8277 = act_8278 & 1'h1;
  assign act_8278 = v_1352 | v_1346;
  assign v_8279 = v_8280 & 1'h1;
  assign v_8280 = v_8281 & v_8282;
  assign v_8281 = ~act_8278;
  assign v_8282 = v_8283 | v_8288;
  assign v_8283 = v_8284 | v_8286;
  assign v_8284 = mux_8284(v_8285);
  assign v_8285 = v_8275 & 1'h1;
  assign v_8286 = mux_8286(v_8287);
  assign v_8287 = ~v_8285;
  assign v_8288 = ~v_8275;
  assign v_8289 = v_8290 | v_8291;
  assign v_8290 = mux_8290(v_8277);
  assign v_8291 = mux_8291(v_8279);
  assign v_8293 = v_8294 | v_8296;
  assign v_8294 = act_8295 & 1'h1;
  assign act_8295 = v_1366 | v_1360;
  assign v_8296 = v_8297 & 1'h1;
  assign v_8297 = v_8298 & v_8299;
  assign v_8298 = ~act_8295;
  assign v_8299 = v_8300 | v_8304;
  assign v_8300 = v_8301 | v_8302;
  assign v_8301 = mux_8301(v_8272);
  assign v_8302 = mux_8302(v_8303);
  assign v_8303 = ~v_8272;
  assign v_8304 = ~v_8292;
  assign v_8305 = v_8306 | v_8307;
  assign v_8306 = mux_8306(v_8294);
  assign v_8307 = mux_8307(v_8296);
  assign v_8308 = v_8309 & 1'h1;
  assign v_8309 = v_8310 & v_8311;
  assign v_8310 = ~act_8271;
  assign v_8311 = v_8312 | v_8317;
  assign v_8312 = v_8313 | v_8315;
  assign v_8313 = mux_8313(v_8314);
  assign v_8314 = v_8268 & 1'h1;
  assign v_8315 = mux_8315(v_8316);
  assign v_8316 = ~v_8314;
  assign v_8317 = ~v_8268;
  assign v_8318 = v_8319 | v_8320;
  assign v_8319 = mux_8319(v_8270);
  assign v_8320 = mux_8320(v_8308);
  assign v_8322 = v_8323 | v_8361;
  assign v_8323 = act_8324 & 1'h1;
  assign act_8324 = v_8325 | v_8338;
  assign v_8325 = v_8326 & 1'h1;
  assign v_8326 = v_8327 & v_8345;
  assign v_8327 = ~v_8328;
  assign v_8329 = v_8330 | v_8332;
  assign v_8330 = act_8331 & 1'h1;
  assign act_8331 = v_1380 | v_1374;
  assign v_8332 = v_8333 & 1'h1;
  assign v_8333 = v_8334 & v_8335;
  assign v_8334 = ~act_8331;
  assign v_8335 = v_8336 | v_8341;
  assign v_8336 = v_8337 | v_8339;
  assign v_8337 = mux_8337(v_8338);
  assign v_8338 = v_8328 & 1'h1;
  assign v_8339 = mux_8339(v_8340);
  assign v_8340 = ~v_8338;
  assign v_8341 = ~v_8328;
  assign v_8342 = v_8343 | v_8344;
  assign v_8343 = mux_8343(v_8330);
  assign v_8344 = mux_8344(v_8332);
  assign v_8346 = v_8347 | v_8349;
  assign v_8347 = act_8348 & 1'h1;
  assign act_8348 = v_1394 | v_1388;
  assign v_8349 = v_8350 & 1'h1;
  assign v_8350 = v_8351 & v_8352;
  assign v_8351 = ~act_8348;
  assign v_8352 = v_8353 | v_8357;
  assign v_8353 = v_8354 | v_8355;
  assign v_8354 = mux_8354(v_8325);
  assign v_8355 = mux_8355(v_8356);
  assign v_8356 = ~v_8325;
  assign v_8357 = ~v_8345;
  assign v_8358 = v_8359 | v_8360;
  assign v_8359 = mux_8359(v_8347);
  assign v_8360 = mux_8360(v_8349);
  assign v_8361 = v_8362 & 1'h1;
  assign v_8362 = v_8363 & v_8364;
  assign v_8363 = ~act_8324;
  assign v_8364 = v_8365 | v_8369;
  assign v_8365 = v_8366 | v_8367;
  assign v_8366 = mux_8366(v_8265);
  assign v_8367 = mux_8367(v_8368);
  assign v_8368 = ~v_8265;
  assign v_8369 = ~v_8321;
  assign v_8370 = v_8371 | v_8372;
  assign v_8371 = mux_8371(v_8323);
  assign v_8372 = mux_8372(v_8361);
  assign v_8373 = v_8374 & 1'h1;
  assign v_8374 = v_8375 & v_8376;
  assign v_8375 = ~act_8264;
  assign v_8376 = v_8377 | v_8382;
  assign v_8377 = v_8378 | v_8380;
  assign v_8378 = mux_8378(v_8379);
  assign v_8379 = v_8261 & 1'h1;
  assign v_8380 = mux_8380(v_8381);
  assign v_8381 = ~v_8379;
  assign v_8382 = ~v_8261;
  assign v_8383 = v_8384 | v_8385;
  assign v_8384 = mux_8384(v_8263);
  assign v_8385 = mux_8385(v_8373);
  assign v_8387 = v_8388 | v_8498;
  assign v_8388 = act_8389 & 1'h1;
  assign act_8389 = v_8390 | v_8439;
  assign v_8390 = v_8391 & 1'h1;
  assign v_8391 = v_8392 & v_8446;
  assign v_8392 = ~v_8393;
  assign v_8394 = v_8395 | v_8433;
  assign v_8395 = act_8396 & 1'h1;
  assign act_8396 = v_8397 | v_8410;
  assign v_8397 = v_8398 & 1'h1;
  assign v_8398 = v_8399 & v_8417;
  assign v_8399 = ~v_8400;
  assign v_8401 = v_8402 | v_8404;
  assign v_8402 = act_8403 & 1'h1;
  assign act_8403 = v_1408 | v_1402;
  assign v_8404 = v_8405 & 1'h1;
  assign v_8405 = v_8406 & v_8407;
  assign v_8406 = ~act_8403;
  assign v_8407 = v_8408 | v_8413;
  assign v_8408 = v_8409 | v_8411;
  assign v_8409 = mux_8409(v_8410);
  assign v_8410 = v_8400 & 1'h1;
  assign v_8411 = mux_8411(v_8412);
  assign v_8412 = ~v_8410;
  assign v_8413 = ~v_8400;
  assign v_8414 = v_8415 | v_8416;
  assign v_8415 = mux_8415(v_8402);
  assign v_8416 = mux_8416(v_8404);
  assign v_8418 = v_8419 | v_8421;
  assign v_8419 = act_8420 & 1'h1;
  assign act_8420 = v_1422 | v_1416;
  assign v_8421 = v_8422 & 1'h1;
  assign v_8422 = v_8423 & v_8424;
  assign v_8423 = ~act_8420;
  assign v_8424 = v_8425 | v_8429;
  assign v_8425 = v_8426 | v_8427;
  assign v_8426 = mux_8426(v_8397);
  assign v_8427 = mux_8427(v_8428);
  assign v_8428 = ~v_8397;
  assign v_8429 = ~v_8417;
  assign v_8430 = v_8431 | v_8432;
  assign v_8431 = mux_8431(v_8419);
  assign v_8432 = mux_8432(v_8421);
  assign v_8433 = v_8434 & 1'h1;
  assign v_8434 = v_8435 & v_8436;
  assign v_8435 = ~act_8396;
  assign v_8436 = v_8437 | v_8442;
  assign v_8437 = v_8438 | v_8440;
  assign v_8438 = mux_8438(v_8439);
  assign v_8439 = v_8393 & 1'h1;
  assign v_8440 = mux_8440(v_8441);
  assign v_8441 = ~v_8439;
  assign v_8442 = ~v_8393;
  assign v_8443 = v_8444 | v_8445;
  assign v_8444 = mux_8444(v_8395);
  assign v_8445 = mux_8445(v_8433);
  assign v_8447 = v_8448 | v_8486;
  assign v_8448 = act_8449 & 1'h1;
  assign act_8449 = v_8450 | v_8463;
  assign v_8450 = v_8451 & 1'h1;
  assign v_8451 = v_8452 & v_8470;
  assign v_8452 = ~v_8453;
  assign v_8454 = v_8455 | v_8457;
  assign v_8455 = act_8456 & 1'h1;
  assign act_8456 = v_1436 | v_1430;
  assign v_8457 = v_8458 & 1'h1;
  assign v_8458 = v_8459 & v_8460;
  assign v_8459 = ~act_8456;
  assign v_8460 = v_8461 | v_8466;
  assign v_8461 = v_8462 | v_8464;
  assign v_8462 = mux_8462(v_8463);
  assign v_8463 = v_8453 & 1'h1;
  assign v_8464 = mux_8464(v_8465);
  assign v_8465 = ~v_8463;
  assign v_8466 = ~v_8453;
  assign v_8467 = v_8468 | v_8469;
  assign v_8468 = mux_8468(v_8455);
  assign v_8469 = mux_8469(v_8457);
  assign v_8471 = v_8472 | v_8474;
  assign v_8472 = act_8473 & 1'h1;
  assign act_8473 = v_1450 | v_1444;
  assign v_8474 = v_8475 & 1'h1;
  assign v_8475 = v_8476 & v_8477;
  assign v_8476 = ~act_8473;
  assign v_8477 = v_8478 | v_8482;
  assign v_8478 = v_8479 | v_8480;
  assign v_8479 = mux_8479(v_8450);
  assign v_8480 = mux_8480(v_8481);
  assign v_8481 = ~v_8450;
  assign v_8482 = ~v_8470;
  assign v_8483 = v_8484 | v_8485;
  assign v_8484 = mux_8484(v_8472);
  assign v_8485 = mux_8485(v_8474);
  assign v_8486 = v_8487 & 1'h1;
  assign v_8487 = v_8488 & v_8489;
  assign v_8488 = ~act_8449;
  assign v_8489 = v_8490 | v_8494;
  assign v_8490 = v_8491 | v_8492;
  assign v_8491 = mux_8491(v_8390);
  assign v_8492 = mux_8492(v_8493);
  assign v_8493 = ~v_8390;
  assign v_8494 = ~v_8446;
  assign v_8495 = v_8496 | v_8497;
  assign v_8496 = mux_8496(v_8448);
  assign v_8497 = mux_8497(v_8486);
  assign v_8498 = v_8499 & 1'h1;
  assign v_8499 = v_8500 & v_8501;
  assign v_8500 = ~act_8389;
  assign v_8501 = v_8502 | v_8506;
  assign v_8502 = v_8503 | v_8504;
  assign v_8503 = mux_8503(v_8258);
  assign v_8504 = mux_8504(v_8505);
  assign v_8505 = ~v_8258;
  assign v_8506 = ~v_8386;
  assign v_8507 = v_8508 | v_8509;
  assign v_8508 = mux_8508(v_8388);
  assign v_8509 = mux_8509(v_8498);
  assign v_8510 = v_8511 & 1'h1;
  assign v_8511 = v_8512 & v_8513;
  assign v_8512 = ~act_8257;
  assign v_8513 = v_8514 | v_8519;
  assign v_8514 = v_8515 | v_8517;
  assign v_8515 = mux_8515(v_8516);
  assign v_8516 = v_8254 & 1'h1;
  assign v_8517 = mux_8517(v_8518);
  assign v_8518 = ~v_8516;
  assign v_8519 = ~v_8254;
  assign v_8520 = v_8521 | v_8522;
  assign v_8521 = mux_8521(v_8256);
  assign v_8522 = mux_8522(v_8510);
  assign v_8524 = v_8525 | v_8779;
  assign v_8525 = act_8526 & 1'h1;
  assign act_8526 = v_8527 | v_8648;
  assign v_8527 = v_8528 & 1'h1;
  assign v_8528 = v_8529 & v_8655;
  assign v_8529 = ~v_8530;
  assign v_8531 = v_8532 | v_8642;
  assign v_8532 = act_8533 & 1'h1;
  assign act_8533 = v_8534 | v_8583;
  assign v_8534 = v_8535 & 1'h1;
  assign v_8535 = v_8536 & v_8590;
  assign v_8536 = ~v_8537;
  assign v_8538 = v_8539 | v_8577;
  assign v_8539 = act_8540 & 1'h1;
  assign act_8540 = v_8541 | v_8554;
  assign v_8541 = v_8542 & 1'h1;
  assign v_8542 = v_8543 & v_8561;
  assign v_8543 = ~v_8544;
  assign v_8545 = v_8546 | v_8548;
  assign v_8546 = act_8547 & 1'h1;
  assign act_8547 = v_1464 | v_1458;
  assign v_8548 = v_8549 & 1'h1;
  assign v_8549 = v_8550 & v_8551;
  assign v_8550 = ~act_8547;
  assign v_8551 = v_8552 | v_8557;
  assign v_8552 = v_8553 | v_8555;
  assign v_8553 = mux_8553(v_8554);
  assign v_8554 = v_8544 & 1'h1;
  assign v_8555 = mux_8555(v_8556);
  assign v_8556 = ~v_8554;
  assign v_8557 = ~v_8544;
  assign v_8558 = v_8559 | v_8560;
  assign v_8559 = mux_8559(v_8546);
  assign v_8560 = mux_8560(v_8548);
  assign v_8562 = v_8563 | v_8565;
  assign v_8563 = act_8564 & 1'h1;
  assign act_8564 = v_1478 | v_1472;
  assign v_8565 = v_8566 & 1'h1;
  assign v_8566 = v_8567 & v_8568;
  assign v_8567 = ~act_8564;
  assign v_8568 = v_8569 | v_8573;
  assign v_8569 = v_8570 | v_8571;
  assign v_8570 = mux_8570(v_8541);
  assign v_8571 = mux_8571(v_8572);
  assign v_8572 = ~v_8541;
  assign v_8573 = ~v_8561;
  assign v_8574 = v_8575 | v_8576;
  assign v_8575 = mux_8575(v_8563);
  assign v_8576 = mux_8576(v_8565);
  assign v_8577 = v_8578 & 1'h1;
  assign v_8578 = v_8579 & v_8580;
  assign v_8579 = ~act_8540;
  assign v_8580 = v_8581 | v_8586;
  assign v_8581 = v_8582 | v_8584;
  assign v_8582 = mux_8582(v_8583);
  assign v_8583 = v_8537 & 1'h1;
  assign v_8584 = mux_8584(v_8585);
  assign v_8585 = ~v_8583;
  assign v_8586 = ~v_8537;
  assign v_8587 = v_8588 | v_8589;
  assign v_8588 = mux_8588(v_8539);
  assign v_8589 = mux_8589(v_8577);
  assign v_8591 = v_8592 | v_8630;
  assign v_8592 = act_8593 & 1'h1;
  assign act_8593 = v_8594 | v_8607;
  assign v_8594 = v_8595 & 1'h1;
  assign v_8595 = v_8596 & v_8614;
  assign v_8596 = ~v_8597;
  assign v_8598 = v_8599 | v_8601;
  assign v_8599 = act_8600 & 1'h1;
  assign act_8600 = v_1492 | v_1486;
  assign v_8601 = v_8602 & 1'h1;
  assign v_8602 = v_8603 & v_8604;
  assign v_8603 = ~act_8600;
  assign v_8604 = v_8605 | v_8610;
  assign v_8605 = v_8606 | v_8608;
  assign v_8606 = mux_8606(v_8607);
  assign v_8607 = v_8597 & 1'h1;
  assign v_8608 = mux_8608(v_8609);
  assign v_8609 = ~v_8607;
  assign v_8610 = ~v_8597;
  assign v_8611 = v_8612 | v_8613;
  assign v_8612 = mux_8612(v_8599);
  assign v_8613 = mux_8613(v_8601);
  assign v_8615 = v_8616 | v_8618;
  assign v_8616 = act_8617 & 1'h1;
  assign act_8617 = v_1506 | v_1500;
  assign v_8618 = v_8619 & 1'h1;
  assign v_8619 = v_8620 & v_8621;
  assign v_8620 = ~act_8617;
  assign v_8621 = v_8622 | v_8626;
  assign v_8622 = v_8623 | v_8624;
  assign v_8623 = mux_8623(v_8594);
  assign v_8624 = mux_8624(v_8625);
  assign v_8625 = ~v_8594;
  assign v_8626 = ~v_8614;
  assign v_8627 = v_8628 | v_8629;
  assign v_8628 = mux_8628(v_8616);
  assign v_8629 = mux_8629(v_8618);
  assign v_8630 = v_8631 & 1'h1;
  assign v_8631 = v_8632 & v_8633;
  assign v_8632 = ~act_8593;
  assign v_8633 = v_8634 | v_8638;
  assign v_8634 = v_8635 | v_8636;
  assign v_8635 = mux_8635(v_8534);
  assign v_8636 = mux_8636(v_8637);
  assign v_8637 = ~v_8534;
  assign v_8638 = ~v_8590;
  assign v_8639 = v_8640 | v_8641;
  assign v_8640 = mux_8640(v_8592);
  assign v_8641 = mux_8641(v_8630);
  assign v_8642 = v_8643 & 1'h1;
  assign v_8643 = v_8644 & v_8645;
  assign v_8644 = ~act_8533;
  assign v_8645 = v_8646 | v_8651;
  assign v_8646 = v_8647 | v_8649;
  assign v_8647 = mux_8647(v_8648);
  assign v_8648 = v_8530 & 1'h1;
  assign v_8649 = mux_8649(v_8650);
  assign v_8650 = ~v_8648;
  assign v_8651 = ~v_8530;
  assign v_8652 = v_8653 | v_8654;
  assign v_8653 = mux_8653(v_8532);
  assign v_8654 = mux_8654(v_8642);
  assign v_8656 = v_8657 | v_8767;
  assign v_8657 = act_8658 & 1'h1;
  assign act_8658 = v_8659 | v_8708;
  assign v_8659 = v_8660 & 1'h1;
  assign v_8660 = v_8661 & v_8715;
  assign v_8661 = ~v_8662;
  assign v_8663 = v_8664 | v_8702;
  assign v_8664 = act_8665 & 1'h1;
  assign act_8665 = v_8666 | v_8679;
  assign v_8666 = v_8667 & 1'h1;
  assign v_8667 = v_8668 & v_8686;
  assign v_8668 = ~v_8669;
  assign v_8670 = v_8671 | v_8673;
  assign v_8671 = act_8672 & 1'h1;
  assign act_8672 = v_1520 | v_1514;
  assign v_8673 = v_8674 & 1'h1;
  assign v_8674 = v_8675 & v_8676;
  assign v_8675 = ~act_8672;
  assign v_8676 = v_8677 | v_8682;
  assign v_8677 = v_8678 | v_8680;
  assign v_8678 = mux_8678(v_8679);
  assign v_8679 = v_8669 & 1'h1;
  assign v_8680 = mux_8680(v_8681);
  assign v_8681 = ~v_8679;
  assign v_8682 = ~v_8669;
  assign v_8683 = v_8684 | v_8685;
  assign v_8684 = mux_8684(v_8671);
  assign v_8685 = mux_8685(v_8673);
  assign v_8687 = v_8688 | v_8690;
  assign v_8688 = act_8689 & 1'h1;
  assign act_8689 = v_1534 | v_1528;
  assign v_8690 = v_8691 & 1'h1;
  assign v_8691 = v_8692 & v_8693;
  assign v_8692 = ~act_8689;
  assign v_8693 = v_8694 | v_8698;
  assign v_8694 = v_8695 | v_8696;
  assign v_8695 = mux_8695(v_8666);
  assign v_8696 = mux_8696(v_8697);
  assign v_8697 = ~v_8666;
  assign v_8698 = ~v_8686;
  assign v_8699 = v_8700 | v_8701;
  assign v_8700 = mux_8700(v_8688);
  assign v_8701 = mux_8701(v_8690);
  assign v_8702 = v_8703 & 1'h1;
  assign v_8703 = v_8704 & v_8705;
  assign v_8704 = ~act_8665;
  assign v_8705 = v_8706 | v_8711;
  assign v_8706 = v_8707 | v_8709;
  assign v_8707 = mux_8707(v_8708);
  assign v_8708 = v_8662 & 1'h1;
  assign v_8709 = mux_8709(v_8710);
  assign v_8710 = ~v_8708;
  assign v_8711 = ~v_8662;
  assign v_8712 = v_8713 | v_8714;
  assign v_8713 = mux_8713(v_8664);
  assign v_8714 = mux_8714(v_8702);
  assign v_8716 = v_8717 | v_8755;
  assign v_8717 = act_8718 & 1'h1;
  assign act_8718 = v_8719 | v_8732;
  assign v_8719 = v_8720 & 1'h1;
  assign v_8720 = v_8721 & v_8739;
  assign v_8721 = ~v_8722;
  assign v_8723 = v_8724 | v_8726;
  assign v_8724 = act_8725 & 1'h1;
  assign act_8725 = v_1548 | v_1542;
  assign v_8726 = v_8727 & 1'h1;
  assign v_8727 = v_8728 & v_8729;
  assign v_8728 = ~act_8725;
  assign v_8729 = v_8730 | v_8735;
  assign v_8730 = v_8731 | v_8733;
  assign v_8731 = mux_8731(v_8732);
  assign v_8732 = v_8722 & 1'h1;
  assign v_8733 = mux_8733(v_8734);
  assign v_8734 = ~v_8732;
  assign v_8735 = ~v_8722;
  assign v_8736 = v_8737 | v_8738;
  assign v_8737 = mux_8737(v_8724);
  assign v_8738 = mux_8738(v_8726);
  assign v_8740 = v_8741 | v_8743;
  assign v_8741 = act_8742 & 1'h1;
  assign act_8742 = v_1562 | v_1556;
  assign v_8743 = v_8744 & 1'h1;
  assign v_8744 = v_8745 & v_8746;
  assign v_8745 = ~act_8742;
  assign v_8746 = v_8747 | v_8751;
  assign v_8747 = v_8748 | v_8749;
  assign v_8748 = mux_8748(v_8719);
  assign v_8749 = mux_8749(v_8750);
  assign v_8750 = ~v_8719;
  assign v_8751 = ~v_8739;
  assign v_8752 = v_8753 | v_8754;
  assign v_8753 = mux_8753(v_8741);
  assign v_8754 = mux_8754(v_8743);
  assign v_8755 = v_8756 & 1'h1;
  assign v_8756 = v_8757 & v_8758;
  assign v_8757 = ~act_8718;
  assign v_8758 = v_8759 | v_8763;
  assign v_8759 = v_8760 | v_8761;
  assign v_8760 = mux_8760(v_8659);
  assign v_8761 = mux_8761(v_8762);
  assign v_8762 = ~v_8659;
  assign v_8763 = ~v_8715;
  assign v_8764 = v_8765 | v_8766;
  assign v_8765 = mux_8765(v_8717);
  assign v_8766 = mux_8766(v_8755);
  assign v_8767 = v_8768 & 1'h1;
  assign v_8768 = v_8769 & v_8770;
  assign v_8769 = ~act_8658;
  assign v_8770 = v_8771 | v_8775;
  assign v_8771 = v_8772 | v_8773;
  assign v_8772 = mux_8772(v_8527);
  assign v_8773 = mux_8773(v_8774);
  assign v_8774 = ~v_8527;
  assign v_8775 = ~v_8655;
  assign v_8776 = v_8777 | v_8778;
  assign v_8777 = mux_8777(v_8657);
  assign v_8778 = mux_8778(v_8767);
  assign v_8779 = v_8780 & 1'h1;
  assign v_8780 = v_8781 & v_8782;
  assign v_8781 = ~act_8526;
  assign v_8782 = v_8783 | v_8787;
  assign v_8783 = v_8784 | v_8785;
  assign v_8784 = mux_8784(v_8251);
  assign v_8785 = mux_8785(v_8786);
  assign v_8786 = ~v_8251;
  assign v_8787 = ~v_8523;
  assign v_8788 = v_8789 | v_8790;
  assign v_8789 = mux_8789(v_8525);
  assign v_8790 = mux_8790(v_8779);
  assign v_8791 = v_8792 & 1'h1;
  assign v_8792 = v_8793 & v_8794;
  assign v_8793 = ~act_8250;
  assign v_8794 = v_8795 | v_8799;
  assign v_8795 = v_8796 | v_8797;
  assign v_8796 = mux_8796(v_7687);
  assign v_8797 = mux_8797(v_8798);
  assign v_8798 = ~v_7687;
  assign v_8799 = ~v_8247;
  assign v_8800 = v_8801 | v_8802;
  assign v_8801 = mux_8801(v_8249);
  assign v_8802 = mux_8802(v_8791);
  assign v_8803 = v_8804 & 1'h1;
  assign v_8804 = v_8805 & v_8806;
  assign v_8805 = ~act_7686;
  assign v_8806 = v_8807 | v_8812;
  assign v_8807 = v_8808 | v_8810;
  assign v_8808 = mux_8808(v_8809);
  assign v_8809 = v_7683 & 1'h1;
  assign v_8810 = mux_8810(v_8811);
  assign v_8811 = ~v_8809;
  assign v_8812 = ~v_7683;
  assign v_8813 = v_8814 | v_8815;
  assign v_8814 = mux_8814(v_7685);
  assign v_8815 = mux_8815(v_8803);
  assign v_8817 = v_8818 | v_9936;
  assign v_8818 = act_8819 & 1'h1;
  assign act_8819 = v_8820 | v_9373;
  assign v_8820 = v_8821 & 1'h1;
  assign v_8821 = v_8822 & v_9380;
  assign v_8822 = ~v_8823;
  assign v_8824 = v_8825 | v_9367;
  assign v_8825 = act_8826 & 1'h1;
  assign act_8826 = v_8827 | v_9092;
  assign v_8827 = v_8828 & 1'h1;
  assign v_8828 = v_8829 & v_9099;
  assign v_8829 = ~v_8830;
  assign v_8831 = v_8832 | v_9086;
  assign v_8832 = act_8833 & 1'h1;
  assign act_8833 = v_8834 | v_8955;
  assign v_8834 = v_8835 & 1'h1;
  assign v_8835 = v_8836 & v_8962;
  assign v_8836 = ~v_8837;
  assign v_8838 = v_8839 | v_8949;
  assign v_8839 = act_8840 & 1'h1;
  assign act_8840 = v_8841 | v_8890;
  assign v_8841 = v_8842 & 1'h1;
  assign v_8842 = v_8843 & v_8897;
  assign v_8843 = ~v_8844;
  assign v_8845 = v_8846 | v_8884;
  assign v_8846 = act_8847 & 1'h1;
  assign act_8847 = v_8848 | v_8861;
  assign v_8848 = v_8849 & 1'h1;
  assign v_8849 = v_8850 & v_8868;
  assign v_8850 = ~v_8851;
  assign v_8852 = v_8853 | v_8855;
  assign v_8853 = act_8854 & 1'h1;
  assign act_8854 = v_1576 | v_1570;
  assign v_8855 = v_8856 & 1'h1;
  assign v_8856 = v_8857 & v_8858;
  assign v_8857 = ~act_8854;
  assign v_8858 = v_8859 | v_8864;
  assign v_8859 = v_8860 | v_8862;
  assign v_8860 = mux_8860(v_8861);
  assign v_8861 = v_8851 & 1'h1;
  assign v_8862 = mux_8862(v_8863);
  assign v_8863 = ~v_8861;
  assign v_8864 = ~v_8851;
  assign v_8865 = v_8866 | v_8867;
  assign v_8866 = mux_8866(v_8853);
  assign v_8867 = mux_8867(v_8855);
  assign v_8869 = v_8870 | v_8872;
  assign v_8870 = act_8871 & 1'h1;
  assign act_8871 = v_1590 | v_1584;
  assign v_8872 = v_8873 & 1'h1;
  assign v_8873 = v_8874 & v_8875;
  assign v_8874 = ~act_8871;
  assign v_8875 = v_8876 | v_8880;
  assign v_8876 = v_8877 | v_8878;
  assign v_8877 = mux_8877(v_8848);
  assign v_8878 = mux_8878(v_8879);
  assign v_8879 = ~v_8848;
  assign v_8880 = ~v_8868;
  assign v_8881 = v_8882 | v_8883;
  assign v_8882 = mux_8882(v_8870);
  assign v_8883 = mux_8883(v_8872);
  assign v_8884 = v_8885 & 1'h1;
  assign v_8885 = v_8886 & v_8887;
  assign v_8886 = ~act_8847;
  assign v_8887 = v_8888 | v_8893;
  assign v_8888 = v_8889 | v_8891;
  assign v_8889 = mux_8889(v_8890);
  assign v_8890 = v_8844 & 1'h1;
  assign v_8891 = mux_8891(v_8892);
  assign v_8892 = ~v_8890;
  assign v_8893 = ~v_8844;
  assign v_8894 = v_8895 | v_8896;
  assign v_8895 = mux_8895(v_8846);
  assign v_8896 = mux_8896(v_8884);
  assign v_8898 = v_8899 | v_8937;
  assign v_8899 = act_8900 & 1'h1;
  assign act_8900 = v_8901 | v_8914;
  assign v_8901 = v_8902 & 1'h1;
  assign v_8902 = v_8903 & v_8921;
  assign v_8903 = ~v_8904;
  assign v_8905 = v_8906 | v_8908;
  assign v_8906 = act_8907 & 1'h1;
  assign act_8907 = v_1604 | v_1598;
  assign v_8908 = v_8909 & 1'h1;
  assign v_8909 = v_8910 & v_8911;
  assign v_8910 = ~act_8907;
  assign v_8911 = v_8912 | v_8917;
  assign v_8912 = v_8913 | v_8915;
  assign v_8913 = mux_8913(v_8914);
  assign v_8914 = v_8904 & 1'h1;
  assign v_8915 = mux_8915(v_8916);
  assign v_8916 = ~v_8914;
  assign v_8917 = ~v_8904;
  assign v_8918 = v_8919 | v_8920;
  assign v_8919 = mux_8919(v_8906);
  assign v_8920 = mux_8920(v_8908);
  assign v_8922 = v_8923 | v_8925;
  assign v_8923 = act_8924 & 1'h1;
  assign act_8924 = v_1618 | v_1612;
  assign v_8925 = v_8926 & 1'h1;
  assign v_8926 = v_8927 & v_8928;
  assign v_8927 = ~act_8924;
  assign v_8928 = v_8929 | v_8933;
  assign v_8929 = v_8930 | v_8931;
  assign v_8930 = mux_8930(v_8901);
  assign v_8931 = mux_8931(v_8932);
  assign v_8932 = ~v_8901;
  assign v_8933 = ~v_8921;
  assign v_8934 = v_8935 | v_8936;
  assign v_8935 = mux_8935(v_8923);
  assign v_8936 = mux_8936(v_8925);
  assign v_8937 = v_8938 & 1'h1;
  assign v_8938 = v_8939 & v_8940;
  assign v_8939 = ~act_8900;
  assign v_8940 = v_8941 | v_8945;
  assign v_8941 = v_8942 | v_8943;
  assign v_8942 = mux_8942(v_8841);
  assign v_8943 = mux_8943(v_8944);
  assign v_8944 = ~v_8841;
  assign v_8945 = ~v_8897;
  assign v_8946 = v_8947 | v_8948;
  assign v_8947 = mux_8947(v_8899);
  assign v_8948 = mux_8948(v_8937);
  assign v_8949 = v_8950 & 1'h1;
  assign v_8950 = v_8951 & v_8952;
  assign v_8951 = ~act_8840;
  assign v_8952 = v_8953 | v_8958;
  assign v_8953 = v_8954 | v_8956;
  assign v_8954 = mux_8954(v_8955);
  assign v_8955 = v_8837 & 1'h1;
  assign v_8956 = mux_8956(v_8957);
  assign v_8957 = ~v_8955;
  assign v_8958 = ~v_8837;
  assign v_8959 = v_8960 | v_8961;
  assign v_8960 = mux_8960(v_8839);
  assign v_8961 = mux_8961(v_8949);
  assign v_8963 = v_8964 | v_9074;
  assign v_8964 = act_8965 & 1'h1;
  assign act_8965 = v_8966 | v_9015;
  assign v_8966 = v_8967 & 1'h1;
  assign v_8967 = v_8968 & v_9022;
  assign v_8968 = ~v_8969;
  assign v_8970 = v_8971 | v_9009;
  assign v_8971 = act_8972 & 1'h1;
  assign act_8972 = v_8973 | v_8986;
  assign v_8973 = v_8974 & 1'h1;
  assign v_8974 = v_8975 & v_8993;
  assign v_8975 = ~v_8976;
  assign v_8977 = v_8978 | v_8980;
  assign v_8978 = act_8979 & 1'h1;
  assign act_8979 = v_1632 | v_1626;
  assign v_8980 = v_8981 & 1'h1;
  assign v_8981 = v_8982 & v_8983;
  assign v_8982 = ~act_8979;
  assign v_8983 = v_8984 | v_8989;
  assign v_8984 = v_8985 | v_8987;
  assign v_8985 = mux_8985(v_8986);
  assign v_8986 = v_8976 & 1'h1;
  assign v_8987 = mux_8987(v_8988);
  assign v_8988 = ~v_8986;
  assign v_8989 = ~v_8976;
  assign v_8990 = v_8991 | v_8992;
  assign v_8991 = mux_8991(v_8978);
  assign v_8992 = mux_8992(v_8980);
  assign v_8994 = v_8995 | v_8997;
  assign v_8995 = act_8996 & 1'h1;
  assign act_8996 = v_1646 | v_1640;
  assign v_8997 = v_8998 & 1'h1;
  assign v_8998 = v_8999 & v_9000;
  assign v_8999 = ~act_8996;
  assign v_9000 = v_9001 | v_9005;
  assign v_9001 = v_9002 | v_9003;
  assign v_9002 = mux_9002(v_8973);
  assign v_9003 = mux_9003(v_9004);
  assign v_9004 = ~v_8973;
  assign v_9005 = ~v_8993;
  assign v_9006 = v_9007 | v_9008;
  assign v_9007 = mux_9007(v_8995);
  assign v_9008 = mux_9008(v_8997);
  assign v_9009 = v_9010 & 1'h1;
  assign v_9010 = v_9011 & v_9012;
  assign v_9011 = ~act_8972;
  assign v_9012 = v_9013 | v_9018;
  assign v_9013 = v_9014 | v_9016;
  assign v_9014 = mux_9014(v_9015);
  assign v_9015 = v_8969 & 1'h1;
  assign v_9016 = mux_9016(v_9017);
  assign v_9017 = ~v_9015;
  assign v_9018 = ~v_8969;
  assign v_9019 = v_9020 | v_9021;
  assign v_9020 = mux_9020(v_8971);
  assign v_9021 = mux_9021(v_9009);
  assign v_9023 = v_9024 | v_9062;
  assign v_9024 = act_9025 & 1'h1;
  assign act_9025 = v_9026 | v_9039;
  assign v_9026 = v_9027 & 1'h1;
  assign v_9027 = v_9028 & v_9046;
  assign v_9028 = ~v_9029;
  assign v_9030 = v_9031 | v_9033;
  assign v_9031 = act_9032 & 1'h1;
  assign act_9032 = v_1660 | v_1654;
  assign v_9033 = v_9034 & 1'h1;
  assign v_9034 = v_9035 & v_9036;
  assign v_9035 = ~act_9032;
  assign v_9036 = v_9037 | v_9042;
  assign v_9037 = v_9038 | v_9040;
  assign v_9038 = mux_9038(v_9039);
  assign v_9039 = v_9029 & 1'h1;
  assign v_9040 = mux_9040(v_9041);
  assign v_9041 = ~v_9039;
  assign v_9042 = ~v_9029;
  assign v_9043 = v_9044 | v_9045;
  assign v_9044 = mux_9044(v_9031);
  assign v_9045 = mux_9045(v_9033);
  assign v_9047 = v_9048 | v_9050;
  assign v_9048 = act_9049 & 1'h1;
  assign act_9049 = v_1674 | v_1668;
  assign v_9050 = v_9051 & 1'h1;
  assign v_9051 = v_9052 & v_9053;
  assign v_9052 = ~act_9049;
  assign v_9053 = v_9054 | v_9058;
  assign v_9054 = v_9055 | v_9056;
  assign v_9055 = mux_9055(v_9026);
  assign v_9056 = mux_9056(v_9057);
  assign v_9057 = ~v_9026;
  assign v_9058 = ~v_9046;
  assign v_9059 = v_9060 | v_9061;
  assign v_9060 = mux_9060(v_9048);
  assign v_9061 = mux_9061(v_9050);
  assign v_9062 = v_9063 & 1'h1;
  assign v_9063 = v_9064 & v_9065;
  assign v_9064 = ~act_9025;
  assign v_9065 = v_9066 | v_9070;
  assign v_9066 = v_9067 | v_9068;
  assign v_9067 = mux_9067(v_8966);
  assign v_9068 = mux_9068(v_9069);
  assign v_9069 = ~v_8966;
  assign v_9070 = ~v_9022;
  assign v_9071 = v_9072 | v_9073;
  assign v_9072 = mux_9072(v_9024);
  assign v_9073 = mux_9073(v_9062);
  assign v_9074 = v_9075 & 1'h1;
  assign v_9075 = v_9076 & v_9077;
  assign v_9076 = ~act_8965;
  assign v_9077 = v_9078 | v_9082;
  assign v_9078 = v_9079 | v_9080;
  assign v_9079 = mux_9079(v_8834);
  assign v_9080 = mux_9080(v_9081);
  assign v_9081 = ~v_8834;
  assign v_9082 = ~v_8962;
  assign v_9083 = v_9084 | v_9085;
  assign v_9084 = mux_9084(v_8964);
  assign v_9085 = mux_9085(v_9074);
  assign v_9086 = v_9087 & 1'h1;
  assign v_9087 = v_9088 & v_9089;
  assign v_9088 = ~act_8833;
  assign v_9089 = v_9090 | v_9095;
  assign v_9090 = v_9091 | v_9093;
  assign v_9091 = mux_9091(v_9092);
  assign v_9092 = v_8830 & 1'h1;
  assign v_9093 = mux_9093(v_9094);
  assign v_9094 = ~v_9092;
  assign v_9095 = ~v_8830;
  assign v_9096 = v_9097 | v_9098;
  assign v_9097 = mux_9097(v_8832);
  assign v_9098 = mux_9098(v_9086);
  assign v_9100 = v_9101 | v_9355;
  assign v_9101 = act_9102 & 1'h1;
  assign act_9102 = v_9103 | v_9224;
  assign v_9103 = v_9104 & 1'h1;
  assign v_9104 = v_9105 & v_9231;
  assign v_9105 = ~v_9106;
  assign v_9107 = v_9108 | v_9218;
  assign v_9108 = act_9109 & 1'h1;
  assign act_9109 = v_9110 | v_9159;
  assign v_9110 = v_9111 & 1'h1;
  assign v_9111 = v_9112 & v_9166;
  assign v_9112 = ~v_9113;
  assign v_9114 = v_9115 | v_9153;
  assign v_9115 = act_9116 & 1'h1;
  assign act_9116 = v_9117 | v_9130;
  assign v_9117 = v_9118 & 1'h1;
  assign v_9118 = v_9119 & v_9137;
  assign v_9119 = ~v_9120;
  assign v_9121 = v_9122 | v_9124;
  assign v_9122 = act_9123 & 1'h1;
  assign act_9123 = v_1688 | v_1682;
  assign v_9124 = v_9125 & 1'h1;
  assign v_9125 = v_9126 & v_9127;
  assign v_9126 = ~act_9123;
  assign v_9127 = v_9128 | v_9133;
  assign v_9128 = v_9129 | v_9131;
  assign v_9129 = mux_9129(v_9130);
  assign v_9130 = v_9120 & 1'h1;
  assign v_9131 = mux_9131(v_9132);
  assign v_9132 = ~v_9130;
  assign v_9133 = ~v_9120;
  assign v_9134 = v_9135 | v_9136;
  assign v_9135 = mux_9135(v_9122);
  assign v_9136 = mux_9136(v_9124);
  assign v_9138 = v_9139 | v_9141;
  assign v_9139 = act_9140 & 1'h1;
  assign act_9140 = v_1702 | v_1696;
  assign v_9141 = v_9142 & 1'h1;
  assign v_9142 = v_9143 & v_9144;
  assign v_9143 = ~act_9140;
  assign v_9144 = v_9145 | v_9149;
  assign v_9145 = v_9146 | v_9147;
  assign v_9146 = mux_9146(v_9117);
  assign v_9147 = mux_9147(v_9148);
  assign v_9148 = ~v_9117;
  assign v_9149 = ~v_9137;
  assign v_9150 = v_9151 | v_9152;
  assign v_9151 = mux_9151(v_9139);
  assign v_9152 = mux_9152(v_9141);
  assign v_9153 = v_9154 & 1'h1;
  assign v_9154 = v_9155 & v_9156;
  assign v_9155 = ~act_9116;
  assign v_9156 = v_9157 | v_9162;
  assign v_9157 = v_9158 | v_9160;
  assign v_9158 = mux_9158(v_9159);
  assign v_9159 = v_9113 & 1'h1;
  assign v_9160 = mux_9160(v_9161);
  assign v_9161 = ~v_9159;
  assign v_9162 = ~v_9113;
  assign v_9163 = v_9164 | v_9165;
  assign v_9164 = mux_9164(v_9115);
  assign v_9165 = mux_9165(v_9153);
  assign v_9167 = v_9168 | v_9206;
  assign v_9168 = act_9169 & 1'h1;
  assign act_9169 = v_9170 | v_9183;
  assign v_9170 = v_9171 & 1'h1;
  assign v_9171 = v_9172 & v_9190;
  assign v_9172 = ~v_9173;
  assign v_9174 = v_9175 | v_9177;
  assign v_9175 = act_9176 & 1'h1;
  assign act_9176 = v_1716 | v_1710;
  assign v_9177 = v_9178 & 1'h1;
  assign v_9178 = v_9179 & v_9180;
  assign v_9179 = ~act_9176;
  assign v_9180 = v_9181 | v_9186;
  assign v_9181 = v_9182 | v_9184;
  assign v_9182 = mux_9182(v_9183);
  assign v_9183 = v_9173 & 1'h1;
  assign v_9184 = mux_9184(v_9185);
  assign v_9185 = ~v_9183;
  assign v_9186 = ~v_9173;
  assign v_9187 = v_9188 | v_9189;
  assign v_9188 = mux_9188(v_9175);
  assign v_9189 = mux_9189(v_9177);
  assign v_9191 = v_9192 | v_9194;
  assign v_9192 = act_9193 & 1'h1;
  assign act_9193 = v_1730 | v_1724;
  assign v_9194 = v_9195 & 1'h1;
  assign v_9195 = v_9196 & v_9197;
  assign v_9196 = ~act_9193;
  assign v_9197 = v_9198 | v_9202;
  assign v_9198 = v_9199 | v_9200;
  assign v_9199 = mux_9199(v_9170);
  assign v_9200 = mux_9200(v_9201);
  assign v_9201 = ~v_9170;
  assign v_9202 = ~v_9190;
  assign v_9203 = v_9204 | v_9205;
  assign v_9204 = mux_9204(v_9192);
  assign v_9205 = mux_9205(v_9194);
  assign v_9206 = v_9207 & 1'h1;
  assign v_9207 = v_9208 & v_9209;
  assign v_9208 = ~act_9169;
  assign v_9209 = v_9210 | v_9214;
  assign v_9210 = v_9211 | v_9212;
  assign v_9211 = mux_9211(v_9110);
  assign v_9212 = mux_9212(v_9213);
  assign v_9213 = ~v_9110;
  assign v_9214 = ~v_9166;
  assign v_9215 = v_9216 | v_9217;
  assign v_9216 = mux_9216(v_9168);
  assign v_9217 = mux_9217(v_9206);
  assign v_9218 = v_9219 & 1'h1;
  assign v_9219 = v_9220 & v_9221;
  assign v_9220 = ~act_9109;
  assign v_9221 = v_9222 | v_9227;
  assign v_9222 = v_9223 | v_9225;
  assign v_9223 = mux_9223(v_9224);
  assign v_9224 = v_9106 & 1'h1;
  assign v_9225 = mux_9225(v_9226);
  assign v_9226 = ~v_9224;
  assign v_9227 = ~v_9106;
  assign v_9228 = v_9229 | v_9230;
  assign v_9229 = mux_9229(v_9108);
  assign v_9230 = mux_9230(v_9218);
  assign v_9232 = v_9233 | v_9343;
  assign v_9233 = act_9234 & 1'h1;
  assign act_9234 = v_9235 | v_9284;
  assign v_9235 = v_9236 & 1'h1;
  assign v_9236 = v_9237 & v_9291;
  assign v_9237 = ~v_9238;
  assign v_9239 = v_9240 | v_9278;
  assign v_9240 = act_9241 & 1'h1;
  assign act_9241 = v_9242 | v_9255;
  assign v_9242 = v_9243 & 1'h1;
  assign v_9243 = v_9244 & v_9262;
  assign v_9244 = ~v_9245;
  assign v_9246 = v_9247 | v_9249;
  assign v_9247 = act_9248 & 1'h1;
  assign act_9248 = v_1744 | v_1738;
  assign v_9249 = v_9250 & 1'h1;
  assign v_9250 = v_9251 & v_9252;
  assign v_9251 = ~act_9248;
  assign v_9252 = v_9253 | v_9258;
  assign v_9253 = v_9254 | v_9256;
  assign v_9254 = mux_9254(v_9255);
  assign v_9255 = v_9245 & 1'h1;
  assign v_9256 = mux_9256(v_9257);
  assign v_9257 = ~v_9255;
  assign v_9258 = ~v_9245;
  assign v_9259 = v_9260 | v_9261;
  assign v_9260 = mux_9260(v_9247);
  assign v_9261 = mux_9261(v_9249);
  assign v_9263 = v_9264 | v_9266;
  assign v_9264 = act_9265 & 1'h1;
  assign act_9265 = v_1758 | v_1752;
  assign v_9266 = v_9267 & 1'h1;
  assign v_9267 = v_9268 & v_9269;
  assign v_9268 = ~act_9265;
  assign v_9269 = v_9270 | v_9274;
  assign v_9270 = v_9271 | v_9272;
  assign v_9271 = mux_9271(v_9242);
  assign v_9272 = mux_9272(v_9273);
  assign v_9273 = ~v_9242;
  assign v_9274 = ~v_9262;
  assign v_9275 = v_9276 | v_9277;
  assign v_9276 = mux_9276(v_9264);
  assign v_9277 = mux_9277(v_9266);
  assign v_9278 = v_9279 & 1'h1;
  assign v_9279 = v_9280 & v_9281;
  assign v_9280 = ~act_9241;
  assign v_9281 = v_9282 | v_9287;
  assign v_9282 = v_9283 | v_9285;
  assign v_9283 = mux_9283(v_9284);
  assign v_9284 = v_9238 & 1'h1;
  assign v_9285 = mux_9285(v_9286);
  assign v_9286 = ~v_9284;
  assign v_9287 = ~v_9238;
  assign v_9288 = v_9289 | v_9290;
  assign v_9289 = mux_9289(v_9240);
  assign v_9290 = mux_9290(v_9278);
  assign v_9292 = v_9293 | v_9331;
  assign v_9293 = act_9294 & 1'h1;
  assign act_9294 = v_9295 | v_9308;
  assign v_9295 = v_9296 & 1'h1;
  assign v_9296 = v_9297 & v_9315;
  assign v_9297 = ~v_9298;
  assign v_9299 = v_9300 | v_9302;
  assign v_9300 = act_9301 & 1'h1;
  assign act_9301 = v_1772 | v_1766;
  assign v_9302 = v_9303 & 1'h1;
  assign v_9303 = v_9304 & v_9305;
  assign v_9304 = ~act_9301;
  assign v_9305 = v_9306 | v_9311;
  assign v_9306 = v_9307 | v_9309;
  assign v_9307 = mux_9307(v_9308);
  assign v_9308 = v_9298 & 1'h1;
  assign v_9309 = mux_9309(v_9310);
  assign v_9310 = ~v_9308;
  assign v_9311 = ~v_9298;
  assign v_9312 = v_9313 | v_9314;
  assign v_9313 = mux_9313(v_9300);
  assign v_9314 = mux_9314(v_9302);
  assign v_9316 = v_9317 | v_9319;
  assign v_9317 = act_9318 & 1'h1;
  assign act_9318 = v_1786 | v_1780;
  assign v_9319 = v_9320 & 1'h1;
  assign v_9320 = v_9321 & v_9322;
  assign v_9321 = ~act_9318;
  assign v_9322 = v_9323 | v_9327;
  assign v_9323 = v_9324 | v_9325;
  assign v_9324 = mux_9324(v_9295);
  assign v_9325 = mux_9325(v_9326);
  assign v_9326 = ~v_9295;
  assign v_9327 = ~v_9315;
  assign v_9328 = v_9329 | v_9330;
  assign v_9329 = mux_9329(v_9317);
  assign v_9330 = mux_9330(v_9319);
  assign v_9331 = v_9332 & 1'h1;
  assign v_9332 = v_9333 & v_9334;
  assign v_9333 = ~act_9294;
  assign v_9334 = v_9335 | v_9339;
  assign v_9335 = v_9336 | v_9337;
  assign v_9336 = mux_9336(v_9235);
  assign v_9337 = mux_9337(v_9338);
  assign v_9338 = ~v_9235;
  assign v_9339 = ~v_9291;
  assign v_9340 = v_9341 | v_9342;
  assign v_9341 = mux_9341(v_9293);
  assign v_9342 = mux_9342(v_9331);
  assign v_9343 = v_9344 & 1'h1;
  assign v_9344 = v_9345 & v_9346;
  assign v_9345 = ~act_9234;
  assign v_9346 = v_9347 | v_9351;
  assign v_9347 = v_9348 | v_9349;
  assign v_9348 = mux_9348(v_9103);
  assign v_9349 = mux_9349(v_9350);
  assign v_9350 = ~v_9103;
  assign v_9351 = ~v_9231;
  assign v_9352 = v_9353 | v_9354;
  assign v_9353 = mux_9353(v_9233);
  assign v_9354 = mux_9354(v_9343);
  assign v_9355 = v_9356 & 1'h1;
  assign v_9356 = v_9357 & v_9358;
  assign v_9357 = ~act_9102;
  assign v_9358 = v_9359 | v_9363;
  assign v_9359 = v_9360 | v_9361;
  assign v_9360 = mux_9360(v_8827);
  assign v_9361 = mux_9361(v_9362);
  assign v_9362 = ~v_8827;
  assign v_9363 = ~v_9099;
  assign v_9364 = v_9365 | v_9366;
  assign v_9365 = mux_9365(v_9101);
  assign v_9366 = mux_9366(v_9355);
  assign v_9367 = v_9368 & 1'h1;
  assign v_9368 = v_9369 & v_9370;
  assign v_9369 = ~act_8826;
  assign v_9370 = v_9371 | v_9376;
  assign v_9371 = v_9372 | v_9374;
  assign v_9372 = mux_9372(v_9373);
  assign v_9373 = v_8823 & 1'h1;
  assign v_9374 = mux_9374(v_9375);
  assign v_9375 = ~v_9373;
  assign v_9376 = ~v_8823;
  assign v_9377 = v_9378 | v_9379;
  assign v_9378 = mux_9378(v_8825);
  assign v_9379 = mux_9379(v_9367);
  assign v_9381 = v_9382 | v_9924;
  assign v_9382 = act_9383 & 1'h1;
  assign act_9383 = v_9384 | v_9649;
  assign v_9384 = v_9385 & 1'h1;
  assign v_9385 = v_9386 & v_9656;
  assign v_9386 = ~v_9387;
  assign v_9388 = v_9389 | v_9643;
  assign v_9389 = act_9390 & 1'h1;
  assign act_9390 = v_9391 | v_9512;
  assign v_9391 = v_9392 & 1'h1;
  assign v_9392 = v_9393 & v_9519;
  assign v_9393 = ~v_9394;
  assign v_9395 = v_9396 | v_9506;
  assign v_9396 = act_9397 & 1'h1;
  assign act_9397 = v_9398 | v_9447;
  assign v_9398 = v_9399 & 1'h1;
  assign v_9399 = v_9400 & v_9454;
  assign v_9400 = ~v_9401;
  assign v_9402 = v_9403 | v_9441;
  assign v_9403 = act_9404 & 1'h1;
  assign act_9404 = v_9405 | v_9418;
  assign v_9405 = v_9406 & 1'h1;
  assign v_9406 = v_9407 & v_9425;
  assign v_9407 = ~v_9408;
  assign v_9409 = v_9410 | v_9412;
  assign v_9410 = act_9411 & 1'h1;
  assign act_9411 = v_1800 | v_1794;
  assign v_9412 = v_9413 & 1'h1;
  assign v_9413 = v_9414 & v_9415;
  assign v_9414 = ~act_9411;
  assign v_9415 = v_9416 | v_9421;
  assign v_9416 = v_9417 | v_9419;
  assign v_9417 = mux_9417(v_9418);
  assign v_9418 = v_9408 & 1'h1;
  assign v_9419 = mux_9419(v_9420);
  assign v_9420 = ~v_9418;
  assign v_9421 = ~v_9408;
  assign v_9422 = v_9423 | v_9424;
  assign v_9423 = mux_9423(v_9410);
  assign v_9424 = mux_9424(v_9412);
  assign v_9426 = v_9427 | v_9429;
  assign v_9427 = act_9428 & 1'h1;
  assign act_9428 = v_1814 | v_1808;
  assign v_9429 = v_9430 & 1'h1;
  assign v_9430 = v_9431 & v_9432;
  assign v_9431 = ~act_9428;
  assign v_9432 = v_9433 | v_9437;
  assign v_9433 = v_9434 | v_9435;
  assign v_9434 = mux_9434(v_9405);
  assign v_9435 = mux_9435(v_9436);
  assign v_9436 = ~v_9405;
  assign v_9437 = ~v_9425;
  assign v_9438 = v_9439 | v_9440;
  assign v_9439 = mux_9439(v_9427);
  assign v_9440 = mux_9440(v_9429);
  assign v_9441 = v_9442 & 1'h1;
  assign v_9442 = v_9443 & v_9444;
  assign v_9443 = ~act_9404;
  assign v_9444 = v_9445 | v_9450;
  assign v_9445 = v_9446 | v_9448;
  assign v_9446 = mux_9446(v_9447);
  assign v_9447 = v_9401 & 1'h1;
  assign v_9448 = mux_9448(v_9449);
  assign v_9449 = ~v_9447;
  assign v_9450 = ~v_9401;
  assign v_9451 = v_9452 | v_9453;
  assign v_9452 = mux_9452(v_9403);
  assign v_9453 = mux_9453(v_9441);
  assign v_9455 = v_9456 | v_9494;
  assign v_9456 = act_9457 & 1'h1;
  assign act_9457 = v_9458 | v_9471;
  assign v_9458 = v_9459 & 1'h1;
  assign v_9459 = v_9460 & v_9478;
  assign v_9460 = ~v_9461;
  assign v_9462 = v_9463 | v_9465;
  assign v_9463 = act_9464 & 1'h1;
  assign act_9464 = v_1828 | v_1822;
  assign v_9465 = v_9466 & 1'h1;
  assign v_9466 = v_9467 & v_9468;
  assign v_9467 = ~act_9464;
  assign v_9468 = v_9469 | v_9474;
  assign v_9469 = v_9470 | v_9472;
  assign v_9470 = mux_9470(v_9471);
  assign v_9471 = v_9461 & 1'h1;
  assign v_9472 = mux_9472(v_9473);
  assign v_9473 = ~v_9471;
  assign v_9474 = ~v_9461;
  assign v_9475 = v_9476 | v_9477;
  assign v_9476 = mux_9476(v_9463);
  assign v_9477 = mux_9477(v_9465);
  assign v_9479 = v_9480 | v_9482;
  assign v_9480 = act_9481 & 1'h1;
  assign act_9481 = v_1842 | v_1836;
  assign v_9482 = v_9483 & 1'h1;
  assign v_9483 = v_9484 & v_9485;
  assign v_9484 = ~act_9481;
  assign v_9485 = v_9486 | v_9490;
  assign v_9486 = v_9487 | v_9488;
  assign v_9487 = mux_9487(v_9458);
  assign v_9488 = mux_9488(v_9489);
  assign v_9489 = ~v_9458;
  assign v_9490 = ~v_9478;
  assign v_9491 = v_9492 | v_9493;
  assign v_9492 = mux_9492(v_9480);
  assign v_9493 = mux_9493(v_9482);
  assign v_9494 = v_9495 & 1'h1;
  assign v_9495 = v_9496 & v_9497;
  assign v_9496 = ~act_9457;
  assign v_9497 = v_9498 | v_9502;
  assign v_9498 = v_9499 | v_9500;
  assign v_9499 = mux_9499(v_9398);
  assign v_9500 = mux_9500(v_9501);
  assign v_9501 = ~v_9398;
  assign v_9502 = ~v_9454;
  assign v_9503 = v_9504 | v_9505;
  assign v_9504 = mux_9504(v_9456);
  assign v_9505 = mux_9505(v_9494);
  assign v_9506 = v_9507 & 1'h1;
  assign v_9507 = v_9508 & v_9509;
  assign v_9508 = ~act_9397;
  assign v_9509 = v_9510 | v_9515;
  assign v_9510 = v_9511 | v_9513;
  assign v_9511 = mux_9511(v_9512);
  assign v_9512 = v_9394 & 1'h1;
  assign v_9513 = mux_9513(v_9514);
  assign v_9514 = ~v_9512;
  assign v_9515 = ~v_9394;
  assign v_9516 = v_9517 | v_9518;
  assign v_9517 = mux_9517(v_9396);
  assign v_9518 = mux_9518(v_9506);
  assign v_9520 = v_9521 | v_9631;
  assign v_9521 = act_9522 & 1'h1;
  assign act_9522 = v_9523 | v_9572;
  assign v_9523 = v_9524 & 1'h1;
  assign v_9524 = v_9525 & v_9579;
  assign v_9525 = ~v_9526;
  assign v_9527 = v_9528 | v_9566;
  assign v_9528 = act_9529 & 1'h1;
  assign act_9529 = v_9530 | v_9543;
  assign v_9530 = v_9531 & 1'h1;
  assign v_9531 = v_9532 & v_9550;
  assign v_9532 = ~v_9533;
  assign v_9534 = v_9535 | v_9537;
  assign v_9535 = act_9536 & 1'h1;
  assign act_9536 = v_1856 | v_1850;
  assign v_9537 = v_9538 & 1'h1;
  assign v_9538 = v_9539 & v_9540;
  assign v_9539 = ~act_9536;
  assign v_9540 = v_9541 | v_9546;
  assign v_9541 = v_9542 | v_9544;
  assign v_9542 = mux_9542(v_9543);
  assign v_9543 = v_9533 & 1'h1;
  assign v_9544 = mux_9544(v_9545);
  assign v_9545 = ~v_9543;
  assign v_9546 = ~v_9533;
  assign v_9547 = v_9548 | v_9549;
  assign v_9548 = mux_9548(v_9535);
  assign v_9549 = mux_9549(v_9537);
  assign v_9551 = v_9552 | v_9554;
  assign v_9552 = act_9553 & 1'h1;
  assign act_9553 = v_1870 | v_1864;
  assign v_9554 = v_9555 & 1'h1;
  assign v_9555 = v_9556 & v_9557;
  assign v_9556 = ~act_9553;
  assign v_9557 = v_9558 | v_9562;
  assign v_9558 = v_9559 | v_9560;
  assign v_9559 = mux_9559(v_9530);
  assign v_9560 = mux_9560(v_9561);
  assign v_9561 = ~v_9530;
  assign v_9562 = ~v_9550;
  assign v_9563 = v_9564 | v_9565;
  assign v_9564 = mux_9564(v_9552);
  assign v_9565 = mux_9565(v_9554);
  assign v_9566 = v_9567 & 1'h1;
  assign v_9567 = v_9568 & v_9569;
  assign v_9568 = ~act_9529;
  assign v_9569 = v_9570 | v_9575;
  assign v_9570 = v_9571 | v_9573;
  assign v_9571 = mux_9571(v_9572);
  assign v_9572 = v_9526 & 1'h1;
  assign v_9573 = mux_9573(v_9574);
  assign v_9574 = ~v_9572;
  assign v_9575 = ~v_9526;
  assign v_9576 = v_9577 | v_9578;
  assign v_9577 = mux_9577(v_9528);
  assign v_9578 = mux_9578(v_9566);
  assign v_9580 = v_9581 | v_9619;
  assign v_9581 = act_9582 & 1'h1;
  assign act_9582 = v_9583 | v_9596;
  assign v_9583 = v_9584 & 1'h1;
  assign v_9584 = v_9585 & v_9603;
  assign v_9585 = ~v_9586;
  assign v_9587 = v_9588 | v_9590;
  assign v_9588 = act_9589 & 1'h1;
  assign act_9589 = v_1884 | v_1878;
  assign v_9590 = v_9591 & 1'h1;
  assign v_9591 = v_9592 & v_9593;
  assign v_9592 = ~act_9589;
  assign v_9593 = v_9594 | v_9599;
  assign v_9594 = v_9595 | v_9597;
  assign v_9595 = mux_9595(v_9596);
  assign v_9596 = v_9586 & 1'h1;
  assign v_9597 = mux_9597(v_9598);
  assign v_9598 = ~v_9596;
  assign v_9599 = ~v_9586;
  assign v_9600 = v_9601 | v_9602;
  assign v_9601 = mux_9601(v_9588);
  assign v_9602 = mux_9602(v_9590);
  assign v_9604 = v_9605 | v_9607;
  assign v_9605 = act_9606 & 1'h1;
  assign act_9606 = v_1898 | v_1892;
  assign v_9607 = v_9608 & 1'h1;
  assign v_9608 = v_9609 & v_9610;
  assign v_9609 = ~act_9606;
  assign v_9610 = v_9611 | v_9615;
  assign v_9611 = v_9612 | v_9613;
  assign v_9612 = mux_9612(v_9583);
  assign v_9613 = mux_9613(v_9614);
  assign v_9614 = ~v_9583;
  assign v_9615 = ~v_9603;
  assign v_9616 = v_9617 | v_9618;
  assign v_9617 = mux_9617(v_9605);
  assign v_9618 = mux_9618(v_9607);
  assign v_9619 = v_9620 & 1'h1;
  assign v_9620 = v_9621 & v_9622;
  assign v_9621 = ~act_9582;
  assign v_9622 = v_9623 | v_9627;
  assign v_9623 = v_9624 | v_9625;
  assign v_9624 = mux_9624(v_9523);
  assign v_9625 = mux_9625(v_9626);
  assign v_9626 = ~v_9523;
  assign v_9627 = ~v_9579;
  assign v_9628 = v_9629 | v_9630;
  assign v_9629 = mux_9629(v_9581);
  assign v_9630 = mux_9630(v_9619);
  assign v_9631 = v_9632 & 1'h1;
  assign v_9632 = v_9633 & v_9634;
  assign v_9633 = ~act_9522;
  assign v_9634 = v_9635 | v_9639;
  assign v_9635 = v_9636 | v_9637;
  assign v_9636 = mux_9636(v_9391);
  assign v_9637 = mux_9637(v_9638);
  assign v_9638 = ~v_9391;
  assign v_9639 = ~v_9519;
  assign v_9640 = v_9641 | v_9642;
  assign v_9641 = mux_9641(v_9521);
  assign v_9642 = mux_9642(v_9631);
  assign v_9643 = v_9644 & 1'h1;
  assign v_9644 = v_9645 & v_9646;
  assign v_9645 = ~act_9390;
  assign v_9646 = v_9647 | v_9652;
  assign v_9647 = v_9648 | v_9650;
  assign v_9648 = mux_9648(v_9649);
  assign v_9649 = v_9387 & 1'h1;
  assign v_9650 = mux_9650(v_9651);
  assign v_9651 = ~v_9649;
  assign v_9652 = ~v_9387;
  assign v_9653 = v_9654 | v_9655;
  assign v_9654 = mux_9654(v_9389);
  assign v_9655 = mux_9655(v_9643);
  assign v_9657 = v_9658 | v_9912;
  assign v_9658 = act_9659 & 1'h1;
  assign act_9659 = v_9660 | v_9781;
  assign v_9660 = v_9661 & 1'h1;
  assign v_9661 = v_9662 & v_9788;
  assign v_9662 = ~v_9663;
  assign v_9664 = v_9665 | v_9775;
  assign v_9665 = act_9666 & 1'h1;
  assign act_9666 = v_9667 | v_9716;
  assign v_9667 = v_9668 & 1'h1;
  assign v_9668 = v_9669 & v_9723;
  assign v_9669 = ~v_9670;
  assign v_9671 = v_9672 | v_9710;
  assign v_9672 = act_9673 & 1'h1;
  assign act_9673 = v_9674 | v_9687;
  assign v_9674 = v_9675 & 1'h1;
  assign v_9675 = v_9676 & v_9694;
  assign v_9676 = ~v_9677;
  assign v_9678 = v_9679 | v_9681;
  assign v_9679 = act_9680 & 1'h1;
  assign act_9680 = v_1912 | v_1906;
  assign v_9681 = v_9682 & 1'h1;
  assign v_9682 = v_9683 & v_9684;
  assign v_9683 = ~act_9680;
  assign v_9684 = v_9685 | v_9690;
  assign v_9685 = v_9686 | v_9688;
  assign v_9686 = mux_9686(v_9687);
  assign v_9687 = v_9677 & 1'h1;
  assign v_9688 = mux_9688(v_9689);
  assign v_9689 = ~v_9687;
  assign v_9690 = ~v_9677;
  assign v_9691 = v_9692 | v_9693;
  assign v_9692 = mux_9692(v_9679);
  assign v_9693 = mux_9693(v_9681);
  assign v_9695 = v_9696 | v_9698;
  assign v_9696 = act_9697 & 1'h1;
  assign act_9697 = v_1926 | v_1920;
  assign v_9698 = v_9699 & 1'h1;
  assign v_9699 = v_9700 & v_9701;
  assign v_9700 = ~act_9697;
  assign v_9701 = v_9702 | v_9706;
  assign v_9702 = v_9703 | v_9704;
  assign v_9703 = mux_9703(v_9674);
  assign v_9704 = mux_9704(v_9705);
  assign v_9705 = ~v_9674;
  assign v_9706 = ~v_9694;
  assign v_9707 = v_9708 | v_9709;
  assign v_9708 = mux_9708(v_9696);
  assign v_9709 = mux_9709(v_9698);
  assign v_9710 = v_9711 & 1'h1;
  assign v_9711 = v_9712 & v_9713;
  assign v_9712 = ~act_9673;
  assign v_9713 = v_9714 | v_9719;
  assign v_9714 = v_9715 | v_9717;
  assign v_9715 = mux_9715(v_9716);
  assign v_9716 = v_9670 & 1'h1;
  assign v_9717 = mux_9717(v_9718);
  assign v_9718 = ~v_9716;
  assign v_9719 = ~v_9670;
  assign v_9720 = v_9721 | v_9722;
  assign v_9721 = mux_9721(v_9672);
  assign v_9722 = mux_9722(v_9710);
  assign v_9724 = v_9725 | v_9763;
  assign v_9725 = act_9726 & 1'h1;
  assign act_9726 = v_9727 | v_9740;
  assign v_9727 = v_9728 & 1'h1;
  assign v_9728 = v_9729 & v_9747;
  assign v_9729 = ~v_9730;
  assign v_9731 = v_9732 | v_9734;
  assign v_9732 = act_9733 & 1'h1;
  assign act_9733 = v_1940 | v_1934;
  assign v_9734 = v_9735 & 1'h1;
  assign v_9735 = v_9736 & v_9737;
  assign v_9736 = ~act_9733;
  assign v_9737 = v_9738 | v_9743;
  assign v_9738 = v_9739 | v_9741;
  assign v_9739 = mux_9739(v_9740);
  assign v_9740 = v_9730 & 1'h1;
  assign v_9741 = mux_9741(v_9742);
  assign v_9742 = ~v_9740;
  assign v_9743 = ~v_9730;
  assign v_9744 = v_9745 | v_9746;
  assign v_9745 = mux_9745(v_9732);
  assign v_9746 = mux_9746(v_9734);
  assign v_9748 = v_9749 | v_9751;
  assign v_9749 = act_9750 & 1'h1;
  assign act_9750 = v_1954 | v_1948;
  assign v_9751 = v_9752 & 1'h1;
  assign v_9752 = v_9753 & v_9754;
  assign v_9753 = ~act_9750;
  assign v_9754 = v_9755 | v_9759;
  assign v_9755 = v_9756 | v_9757;
  assign v_9756 = mux_9756(v_9727);
  assign v_9757 = mux_9757(v_9758);
  assign v_9758 = ~v_9727;
  assign v_9759 = ~v_9747;
  assign v_9760 = v_9761 | v_9762;
  assign v_9761 = mux_9761(v_9749);
  assign v_9762 = mux_9762(v_9751);
  assign v_9763 = v_9764 & 1'h1;
  assign v_9764 = v_9765 & v_9766;
  assign v_9765 = ~act_9726;
  assign v_9766 = v_9767 | v_9771;
  assign v_9767 = v_9768 | v_9769;
  assign v_9768 = mux_9768(v_9667);
  assign v_9769 = mux_9769(v_9770);
  assign v_9770 = ~v_9667;
  assign v_9771 = ~v_9723;
  assign v_9772 = v_9773 | v_9774;
  assign v_9773 = mux_9773(v_9725);
  assign v_9774 = mux_9774(v_9763);
  assign v_9775 = v_9776 & 1'h1;
  assign v_9776 = v_9777 & v_9778;
  assign v_9777 = ~act_9666;
  assign v_9778 = v_9779 | v_9784;
  assign v_9779 = v_9780 | v_9782;
  assign v_9780 = mux_9780(v_9781);
  assign v_9781 = v_9663 & 1'h1;
  assign v_9782 = mux_9782(v_9783);
  assign v_9783 = ~v_9781;
  assign v_9784 = ~v_9663;
  assign v_9785 = v_9786 | v_9787;
  assign v_9786 = mux_9786(v_9665);
  assign v_9787 = mux_9787(v_9775);
  assign v_9789 = v_9790 | v_9900;
  assign v_9790 = act_9791 & 1'h1;
  assign act_9791 = v_9792 | v_9841;
  assign v_9792 = v_9793 & 1'h1;
  assign v_9793 = v_9794 & v_9848;
  assign v_9794 = ~v_9795;
  assign v_9796 = v_9797 | v_9835;
  assign v_9797 = act_9798 & 1'h1;
  assign act_9798 = v_9799 | v_9812;
  assign v_9799 = v_9800 & 1'h1;
  assign v_9800 = v_9801 & v_9819;
  assign v_9801 = ~v_9802;
  assign v_9803 = v_9804 | v_9806;
  assign v_9804 = act_9805 & 1'h1;
  assign act_9805 = v_1968 | v_1962;
  assign v_9806 = v_9807 & 1'h1;
  assign v_9807 = v_9808 & v_9809;
  assign v_9808 = ~act_9805;
  assign v_9809 = v_9810 | v_9815;
  assign v_9810 = v_9811 | v_9813;
  assign v_9811 = mux_9811(v_9812);
  assign v_9812 = v_9802 & 1'h1;
  assign v_9813 = mux_9813(v_9814);
  assign v_9814 = ~v_9812;
  assign v_9815 = ~v_9802;
  assign v_9816 = v_9817 | v_9818;
  assign v_9817 = mux_9817(v_9804);
  assign v_9818 = mux_9818(v_9806);
  assign v_9820 = v_9821 | v_9823;
  assign v_9821 = act_9822 & 1'h1;
  assign act_9822 = v_1982 | v_1976;
  assign v_9823 = v_9824 & 1'h1;
  assign v_9824 = v_9825 & v_9826;
  assign v_9825 = ~act_9822;
  assign v_9826 = v_9827 | v_9831;
  assign v_9827 = v_9828 | v_9829;
  assign v_9828 = mux_9828(v_9799);
  assign v_9829 = mux_9829(v_9830);
  assign v_9830 = ~v_9799;
  assign v_9831 = ~v_9819;
  assign v_9832 = v_9833 | v_9834;
  assign v_9833 = mux_9833(v_9821);
  assign v_9834 = mux_9834(v_9823);
  assign v_9835 = v_9836 & 1'h1;
  assign v_9836 = v_9837 & v_9838;
  assign v_9837 = ~act_9798;
  assign v_9838 = v_9839 | v_9844;
  assign v_9839 = v_9840 | v_9842;
  assign v_9840 = mux_9840(v_9841);
  assign v_9841 = v_9795 & 1'h1;
  assign v_9842 = mux_9842(v_9843);
  assign v_9843 = ~v_9841;
  assign v_9844 = ~v_9795;
  assign v_9845 = v_9846 | v_9847;
  assign v_9846 = mux_9846(v_9797);
  assign v_9847 = mux_9847(v_9835);
  assign v_9849 = v_9850 | v_9888;
  assign v_9850 = act_9851 & 1'h1;
  assign act_9851 = v_9852 | v_9865;
  assign v_9852 = v_9853 & 1'h1;
  assign v_9853 = v_9854 & v_9872;
  assign v_9854 = ~v_9855;
  assign v_9856 = v_9857 | v_9859;
  assign v_9857 = act_9858 & 1'h1;
  assign act_9858 = v_1996 | v_1990;
  assign v_9859 = v_9860 & 1'h1;
  assign v_9860 = v_9861 & v_9862;
  assign v_9861 = ~act_9858;
  assign v_9862 = v_9863 | v_9868;
  assign v_9863 = v_9864 | v_9866;
  assign v_9864 = mux_9864(v_9865);
  assign v_9865 = v_9855 & 1'h1;
  assign v_9866 = mux_9866(v_9867);
  assign v_9867 = ~v_9865;
  assign v_9868 = ~v_9855;
  assign v_9869 = v_9870 | v_9871;
  assign v_9870 = mux_9870(v_9857);
  assign v_9871 = mux_9871(v_9859);
  assign v_9873 = v_9874 | v_9876;
  assign v_9874 = act_9875 & 1'h1;
  assign act_9875 = v_2010 | v_2004;
  assign v_9876 = v_9877 & 1'h1;
  assign v_9877 = v_9878 & v_9879;
  assign v_9878 = ~act_9875;
  assign v_9879 = v_9880 | v_9884;
  assign v_9880 = v_9881 | v_9882;
  assign v_9881 = mux_9881(v_9852);
  assign v_9882 = mux_9882(v_9883);
  assign v_9883 = ~v_9852;
  assign v_9884 = ~v_9872;
  assign v_9885 = v_9886 | v_9887;
  assign v_9886 = mux_9886(v_9874);
  assign v_9887 = mux_9887(v_9876);
  assign v_9888 = v_9889 & 1'h1;
  assign v_9889 = v_9890 & v_9891;
  assign v_9890 = ~act_9851;
  assign v_9891 = v_9892 | v_9896;
  assign v_9892 = v_9893 | v_9894;
  assign v_9893 = mux_9893(v_9792);
  assign v_9894 = mux_9894(v_9895);
  assign v_9895 = ~v_9792;
  assign v_9896 = ~v_9848;
  assign v_9897 = v_9898 | v_9899;
  assign v_9898 = mux_9898(v_9850);
  assign v_9899 = mux_9899(v_9888);
  assign v_9900 = v_9901 & 1'h1;
  assign v_9901 = v_9902 & v_9903;
  assign v_9902 = ~act_9791;
  assign v_9903 = v_9904 | v_9908;
  assign v_9904 = v_9905 | v_9906;
  assign v_9905 = mux_9905(v_9660);
  assign v_9906 = mux_9906(v_9907);
  assign v_9907 = ~v_9660;
  assign v_9908 = ~v_9788;
  assign v_9909 = v_9910 | v_9911;
  assign v_9910 = mux_9910(v_9790);
  assign v_9911 = mux_9911(v_9900);
  assign v_9912 = v_9913 & 1'h1;
  assign v_9913 = v_9914 & v_9915;
  assign v_9914 = ~act_9659;
  assign v_9915 = v_9916 | v_9920;
  assign v_9916 = v_9917 | v_9918;
  assign v_9917 = mux_9917(v_9384);
  assign v_9918 = mux_9918(v_9919);
  assign v_9919 = ~v_9384;
  assign v_9920 = ~v_9656;
  assign v_9921 = v_9922 | v_9923;
  assign v_9922 = mux_9922(v_9658);
  assign v_9923 = mux_9923(v_9912);
  assign v_9924 = v_9925 & 1'h1;
  assign v_9925 = v_9926 & v_9927;
  assign v_9926 = ~act_9383;
  assign v_9927 = v_9928 | v_9932;
  assign v_9928 = v_9929 | v_9930;
  assign v_9929 = mux_9929(v_8820);
  assign v_9930 = mux_9930(v_9931);
  assign v_9931 = ~v_8820;
  assign v_9932 = ~v_9380;
  assign v_9933 = v_9934 | v_9935;
  assign v_9934 = mux_9934(v_9382);
  assign v_9935 = mux_9935(v_9924);
  assign v_9936 = v_9937 & 1'h1;
  assign v_9937 = v_9938 & v_9939;
  assign v_9938 = ~act_8819;
  assign v_9939 = v_9940 | v_9944;
  assign v_9940 = v_9941 | v_9942;
  assign v_9941 = mux_9941(v_7680);
  assign v_9942 = mux_9942(v_9943);
  assign v_9943 = ~v_7680;
  assign v_9944 = ~v_8816;
  assign v_9945 = v_9946 | v_9947;
  assign v_9946 = mux_9946(v_8818);
  assign v_9947 = mux_9947(v_9936);
  assign v_9948 = v_9949 & 1'h1;
  assign v_9949 = v_9950 & v_9951;
  assign v_9950 = ~act_7679;
  assign v_9951 = v_9952 | v_9956;
  assign v_9952 = v_9953 | v_9954;
  assign v_9953 = mux_9953(v_5388);
  assign v_9954 = mux_9954(v_9955);
  assign v_9955 = ~v_5388;
  assign v_9956 = ~v_7676;
  assign v_9957 = v_9958 | v_9959;
  assign v_9958 = mux_9958(v_7678);
  assign v_9959 = mux_9959(v_9948);
  assign v_9960 = v_9961 & 1'h1;
  assign v_9961 = v_9962 & v_9963;
  assign v_9962 = ~act_5387;
  assign v_9963 = v_9964 | v_9968;
  assign v_9964 = v_9965 | v_9966;
  assign v_9965 = mux_9965(v_2808);
  assign v_9966 = mux_9966(v_9967);
  assign v_9967 = ~v_2808;
  assign v_9968 = ~v_5384;
  assign v_9969 = v_9970 | v_9971;
  assign v_9970 = mux_9970(v_5386);
  assign v_9971 = mux_9971(v_9960);
  assign v_9972 = v_9973 & 1'h1;
  assign v_9973 = v_9974 & v_9975;
  assign v_9974 = ~act_2807;
  assign v_9975 = v_9976 | v_9982;
  assign v_9976 = v_9977 | v_9980;
  assign v_9977 = mux_9977(v_9978);
  assign v_9978 = v_9979 & 1'h1;
  assign v_9979 = out_consume_en;
  assign v_9980 = mux_9980(v_9981);
  assign v_9981 = ~v_9978;
  assign v_9982 = ~v_2804;
  assign v_9983 = v_9984 | v_9985;
  assign v_9984 = mux_9984(v_2806);
  assign v_9985 = mux_9985(v_9972);
  assign out_peek = v_9987;
  assign v_9988 = v_9989 | v_9991;
  assign v_9989 = mux_9989(v_9990);
  assign v_9990 = ~act_2807;
  assign v_9991 = v_9992 | v_11778;
  assign v_9992 = mux_9992(v_2808);
  assign v_9994 = v_9995 | v_9997;
  assign v_9995 = mux_9995(v_9996);
  assign v_9996 = ~act_5387;
  assign v_9997 = v_9998 | v_10888;
  assign v_9998 = mux_9998(v_5388);
  assign v_10000 = v_10001 | v_10003;
  assign v_10001 = mux_10001(v_10002);
  assign v_10002 = ~act_7679;
  assign v_10003 = v_10004 | v_10446;
  assign v_10004 = mux_10004(v_7680);
  assign v_10006 = v_10007 | v_10009;
  assign v_10007 = mux_10007(v_10008);
  assign v_10008 = ~act_8819;
  assign v_10009 = v_10010 | v_10228;
  assign v_10010 = mux_10010(v_8820);
  assign v_10012 = v_10013 | v_10015;
  assign v_10013 = mux_10013(v_10014);
  assign v_10014 = ~act_9383;
  assign v_10015 = v_10016 | v_10122;
  assign v_10016 = mux_10016(v_9384);
  assign v_10018 = v_10019 | v_10021;
  assign v_10019 = mux_10019(v_10020);
  assign v_10020 = ~act_9659;
  assign v_10021 = v_10022 | v_10072;
  assign v_10022 = mux_10022(v_9660);
  assign v_10024 = v_10025 | v_10027;
  assign v_10025 = mux_10025(v_10026);
  assign v_10026 = ~act_9791;
  assign v_10027 = v_10028 | v_10050;
  assign v_10028 = mux_10028(v_9792);
  assign v_10030 = v_10031 | v_10033;
  assign v_10031 = mux_10031(v_10032);
  assign v_10032 = ~act_9851;
  assign v_10033 = v_10034 | v_10042;
  assign v_10034 = mux_10034(v_9852);
  assign v_10036 = v_10037 | v_10039;
  assign v_10037 = mux_10037(v_10038);
  assign v_10038 = ~act_9875;
  assign v_10039 = v_10040 | v_10041;
  assign v_10040 = mux_10040(v_2010);
  assign v_10041 = mux_10041(v_2004);
  assign v_10042 = mux_10042(v_9865);
  assign v_10044 = v_10045 | v_10047;
  assign v_10045 = mux_10045(v_10046);
  assign v_10046 = ~act_9858;
  assign v_10047 = v_10048 | v_10049;
  assign v_10048 = mux_10048(v_1996);
  assign v_10049 = mux_10049(v_1990);
  assign v_10050 = mux_10050(v_9841);
  assign v_10052 = v_10053 | v_10055;
  assign v_10053 = mux_10053(v_10054);
  assign v_10054 = ~act_9798;
  assign v_10055 = v_10056 | v_10064;
  assign v_10056 = mux_10056(v_9799);
  assign v_10058 = v_10059 | v_10061;
  assign v_10059 = mux_10059(v_10060);
  assign v_10060 = ~act_9822;
  assign v_10061 = v_10062 | v_10063;
  assign v_10062 = mux_10062(v_1982);
  assign v_10063 = mux_10063(v_1976);
  assign v_10064 = mux_10064(v_9812);
  assign v_10066 = v_10067 | v_10069;
  assign v_10067 = mux_10067(v_10068);
  assign v_10068 = ~act_9805;
  assign v_10069 = v_10070 | v_10071;
  assign v_10070 = mux_10070(v_1968);
  assign v_10071 = mux_10071(v_1962);
  assign v_10072 = mux_10072(v_9781);
  assign v_10074 = v_10075 | v_10077;
  assign v_10075 = mux_10075(v_10076);
  assign v_10076 = ~act_9666;
  assign v_10077 = v_10078 | v_10100;
  assign v_10078 = mux_10078(v_9667);
  assign v_10080 = v_10081 | v_10083;
  assign v_10081 = mux_10081(v_10082);
  assign v_10082 = ~act_9726;
  assign v_10083 = v_10084 | v_10092;
  assign v_10084 = mux_10084(v_9727);
  assign v_10086 = v_10087 | v_10089;
  assign v_10087 = mux_10087(v_10088);
  assign v_10088 = ~act_9750;
  assign v_10089 = v_10090 | v_10091;
  assign v_10090 = mux_10090(v_1954);
  assign v_10091 = mux_10091(v_1948);
  assign v_10092 = mux_10092(v_9740);
  assign v_10094 = v_10095 | v_10097;
  assign v_10095 = mux_10095(v_10096);
  assign v_10096 = ~act_9733;
  assign v_10097 = v_10098 | v_10099;
  assign v_10098 = mux_10098(v_1940);
  assign v_10099 = mux_10099(v_1934);
  assign v_10100 = mux_10100(v_9716);
  assign v_10102 = v_10103 | v_10105;
  assign v_10103 = mux_10103(v_10104);
  assign v_10104 = ~act_9673;
  assign v_10105 = v_10106 | v_10114;
  assign v_10106 = mux_10106(v_9674);
  assign v_10108 = v_10109 | v_10111;
  assign v_10109 = mux_10109(v_10110);
  assign v_10110 = ~act_9697;
  assign v_10111 = v_10112 | v_10113;
  assign v_10112 = mux_10112(v_1926);
  assign v_10113 = mux_10113(v_1920);
  assign v_10114 = mux_10114(v_9687);
  assign v_10116 = v_10117 | v_10119;
  assign v_10117 = mux_10117(v_10118);
  assign v_10118 = ~act_9680;
  assign v_10119 = v_10120 | v_10121;
  assign v_10120 = mux_10120(v_1912);
  assign v_10121 = mux_10121(v_1906);
  assign v_10122 = mux_10122(v_9649);
  assign v_10124 = v_10125 | v_10127;
  assign v_10125 = mux_10125(v_10126);
  assign v_10126 = ~act_9390;
  assign v_10127 = v_10128 | v_10178;
  assign v_10128 = mux_10128(v_9391);
  assign v_10130 = v_10131 | v_10133;
  assign v_10131 = mux_10131(v_10132);
  assign v_10132 = ~act_9522;
  assign v_10133 = v_10134 | v_10156;
  assign v_10134 = mux_10134(v_9523);
  assign v_10136 = v_10137 | v_10139;
  assign v_10137 = mux_10137(v_10138);
  assign v_10138 = ~act_9582;
  assign v_10139 = v_10140 | v_10148;
  assign v_10140 = mux_10140(v_9583);
  assign v_10142 = v_10143 | v_10145;
  assign v_10143 = mux_10143(v_10144);
  assign v_10144 = ~act_9606;
  assign v_10145 = v_10146 | v_10147;
  assign v_10146 = mux_10146(v_1898);
  assign v_10147 = mux_10147(v_1892);
  assign v_10148 = mux_10148(v_9596);
  assign v_10150 = v_10151 | v_10153;
  assign v_10151 = mux_10151(v_10152);
  assign v_10152 = ~act_9589;
  assign v_10153 = v_10154 | v_10155;
  assign v_10154 = mux_10154(v_1884);
  assign v_10155 = mux_10155(v_1878);
  assign v_10156 = mux_10156(v_9572);
  assign v_10158 = v_10159 | v_10161;
  assign v_10159 = mux_10159(v_10160);
  assign v_10160 = ~act_9529;
  assign v_10161 = v_10162 | v_10170;
  assign v_10162 = mux_10162(v_9530);
  assign v_10164 = v_10165 | v_10167;
  assign v_10165 = mux_10165(v_10166);
  assign v_10166 = ~act_9553;
  assign v_10167 = v_10168 | v_10169;
  assign v_10168 = mux_10168(v_1870);
  assign v_10169 = mux_10169(v_1864);
  assign v_10170 = mux_10170(v_9543);
  assign v_10172 = v_10173 | v_10175;
  assign v_10173 = mux_10173(v_10174);
  assign v_10174 = ~act_9536;
  assign v_10175 = v_10176 | v_10177;
  assign v_10176 = mux_10176(v_1856);
  assign v_10177 = mux_10177(v_1850);
  assign v_10178 = mux_10178(v_9512);
  assign v_10180 = v_10181 | v_10183;
  assign v_10181 = mux_10181(v_10182);
  assign v_10182 = ~act_9397;
  assign v_10183 = v_10184 | v_10206;
  assign v_10184 = mux_10184(v_9398);
  assign v_10186 = v_10187 | v_10189;
  assign v_10187 = mux_10187(v_10188);
  assign v_10188 = ~act_9457;
  assign v_10189 = v_10190 | v_10198;
  assign v_10190 = mux_10190(v_9458);
  assign v_10192 = v_10193 | v_10195;
  assign v_10193 = mux_10193(v_10194);
  assign v_10194 = ~act_9481;
  assign v_10195 = v_10196 | v_10197;
  assign v_10196 = mux_10196(v_1842);
  assign v_10197 = mux_10197(v_1836);
  assign v_10198 = mux_10198(v_9471);
  assign v_10200 = v_10201 | v_10203;
  assign v_10201 = mux_10201(v_10202);
  assign v_10202 = ~act_9464;
  assign v_10203 = v_10204 | v_10205;
  assign v_10204 = mux_10204(v_1828);
  assign v_10205 = mux_10205(v_1822);
  assign v_10206 = mux_10206(v_9447);
  assign v_10208 = v_10209 | v_10211;
  assign v_10209 = mux_10209(v_10210);
  assign v_10210 = ~act_9404;
  assign v_10211 = v_10212 | v_10220;
  assign v_10212 = mux_10212(v_9405);
  assign v_10214 = v_10215 | v_10217;
  assign v_10215 = mux_10215(v_10216);
  assign v_10216 = ~act_9428;
  assign v_10217 = v_10218 | v_10219;
  assign v_10218 = mux_10218(v_1814);
  assign v_10219 = mux_10219(v_1808);
  assign v_10220 = mux_10220(v_9418);
  assign v_10222 = v_10223 | v_10225;
  assign v_10223 = mux_10223(v_10224);
  assign v_10224 = ~act_9411;
  assign v_10225 = v_10226 | v_10227;
  assign v_10226 = mux_10226(v_1800);
  assign v_10227 = mux_10227(v_1794);
  assign v_10228 = mux_10228(v_9373);
  assign v_10230 = v_10231 | v_10233;
  assign v_10231 = mux_10231(v_10232);
  assign v_10232 = ~act_8826;
  assign v_10233 = v_10234 | v_10340;
  assign v_10234 = mux_10234(v_8827);
  assign v_10236 = v_10237 | v_10239;
  assign v_10237 = mux_10237(v_10238);
  assign v_10238 = ~act_9102;
  assign v_10239 = v_10240 | v_10290;
  assign v_10240 = mux_10240(v_9103);
  assign v_10242 = v_10243 | v_10245;
  assign v_10243 = mux_10243(v_10244);
  assign v_10244 = ~act_9234;
  assign v_10245 = v_10246 | v_10268;
  assign v_10246 = mux_10246(v_9235);
  assign v_10248 = v_10249 | v_10251;
  assign v_10249 = mux_10249(v_10250);
  assign v_10250 = ~act_9294;
  assign v_10251 = v_10252 | v_10260;
  assign v_10252 = mux_10252(v_9295);
  assign v_10254 = v_10255 | v_10257;
  assign v_10255 = mux_10255(v_10256);
  assign v_10256 = ~act_9318;
  assign v_10257 = v_10258 | v_10259;
  assign v_10258 = mux_10258(v_1786);
  assign v_10259 = mux_10259(v_1780);
  assign v_10260 = mux_10260(v_9308);
  assign v_10262 = v_10263 | v_10265;
  assign v_10263 = mux_10263(v_10264);
  assign v_10264 = ~act_9301;
  assign v_10265 = v_10266 | v_10267;
  assign v_10266 = mux_10266(v_1772);
  assign v_10267 = mux_10267(v_1766);
  assign v_10268 = mux_10268(v_9284);
  assign v_10270 = v_10271 | v_10273;
  assign v_10271 = mux_10271(v_10272);
  assign v_10272 = ~act_9241;
  assign v_10273 = v_10274 | v_10282;
  assign v_10274 = mux_10274(v_9242);
  assign v_10276 = v_10277 | v_10279;
  assign v_10277 = mux_10277(v_10278);
  assign v_10278 = ~act_9265;
  assign v_10279 = v_10280 | v_10281;
  assign v_10280 = mux_10280(v_1758);
  assign v_10281 = mux_10281(v_1752);
  assign v_10282 = mux_10282(v_9255);
  assign v_10284 = v_10285 | v_10287;
  assign v_10285 = mux_10285(v_10286);
  assign v_10286 = ~act_9248;
  assign v_10287 = v_10288 | v_10289;
  assign v_10288 = mux_10288(v_1744);
  assign v_10289 = mux_10289(v_1738);
  assign v_10290 = mux_10290(v_9224);
  assign v_10292 = v_10293 | v_10295;
  assign v_10293 = mux_10293(v_10294);
  assign v_10294 = ~act_9109;
  assign v_10295 = v_10296 | v_10318;
  assign v_10296 = mux_10296(v_9110);
  assign v_10298 = v_10299 | v_10301;
  assign v_10299 = mux_10299(v_10300);
  assign v_10300 = ~act_9169;
  assign v_10301 = v_10302 | v_10310;
  assign v_10302 = mux_10302(v_9170);
  assign v_10304 = v_10305 | v_10307;
  assign v_10305 = mux_10305(v_10306);
  assign v_10306 = ~act_9193;
  assign v_10307 = v_10308 | v_10309;
  assign v_10308 = mux_10308(v_1730);
  assign v_10309 = mux_10309(v_1724);
  assign v_10310 = mux_10310(v_9183);
  assign v_10312 = v_10313 | v_10315;
  assign v_10313 = mux_10313(v_10314);
  assign v_10314 = ~act_9176;
  assign v_10315 = v_10316 | v_10317;
  assign v_10316 = mux_10316(v_1716);
  assign v_10317 = mux_10317(v_1710);
  assign v_10318 = mux_10318(v_9159);
  assign v_10320 = v_10321 | v_10323;
  assign v_10321 = mux_10321(v_10322);
  assign v_10322 = ~act_9116;
  assign v_10323 = v_10324 | v_10332;
  assign v_10324 = mux_10324(v_9117);
  assign v_10326 = v_10327 | v_10329;
  assign v_10327 = mux_10327(v_10328);
  assign v_10328 = ~act_9140;
  assign v_10329 = v_10330 | v_10331;
  assign v_10330 = mux_10330(v_1702);
  assign v_10331 = mux_10331(v_1696);
  assign v_10332 = mux_10332(v_9130);
  assign v_10334 = v_10335 | v_10337;
  assign v_10335 = mux_10335(v_10336);
  assign v_10336 = ~act_9123;
  assign v_10337 = v_10338 | v_10339;
  assign v_10338 = mux_10338(v_1688);
  assign v_10339 = mux_10339(v_1682);
  assign v_10340 = mux_10340(v_9092);
  assign v_10342 = v_10343 | v_10345;
  assign v_10343 = mux_10343(v_10344);
  assign v_10344 = ~act_8833;
  assign v_10345 = v_10346 | v_10396;
  assign v_10346 = mux_10346(v_8834);
  assign v_10348 = v_10349 | v_10351;
  assign v_10349 = mux_10349(v_10350);
  assign v_10350 = ~act_8965;
  assign v_10351 = v_10352 | v_10374;
  assign v_10352 = mux_10352(v_8966);
  assign v_10354 = v_10355 | v_10357;
  assign v_10355 = mux_10355(v_10356);
  assign v_10356 = ~act_9025;
  assign v_10357 = v_10358 | v_10366;
  assign v_10358 = mux_10358(v_9026);
  assign v_10360 = v_10361 | v_10363;
  assign v_10361 = mux_10361(v_10362);
  assign v_10362 = ~act_9049;
  assign v_10363 = v_10364 | v_10365;
  assign v_10364 = mux_10364(v_1674);
  assign v_10365 = mux_10365(v_1668);
  assign v_10366 = mux_10366(v_9039);
  assign v_10368 = v_10369 | v_10371;
  assign v_10369 = mux_10369(v_10370);
  assign v_10370 = ~act_9032;
  assign v_10371 = v_10372 | v_10373;
  assign v_10372 = mux_10372(v_1660);
  assign v_10373 = mux_10373(v_1654);
  assign v_10374 = mux_10374(v_9015);
  assign v_10376 = v_10377 | v_10379;
  assign v_10377 = mux_10377(v_10378);
  assign v_10378 = ~act_8972;
  assign v_10379 = v_10380 | v_10388;
  assign v_10380 = mux_10380(v_8973);
  assign v_10382 = v_10383 | v_10385;
  assign v_10383 = mux_10383(v_10384);
  assign v_10384 = ~act_8996;
  assign v_10385 = v_10386 | v_10387;
  assign v_10386 = mux_10386(v_1646);
  assign v_10387 = mux_10387(v_1640);
  assign v_10388 = mux_10388(v_8986);
  assign v_10390 = v_10391 | v_10393;
  assign v_10391 = mux_10391(v_10392);
  assign v_10392 = ~act_8979;
  assign v_10393 = v_10394 | v_10395;
  assign v_10394 = mux_10394(v_1632);
  assign v_10395 = mux_10395(v_1626);
  assign v_10396 = mux_10396(v_8955);
  assign v_10398 = v_10399 | v_10401;
  assign v_10399 = mux_10399(v_10400);
  assign v_10400 = ~act_8840;
  assign v_10401 = v_10402 | v_10424;
  assign v_10402 = mux_10402(v_8841);
  assign v_10404 = v_10405 | v_10407;
  assign v_10405 = mux_10405(v_10406);
  assign v_10406 = ~act_8900;
  assign v_10407 = v_10408 | v_10416;
  assign v_10408 = mux_10408(v_8901);
  assign v_10410 = v_10411 | v_10413;
  assign v_10411 = mux_10411(v_10412);
  assign v_10412 = ~act_8924;
  assign v_10413 = v_10414 | v_10415;
  assign v_10414 = mux_10414(v_1618);
  assign v_10415 = mux_10415(v_1612);
  assign v_10416 = mux_10416(v_8914);
  assign v_10418 = v_10419 | v_10421;
  assign v_10419 = mux_10419(v_10420);
  assign v_10420 = ~act_8907;
  assign v_10421 = v_10422 | v_10423;
  assign v_10422 = mux_10422(v_1604);
  assign v_10423 = mux_10423(v_1598);
  assign v_10424 = mux_10424(v_8890);
  assign v_10426 = v_10427 | v_10429;
  assign v_10427 = mux_10427(v_10428);
  assign v_10428 = ~act_8847;
  assign v_10429 = v_10430 | v_10438;
  assign v_10430 = mux_10430(v_8848);
  assign v_10432 = v_10433 | v_10435;
  assign v_10433 = mux_10433(v_10434);
  assign v_10434 = ~act_8871;
  assign v_10435 = v_10436 | v_10437;
  assign v_10436 = mux_10436(v_1590);
  assign v_10437 = mux_10437(v_1584);
  assign v_10438 = mux_10438(v_8861);
  assign v_10440 = v_10441 | v_10443;
  assign v_10441 = mux_10441(v_10442);
  assign v_10442 = ~act_8854;
  assign v_10443 = v_10444 | v_10445;
  assign v_10444 = mux_10444(v_1576);
  assign v_10445 = mux_10445(v_1570);
  assign v_10446 = mux_10446(v_8809);
  assign v_10448 = v_10449 | v_10451;
  assign v_10449 = mux_10449(v_10450);
  assign v_10450 = ~act_7686;
  assign v_10451 = v_10452 | v_10670;
  assign v_10452 = mux_10452(v_7687);
  assign v_10454 = v_10455 | v_10457;
  assign v_10455 = mux_10455(v_10456);
  assign v_10456 = ~act_8250;
  assign v_10457 = v_10458 | v_10564;
  assign v_10458 = mux_10458(v_8251);
  assign v_10460 = v_10461 | v_10463;
  assign v_10461 = mux_10461(v_10462);
  assign v_10462 = ~act_8526;
  assign v_10463 = v_10464 | v_10514;
  assign v_10464 = mux_10464(v_8527);
  assign v_10466 = v_10467 | v_10469;
  assign v_10467 = mux_10467(v_10468);
  assign v_10468 = ~act_8658;
  assign v_10469 = v_10470 | v_10492;
  assign v_10470 = mux_10470(v_8659);
  assign v_10472 = v_10473 | v_10475;
  assign v_10473 = mux_10473(v_10474);
  assign v_10474 = ~act_8718;
  assign v_10475 = v_10476 | v_10484;
  assign v_10476 = mux_10476(v_8719);
  assign v_10478 = v_10479 | v_10481;
  assign v_10479 = mux_10479(v_10480);
  assign v_10480 = ~act_8742;
  assign v_10481 = v_10482 | v_10483;
  assign v_10482 = mux_10482(v_1562);
  assign v_10483 = mux_10483(v_1556);
  assign v_10484 = mux_10484(v_8732);
  assign v_10486 = v_10487 | v_10489;
  assign v_10487 = mux_10487(v_10488);
  assign v_10488 = ~act_8725;
  assign v_10489 = v_10490 | v_10491;
  assign v_10490 = mux_10490(v_1548);
  assign v_10491 = mux_10491(v_1542);
  assign v_10492 = mux_10492(v_8708);
  assign v_10494 = v_10495 | v_10497;
  assign v_10495 = mux_10495(v_10496);
  assign v_10496 = ~act_8665;
  assign v_10497 = v_10498 | v_10506;
  assign v_10498 = mux_10498(v_8666);
  assign v_10500 = v_10501 | v_10503;
  assign v_10501 = mux_10501(v_10502);
  assign v_10502 = ~act_8689;
  assign v_10503 = v_10504 | v_10505;
  assign v_10504 = mux_10504(v_1534);
  assign v_10505 = mux_10505(v_1528);
  assign v_10506 = mux_10506(v_8679);
  assign v_10508 = v_10509 | v_10511;
  assign v_10509 = mux_10509(v_10510);
  assign v_10510 = ~act_8672;
  assign v_10511 = v_10512 | v_10513;
  assign v_10512 = mux_10512(v_1520);
  assign v_10513 = mux_10513(v_1514);
  assign v_10514 = mux_10514(v_8648);
  assign v_10516 = v_10517 | v_10519;
  assign v_10517 = mux_10517(v_10518);
  assign v_10518 = ~act_8533;
  assign v_10519 = v_10520 | v_10542;
  assign v_10520 = mux_10520(v_8534);
  assign v_10522 = v_10523 | v_10525;
  assign v_10523 = mux_10523(v_10524);
  assign v_10524 = ~act_8593;
  assign v_10525 = v_10526 | v_10534;
  assign v_10526 = mux_10526(v_8594);
  assign v_10528 = v_10529 | v_10531;
  assign v_10529 = mux_10529(v_10530);
  assign v_10530 = ~act_8617;
  assign v_10531 = v_10532 | v_10533;
  assign v_10532 = mux_10532(v_1506);
  assign v_10533 = mux_10533(v_1500);
  assign v_10534 = mux_10534(v_8607);
  assign v_10536 = v_10537 | v_10539;
  assign v_10537 = mux_10537(v_10538);
  assign v_10538 = ~act_8600;
  assign v_10539 = v_10540 | v_10541;
  assign v_10540 = mux_10540(v_1492);
  assign v_10541 = mux_10541(v_1486);
  assign v_10542 = mux_10542(v_8583);
  assign v_10544 = v_10545 | v_10547;
  assign v_10545 = mux_10545(v_10546);
  assign v_10546 = ~act_8540;
  assign v_10547 = v_10548 | v_10556;
  assign v_10548 = mux_10548(v_8541);
  assign v_10550 = v_10551 | v_10553;
  assign v_10551 = mux_10551(v_10552);
  assign v_10552 = ~act_8564;
  assign v_10553 = v_10554 | v_10555;
  assign v_10554 = mux_10554(v_1478);
  assign v_10555 = mux_10555(v_1472);
  assign v_10556 = mux_10556(v_8554);
  assign v_10558 = v_10559 | v_10561;
  assign v_10559 = mux_10559(v_10560);
  assign v_10560 = ~act_8547;
  assign v_10561 = v_10562 | v_10563;
  assign v_10562 = mux_10562(v_1464);
  assign v_10563 = mux_10563(v_1458);
  assign v_10564 = mux_10564(v_8516);
  assign v_10566 = v_10567 | v_10569;
  assign v_10567 = mux_10567(v_10568);
  assign v_10568 = ~act_8257;
  assign v_10569 = v_10570 | v_10620;
  assign v_10570 = mux_10570(v_8258);
  assign v_10572 = v_10573 | v_10575;
  assign v_10573 = mux_10573(v_10574);
  assign v_10574 = ~act_8389;
  assign v_10575 = v_10576 | v_10598;
  assign v_10576 = mux_10576(v_8390);
  assign v_10578 = v_10579 | v_10581;
  assign v_10579 = mux_10579(v_10580);
  assign v_10580 = ~act_8449;
  assign v_10581 = v_10582 | v_10590;
  assign v_10582 = mux_10582(v_8450);
  assign v_10584 = v_10585 | v_10587;
  assign v_10585 = mux_10585(v_10586);
  assign v_10586 = ~act_8473;
  assign v_10587 = v_10588 | v_10589;
  assign v_10588 = mux_10588(v_1450);
  assign v_10589 = mux_10589(v_1444);
  assign v_10590 = mux_10590(v_8463);
  assign v_10592 = v_10593 | v_10595;
  assign v_10593 = mux_10593(v_10594);
  assign v_10594 = ~act_8456;
  assign v_10595 = v_10596 | v_10597;
  assign v_10596 = mux_10596(v_1436);
  assign v_10597 = mux_10597(v_1430);
  assign v_10598 = mux_10598(v_8439);
  assign v_10600 = v_10601 | v_10603;
  assign v_10601 = mux_10601(v_10602);
  assign v_10602 = ~act_8396;
  assign v_10603 = v_10604 | v_10612;
  assign v_10604 = mux_10604(v_8397);
  assign v_10606 = v_10607 | v_10609;
  assign v_10607 = mux_10607(v_10608);
  assign v_10608 = ~act_8420;
  assign v_10609 = v_10610 | v_10611;
  assign v_10610 = mux_10610(v_1422);
  assign v_10611 = mux_10611(v_1416);
  assign v_10612 = mux_10612(v_8410);
  assign v_10614 = v_10615 | v_10617;
  assign v_10615 = mux_10615(v_10616);
  assign v_10616 = ~act_8403;
  assign v_10617 = v_10618 | v_10619;
  assign v_10618 = mux_10618(v_1408);
  assign v_10619 = mux_10619(v_1402);
  assign v_10620 = mux_10620(v_8379);
  assign v_10622 = v_10623 | v_10625;
  assign v_10623 = mux_10623(v_10624);
  assign v_10624 = ~act_8264;
  assign v_10625 = v_10626 | v_10648;
  assign v_10626 = mux_10626(v_8265);
  assign v_10628 = v_10629 | v_10631;
  assign v_10629 = mux_10629(v_10630);
  assign v_10630 = ~act_8324;
  assign v_10631 = v_10632 | v_10640;
  assign v_10632 = mux_10632(v_8325);
  assign v_10634 = v_10635 | v_10637;
  assign v_10635 = mux_10635(v_10636);
  assign v_10636 = ~act_8348;
  assign v_10637 = v_10638 | v_10639;
  assign v_10638 = mux_10638(v_1394);
  assign v_10639 = mux_10639(v_1388);
  assign v_10640 = mux_10640(v_8338);
  assign v_10642 = v_10643 | v_10645;
  assign v_10643 = mux_10643(v_10644);
  assign v_10644 = ~act_8331;
  assign v_10645 = v_10646 | v_10647;
  assign v_10646 = mux_10646(v_1380);
  assign v_10647 = mux_10647(v_1374);
  assign v_10648 = mux_10648(v_8314);
  assign v_10650 = v_10651 | v_10653;
  assign v_10651 = mux_10651(v_10652);
  assign v_10652 = ~act_8271;
  assign v_10653 = v_10654 | v_10662;
  assign v_10654 = mux_10654(v_8272);
  assign v_10656 = v_10657 | v_10659;
  assign v_10657 = mux_10657(v_10658);
  assign v_10658 = ~act_8295;
  assign v_10659 = v_10660 | v_10661;
  assign v_10660 = mux_10660(v_1366);
  assign v_10661 = mux_10661(v_1360);
  assign v_10662 = mux_10662(v_8285);
  assign v_10664 = v_10665 | v_10667;
  assign v_10665 = mux_10665(v_10666);
  assign v_10666 = ~act_8278;
  assign v_10667 = v_10668 | v_10669;
  assign v_10668 = mux_10668(v_1352);
  assign v_10669 = mux_10669(v_1346);
  assign v_10670 = mux_10670(v_8240);
  assign v_10672 = v_10673 | v_10675;
  assign v_10673 = mux_10673(v_10674);
  assign v_10674 = ~act_7693;
  assign v_10675 = v_10676 | v_10782;
  assign v_10676 = mux_10676(v_7694);
  assign v_10678 = v_10679 | v_10681;
  assign v_10679 = mux_10679(v_10680);
  assign v_10680 = ~act_7969;
  assign v_10681 = v_10682 | v_10732;
  assign v_10682 = mux_10682(v_7970);
  assign v_10684 = v_10685 | v_10687;
  assign v_10685 = mux_10685(v_10686);
  assign v_10686 = ~act_8101;
  assign v_10687 = v_10688 | v_10710;
  assign v_10688 = mux_10688(v_8102);
  assign v_10690 = v_10691 | v_10693;
  assign v_10691 = mux_10691(v_10692);
  assign v_10692 = ~act_8161;
  assign v_10693 = v_10694 | v_10702;
  assign v_10694 = mux_10694(v_8162);
  assign v_10696 = v_10697 | v_10699;
  assign v_10697 = mux_10697(v_10698);
  assign v_10698 = ~act_8185;
  assign v_10699 = v_10700 | v_10701;
  assign v_10700 = mux_10700(v_1338);
  assign v_10701 = mux_10701(v_1332);
  assign v_10702 = mux_10702(v_8175);
  assign v_10704 = v_10705 | v_10707;
  assign v_10705 = mux_10705(v_10706);
  assign v_10706 = ~act_8168;
  assign v_10707 = v_10708 | v_10709;
  assign v_10708 = mux_10708(v_1324);
  assign v_10709 = mux_10709(v_1318);
  assign v_10710 = mux_10710(v_8151);
  assign v_10712 = v_10713 | v_10715;
  assign v_10713 = mux_10713(v_10714);
  assign v_10714 = ~act_8108;
  assign v_10715 = v_10716 | v_10724;
  assign v_10716 = mux_10716(v_8109);
  assign v_10718 = v_10719 | v_10721;
  assign v_10719 = mux_10719(v_10720);
  assign v_10720 = ~act_8132;
  assign v_10721 = v_10722 | v_10723;
  assign v_10722 = mux_10722(v_1310);
  assign v_10723 = mux_10723(v_1304);
  assign v_10724 = mux_10724(v_8122);
  assign v_10726 = v_10727 | v_10729;
  assign v_10727 = mux_10727(v_10728);
  assign v_10728 = ~act_8115;
  assign v_10729 = v_10730 | v_10731;
  assign v_10730 = mux_10730(v_1296);
  assign v_10731 = mux_10731(v_1290);
  assign v_10732 = mux_10732(v_8091);
  assign v_10734 = v_10735 | v_10737;
  assign v_10735 = mux_10735(v_10736);
  assign v_10736 = ~act_7976;
  assign v_10737 = v_10738 | v_10760;
  assign v_10738 = mux_10738(v_7977);
  assign v_10740 = v_10741 | v_10743;
  assign v_10741 = mux_10741(v_10742);
  assign v_10742 = ~act_8036;
  assign v_10743 = v_10744 | v_10752;
  assign v_10744 = mux_10744(v_8037);
  assign v_10746 = v_10747 | v_10749;
  assign v_10747 = mux_10747(v_10748);
  assign v_10748 = ~act_8060;
  assign v_10749 = v_10750 | v_10751;
  assign v_10750 = mux_10750(v_1282);
  assign v_10751 = mux_10751(v_1276);
  assign v_10752 = mux_10752(v_8050);
  assign v_10754 = v_10755 | v_10757;
  assign v_10755 = mux_10755(v_10756);
  assign v_10756 = ~act_8043;
  assign v_10757 = v_10758 | v_10759;
  assign v_10758 = mux_10758(v_1268);
  assign v_10759 = mux_10759(v_1262);
  assign v_10760 = mux_10760(v_8026);
  assign v_10762 = v_10763 | v_10765;
  assign v_10763 = mux_10763(v_10764);
  assign v_10764 = ~act_7983;
  assign v_10765 = v_10766 | v_10774;
  assign v_10766 = mux_10766(v_7984);
  assign v_10768 = v_10769 | v_10771;
  assign v_10769 = mux_10769(v_10770);
  assign v_10770 = ~act_8007;
  assign v_10771 = v_10772 | v_10773;
  assign v_10772 = mux_10772(v_1254);
  assign v_10773 = mux_10773(v_1248);
  assign v_10774 = mux_10774(v_7997);
  assign v_10776 = v_10777 | v_10779;
  assign v_10777 = mux_10777(v_10778);
  assign v_10778 = ~act_7990;
  assign v_10779 = v_10780 | v_10781;
  assign v_10780 = mux_10780(v_1240);
  assign v_10781 = mux_10781(v_1234);
  assign v_10782 = mux_10782(v_7959);
  assign v_10784 = v_10785 | v_10787;
  assign v_10785 = mux_10785(v_10786);
  assign v_10786 = ~act_7700;
  assign v_10787 = v_10788 | v_10838;
  assign v_10788 = mux_10788(v_7701);
  assign v_10790 = v_10791 | v_10793;
  assign v_10791 = mux_10791(v_10792);
  assign v_10792 = ~act_7832;
  assign v_10793 = v_10794 | v_10816;
  assign v_10794 = mux_10794(v_7833);
  assign v_10796 = v_10797 | v_10799;
  assign v_10797 = mux_10797(v_10798);
  assign v_10798 = ~act_7892;
  assign v_10799 = v_10800 | v_10808;
  assign v_10800 = mux_10800(v_7893);
  assign v_10802 = v_10803 | v_10805;
  assign v_10803 = mux_10803(v_10804);
  assign v_10804 = ~act_7916;
  assign v_10805 = v_10806 | v_10807;
  assign v_10806 = mux_10806(v_1226);
  assign v_10807 = mux_10807(v_1220);
  assign v_10808 = mux_10808(v_7906);
  assign v_10810 = v_10811 | v_10813;
  assign v_10811 = mux_10811(v_10812);
  assign v_10812 = ~act_7899;
  assign v_10813 = v_10814 | v_10815;
  assign v_10814 = mux_10814(v_1212);
  assign v_10815 = mux_10815(v_1206);
  assign v_10816 = mux_10816(v_7882);
  assign v_10818 = v_10819 | v_10821;
  assign v_10819 = mux_10819(v_10820);
  assign v_10820 = ~act_7839;
  assign v_10821 = v_10822 | v_10830;
  assign v_10822 = mux_10822(v_7840);
  assign v_10824 = v_10825 | v_10827;
  assign v_10825 = mux_10825(v_10826);
  assign v_10826 = ~act_7863;
  assign v_10827 = v_10828 | v_10829;
  assign v_10828 = mux_10828(v_1198);
  assign v_10829 = mux_10829(v_1192);
  assign v_10830 = mux_10830(v_7853);
  assign v_10832 = v_10833 | v_10835;
  assign v_10833 = mux_10833(v_10834);
  assign v_10834 = ~act_7846;
  assign v_10835 = v_10836 | v_10837;
  assign v_10836 = mux_10836(v_1184);
  assign v_10837 = mux_10837(v_1178);
  assign v_10838 = mux_10838(v_7822);
  assign v_10840 = v_10841 | v_10843;
  assign v_10841 = mux_10841(v_10842);
  assign v_10842 = ~act_7707;
  assign v_10843 = v_10844 | v_10866;
  assign v_10844 = mux_10844(v_7708);
  assign v_10846 = v_10847 | v_10849;
  assign v_10847 = mux_10847(v_10848);
  assign v_10848 = ~act_7767;
  assign v_10849 = v_10850 | v_10858;
  assign v_10850 = mux_10850(v_7768);
  assign v_10852 = v_10853 | v_10855;
  assign v_10853 = mux_10853(v_10854);
  assign v_10854 = ~act_7791;
  assign v_10855 = v_10856 | v_10857;
  assign v_10856 = mux_10856(v_1170);
  assign v_10857 = mux_10857(v_1164);
  assign v_10858 = mux_10858(v_7781);
  assign v_10860 = v_10861 | v_10863;
  assign v_10861 = mux_10861(v_10862);
  assign v_10862 = ~act_7774;
  assign v_10863 = v_10864 | v_10865;
  assign v_10864 = mux_10864(v_1156);
  assign v_10865 = mux_10865(v_1150);
  assign v_10866 = mux_10866(v_7757);
  assign v_10868 = v_10869 | v_10871;
  assign v_10869 = mux_10869(v_10870);
  assign v_10870 = ~act_7714;
  assign v_10871 = v_10872 | v_10880;
  assign v_10872 = mux_10872(v_7715);
  assign v_10874 = v_10875 | v_10877;
  assign v_10875 = mux_10875(v_10876);
  assign v_10876 = ~act_7738;
  assign v_10877 = v_10878 | v_10879;
  assign v_10878 = mux_10878(v_1142);
  assign v_10879 = mux_10879(v_1136);
  assign v_10880 = mux_10880(v_7728);
  assign v_10882 = v_10883 | v_10885;
  assign v_10883 = mux_10883(v_10884);
  assign v_10884 = ~act_7721;
  assign v_10885 = v_10886 | v_10887;
  assign v_10886 = mux_10886(v_1128);
  assign v_10887 = mux_10887(v_1122);
  assign v_10888 = mux_10888(v_7669);
  assign v_10890 = v_10891 | v_10893;
  assign v_10891 = mux_10891(v_10892);
  assign v_10892 = ~act_5394;
  assign v_10893 = v_10894 | v_11336;
  assign v_10894 = mux_10894(v_5395);
  assign v_10896 = v_10897 | v_10899;
  assign v_10897 = mux_10897(v_10898);
  assign v_10898 = ~act_6534;
  assign v_10899 = v_10900 | v_11118;
  assign v_10900 = mux_10900(v_6535);
  assign v_10902 = v_10903 | v_10905;
  assign v_10903 = mux_10903(v_10904);
  assign v_10904 = ~act_7098;
  assign v_10905 = v_10906 | v_11012;
  assign v_10906 = mux_10906(v_7099);
  assign v_10908 = v_10909 | v_10911;
  assign v_10909 = mux_10909(v_10910);
  assign v_10910 = ~act_7374;
  assign v_10911 = v_10912 | v_10962;
  assign v_10912 = mux_10912(v_7375);
  assign v_10914 = v_10915 | v_10917;
  assign v_10915 = mux_10915(v_10916);
  assign v_10916 = ~act_7506;
  assign v_10917 = v_10918 | v_10940;
  assign v_10918 = mux_10918(v_7507);
  assign v_10920 = v_10921 | v_10923;
  assign v_10921 = mux_10921(v_10922);
  assign v_10922 = ~act_7566;
  assign v_10923 = v_10924 | v_10932;
  assign v_10924 = mux_10924(v_7567);
  assign v_10926 = v_10927 | v_10929;
  assign v_10927 = mux_10927(v_10928);
  assign v_10928 = ~act_7590;
  assign v_10929 = v_10930 | v_10931;
  assign v_10930 = mux_10930(v_1114);
  assign v_10931 = mux_10931(v_1108);
  assign v_10932 = mux_10932(v_7580);
  assign v_10934 = v_10935 | v_10937;
  assign v_10935 = mux_10935(v_10936);
  assign v_10936 = ~act_7573;
  assign v_10937 = v_10938 | v_10939;
  assign v_10938 = mux_10938(v_1100);
  assign v_10939 = mux_10939(v_1094);
  assign v_10940 = mux_10940(v_7556);
  assign v_10942 = v_10943 | v_10945;
  assign v_10943 = mux_10943(v_10944);
  assign v_10944 = ~act_7513;
  assign v_10945 = v_10946 | v_10954;
  assign v_10946 = mux_10946(v_7514);
  assign v_10948 = v_10949 | v_10951;
  assign v_10949 = mux_10949(v_10950);
  assign v_10950 = ~act_7537;
  assign v_10951 = v_10952 | v_10953;
  assign v_10952 = mux_10952(v_1086);
  assign v_10953 = mux_10953(v_1080);
  assign v_10954 = mux_10954(v_7527);
  assign v_10956 = v_10957 | v_10959;
  assign v_10957 = mux_10957(v_10958);
  assign v_10958 = ~act_7520;
  assign v_10959 = v_10960 | v_10961;
  assign v_10960 = mux_10960(v_1072);
  assign v_10961 = mux_10961(v_1066);
  assign v_10962 = mux_10962(v_7496);
  assign v_10964 = v_10965 | v_10967;
  assign v_10965 = mux_10965(v_10966);
  assign v_10966 = ~act_7381;
  assign v_10967 = v_10968 | v_10990;
  assign v_10968 = mux_10968(v_7382);
  assign v_10970 = v_10971 | v_10973;
  assign v_10971 = mux_10971(v_10972);
  assign v_10972 = ~act_7441;
  assign v_10973 = v_10974 | v_10982;
  assign v_10974 = mux_10974(v_7442);
  assign v_10976 = v_10977 | v_10979;
  assign v_10977 = mux_10977(v_10978);
  assign v_10978 = ~act_7465;
  assign v_10979 = v_10980 | v_10981;
  assign v_10980 = mux_10980(v_1058);
  assign v_10981 = mux_10981(v_1052);
  assign v_10982 = mux_10982(v_7455);
  assign v_10984 = v_10985 | v_10987;
  assign v_10985 = mux_10985(v_10986);
  assign v_10986 = ~act_7448;
  assign v_10987 = v_10988 | v_10989;
  assign v_10988 = mux_10988(v_1044);
  assign v_10989 = mux_10989(v_1038);
  assign v_10990 = mux_10990(v_7431);
  assign v_10992 = v_10993 | v_10995;
  assign v_10993 = mux_10993(v_10994);
  assign v_10994 = ~act_7388;
  assign v_10995 = v_10996 | v_11004;
  assign v_10996 = mux_10996(v_7389);
  assign v_10998 = v_10999 | v_11001;
  assign v_10999 = mux_10999(v_11000);
  assign v_11000 = ~act_7412;
  assign v_11001 = v_11002 | v_11003;
  assign v_11002 = mux_11002(v_1030);
  assign v_11003 = mux_11003(v_1024);
  assign v_11004 = mux_11004(v_7402);
  assign v_11006 = v_11007 | v_11009;
  assign v_11007 = mux_11007(v_11008);
  assign v_11008 = ~act_7395;
  assign v_11009 = v_11010 | v_11011;
  assign v_11010 = mux_11010(v_1016);
  assign v_11011 = mux_11011(v_1010);
  assign v_11012 = mux_11012(v_7364);
  assign v_11014 = v_11015 | v_11017;
  assign v_11015 = mux_11015(v_11016);
  assign v_11016 = ~act_7105;
  assign v_11017 = v_11018 | v_11068;
  assign v_11018 = mux_11018(v_7106);
  assign v_11020 = v_11021 | v_11023;
  assign v_11021 = mux_11021(v_11022);
  assign v_11022 = ~act_7237;
  assign v_11023 = v_11024 | v_11046;
  assign v_11024 = mux_11024(v_7238);
  assign v_11026 = v_11027 | v_11029;
  assign v_11027 = mux_11027(v_11028);
  assign v_11028 = ~act_7297;
  assign v_11029 = v_11030 | v_11038;
  assign v_11030 = mux_11030(v_7298);
  assign v_11032 = v_11033 | v_11035;
  assign v_11033 = mux_11033(v_11034);
  assign v_11034 = ~act_7321;
  assign v_11035 = v_11036 | v_11037;
  assign v_11036 = mux_11036(v_1002);
  assign v_11037 = mux_11037(v_996);
  assign v_11038 = mux_11038(v_7311);
  assign v_11040 = v_11041 | v_11043;
  assign v_11041 = mux_11041(v_11042);
  assign v_11042 = ~act_7304;
  assign v_11043 = v_11044 | v_11045;
  assign v_11044 = mux_11044(v_988);
  assign v_11045 = mux_11045(v_982);
  assign v_11046 = mux_11046(v_7287);
  assign v_11048 = v_11049 | v_11051;
  assign v_11049 = mux_11049(v_11050);
  assign v_11050 = ~act_7244;
  assign v_11051 = v_11052 | v_11060;
  assign v_11052 = mux_11052(v_7245);
  assign v_11054 = v_11055 | v_11057;
  assign v_11055 = mux_11055(v_11056);
  assign v_11056 = ~act_7268;
  assign v_11057 = v_11058 | v_11059;
  assign v_11058 = mux_11058(v_974);
  assign v_11059 = mux_11059(v_968);
  assign v_11060 = mux_11060(v_7258);
  assign v_11062 = v_11063 | v_11065;
  assign v_11063 = mux_11063(v_11064);
  assign v_11064 = ~act_7251;
  assign v_11065 = v_11066 | v_11067;
  assign v_11066 = mux_11066(v_960);
  assign v_11067 = mux_11067(v_954);
  assign v_11068 = mux_11068(v_7227);
  assign v_11070 = v_11071 | v_11073;
  assign v_11071 = mux_11071(v_11072);
  assign v_11072 = ~act_7112;
  assign v_11073 = v_11074 | v_11096;
  assign v_11074 = mux_11074(v_7113);
  assign v_11076 = v_11077 | v_11079;
  assign v_11077 = mux_11077(v_11078);
  assign v_11078 = ~act_7172;
  assign v_11079 = v_11080 | v_11088;
  assign v_11080 = mux_11080(v_7173);
  assign v_11082 = v_11083 | v_11085;
  assign v_11083 = mux_11083(v_11084);
  assign v_11084 = ~act_7196;
  assign v_11085 = v_11086 | v_11087;
  assign v_11086 = mux_11086(v_946);
  assign v_11087 = mux_11087(v_940);
  assign v_11088 = mux_11088(v_7186);
  assign v_11090 = v_11091 | v_11093;
  assign v_11091 = mux_11091(v_11092);
  assign v_11092 = ~act_7179;
  assign v_11093 = v_11094 | v_11095;
  assign v_11094 = mux_11094(v_932);
  assign v_11095 = mux_11095(v_926);
  assign v_11096 = mux_11096(v_7162);
  assign v_11098 = v_11099 | v_11101;
  assign v_11099 = mux_11099(v_11100);
  assign v_11100 = ~act_7119;
  assign v_11101 = v_11102 | v_11110;
  assign v_11102 = mux_11102(v_7120);
  assign v_11104 = v_11105 | v_11107;
  assign v_11105 = mux_11105(v_11106);
  assign v_11106 = ~act_7143;
  assign v_11107 = v_11108 | v_11109;
  assign v_11108 = mux_11108(v_918);
  assign v_11109 = mux_11109(v_912);
  assign v_11110 = mux_11110(v_7133);
  assign v_11112 = v_11113 | v_11115;
  assign v_11113 = mux_11113(v_11114);
  assign v_11114 = ~act_7126;
  assign v_11115 = v_11116 | v_11117;
  assign v_11116 = mux_11116(v_904);
  assign v_11117 = mux_11117(v_898);
  assign v_11118 = mux_11118(v_7088);
  assign v_11120 = v_11121 | v_11123;
  assign v_11121 = mux_11121(v_11122);
  assign v_11122 = ~act_6541;
  assign v_11123 = v_11124 | v_11230;
  assign v_11124 = mux_11124(v_6542);
  assign v_11126 = v_11127 | v_11129;
  assign v_11127 = mux_11127(v_11128);
  assign v_11128 = ~act_6817;
  assign v_11129 = v_11130 | v_11180;
  assign v_11130 = mux_11130(v_6818);
  assign v_11132 = v_11133 | v_11135;
  assign v_11133 = mux_11133(v_11134);
  assign v_11134 = ~act_6949;
  assign v_11135 = v_11136 | v_11158;
  assign v_11136 = mux_11136(v_6950);
  assign v_11138 = v_11139 | v_11141;
  assign v_11139 = mux_11139(v_11140);
  assign v_11140 = ~act_7009;
  assign v_11141 = v_11142 | v_11150;
  assign v_11142 = mux_11142(v_7010);
  assign v_11144 = v_11145 | v_11147;
  assign v_11145 = mux_11145(v_11146);
  assign v_11146 = ~act_7033;
  assign v_11147 = v_11148 | v_11149;
  assign v_11148 = mux_11148(v_890);
  assign v_11149 = mux_11149(v_884);
  assign v_11150 = mux_11150(v_7023);
  assign v_11152 = v_11153 | v_11155;
  assign v_11153 = mux_11153(v_11154);
  assign v_11154 = ~act_7016;
  assign v_11155 = v_11156 | v_11157;
  assign v_11156 = mux_11156(v_876);
  assign v_11157 = mux_11157(v_870);
  assign v_11158 = mux_11158(v_6999);
  assign v_11160 = v_11161 | v_11163;
  assign v_11161 = mux_11161(v_11162);
  assign v_11162 = ~act_6956;
  assign v_11163 = v_11164 | v_11172;
  assign v_11164 = mux_11164(v_6957);
  assign v_11166 = v_11167 | v_11169;
  assign v_11167 = mux_11167(v_11168);
  assign v_11168 = ~act_6980;
  assign v_11169 = v_11170 | v_11171;
  assign v_11170 = mux_11170(v_862);
  assign v_11171 = mux_11171(v_856);
  assign v_11172 = mux_11172(v_6970);
  assign v_11174 = v_11175 | v_11177;
  assign v_11175 = mux_11175(v_11176);
  assign v_11176 = ~act_6963;
  assign v_11177 = v_11178 | v_11179;
  assign v_11178 = mux_11178(v_848);
  assign v_11179 = mux_11179(v_842);
  assign v_11180 = mux_11180(v_6939);
  assign v_11182 = v_11183 | v_11185;
  assign v_11183 = mux_11183(v_11184);
  assign v_11184 = ~act_6824;
  assign v_11185 = v_11186 | v_11208;
  assign v_11186 = mux_11186(v_6825);
  assign v_11188 = v_11189 | v_11191;
  assign v_11189 = mux_11189(v_11190);
  assign v_11190 = ~act_6884;
  assign v_11191 = v_11192 | v_11200;
  assign v_11192 = mux_11192(v_6885);
  assign v_11194 = v_11195 | v_11197;
  assign v_11195 = mux_11195(v_11196);
  assign v_11196 = ~act_6908;
  assign v_11197 = v_11198 | v_11199;
  assign v_11198 = mux_11198(v_834);
  assign v_11199 = mux_11199(v_828);
  assign v_11200 = mux_11200(v_6898);
  assign v_11202 = v_11203 | v_11205;
  assign v_11203 = mux_11203(v_11204);
  assign v_11204 = ~act_6891;
  assign v_11205 = v_11206 | v_11207;
  assign v_11206 = mux_11206(v_820);
  assign v_11207 = mux_11207(v_814);
  assign v_11208 = mux_11208(v_6874);
  assign v_11210 = v_11211 | v_11213;
  assign v_11211 = mux_11211(v_11212);
  assign v_11212 = ~act_6831;
  assign v_11213 = v_11214 | v_11222;
  assign v_11214 = mux_11214(v_6832);
  assign v_11216 = v_11217 | v_11219;
  assign v_11217 = mux_11217(v_11218);
  assign v_11218 = ~act_6855;
  assign v_11219 = v_11220 | v_11221;
  assign v_11220 = mux_11220(v_806);
  assign v_11221 = mux_11221(v_800);
  assign v_11222 = mux_11222(v_6845);
  assign v_11224 = v_11225 | v_11227;
  assign v_11225 = mux_11225(v_11226);
  assign v_11226 = ~act_6838;
  assign v_11227 = v_11228 | v_11229;
  assign v_11228 = mux_11228(v_792);
  assign v_11229 = mux_11229(v_786);
  assign v_11230 = mux_11230(v_6807);
  assign v_11232 = v_11233 | v_11235;
  assign v_11233 = mux_11233(v_11234);
  assign v_11234 = ~act_6548;
  assign v_11235 = v_11236 | v_11286;
  assign v_11236 = mux_11236(v_6549);
  assign v_11238 = v_11239 | v_11241;
  assign v_11239 = mux_11239(v_11240);
  assign v_11240 = ~act_6680;
  assign v_11241 = v_11242 | v_11264;
  assign v_11242 = mux_11242(v_6681);
  assign v_11244 = v_11245 | v_11247;
  assign v_11245 = mux_11245(v_11246);
  assign v_11246 = ~act_6740;
  assign v_11247 = v_11248 | v_11256;
  assign v_11248 = mux_11248(v_6741);
  assign v_11250 = v_11251 | v_11253;
  assign v_11251 = mux_11251(v_11252);
  assign v_11252 = ~act_6764;
  assign v_11253 = v_11254 | v_11255;
  assign v_11254 = mux_11254(v_778);
  assign v_11255 = mux_11255(v_772);
  assign v_11256 = mux_11256(v_6754);
  assign v_11258 = v_11259 | v_11261;
  assign v_11259 = mux_11259(v_11260);
  assign v_11260 = ~act_6747;
  assign v_11261 = v_11262 | v_11263;
  assign v_11262 = mux_11262(v_764);
  assign v_11263 = mux_11263(v_758);
  assign v_11264 = mux_11264(v_6730);
  assign v_11266 = v_11267 | v_11269;
  assign v_11267 = mux_11267(v_11268);
  assign v_11268 = ~act_6687;
  assign v_11269 = v_11270 | v_11278;
  assign v_11270 = mux_11270(v_6688);
  assign v_11272 = v_11273 | v_11275;
  assign v_11273 = mux_11273(v_11274);
  assign v_11274 = ~act_6711;
  assign v_11275 = v_11276 | v_11277;
  assign v_11276 = mux_11276(v_750);
  assign v_11277 = mux_11277(v_744);
  assign v_11278 = mux_11278(v_6701);
  assign v_11280 = v_11281 | v_11283;
  assign v_11281 = mux_11281(v_11282);
  assign v_11282 = ~act_6694;
  assign v_11283 = v_11284 | v_11285;
  assign v_11284 = mux_11284(v_736);
  assign v_11285 = mux_11285(v_730);
  assign v_11286 = mux_11286(v_6670);
  assign v_11288 = v_11289 | v_11291;
  assign v_11289 = mux_11289(v_11290);
  assign v_11290 = ~act_6555;
  assign v_11291 = v_11292 | v_11314;
  assign v_11292 = mux_11292(v_6556);
  assign v_11294 = v_11295 | v_11297;
  assign v_11295 = mux_11295(v_11296);
  assign v_11296 = ~act_6615;
  assign v_11297 = v_11298 | v_11306;
  assign v_11298 = mux_11298(v_6616);
  assign v_11300 = v_11301 | v_11303;
  assign v_11301 = mux_11301(v_11302);
  assign v_11302 = ~act_6639;
  assign v_11303 = v_11304 | v_11305;
  assign v_11304 = mux_11304(v_722);
  assign v_11305 = mux_11305(v_716);
  assign v_11306 = mux_11306(v_6629);
  assign v_11308 = v_11309 | v_11311;
  assign v_11309 = mux_11309(v_11310);
  assign v_11310 = ~act_6622;
  assign v_11311 = v_11312 | v_11313;
  assign v_11312 = mux_11312(v_708);
  assign v_11313 = mux_11313(v_702);
  assign v_11314 = mux_11314(v_6605);
  assign v_11316 = v_11317 | v_11319;
  assign v_11317 = mux_11317(v_11318);
  assign v_11318 = ~act_6562;
  assign v_11319 = v_11320 | v_11328;
  assign v_11320 = mux_11320(v_6563);
  assign v_11322 = v_11323 | v_11325;
  assign v_11323 = mux_11323(v_11324);
  assign v_11324 = ~act_6586;
  assign v_11325 = v_11326 | v_11327;
  assign v_11326 = mux_11326(v_694);
  assign v_11327 = mux_11327(v_688);
  assign v_11328 = mux_11328(v_6576);
  assign v_11330 = v_11331 | v_11333;
  assign v_11331 = mux_11331(v_11332);
  assign v_11332 = ~act_6569;
  assign v_11333 = v_11334 | v_11335;
  assign v_11334 = mux_11334(v_680);
  assign v_11335 = mux_11335(v_674);
  assign v_11336 = mux_11336(v_6524);
  assign v_11338 = v_11339 | v_11341;
  assign v_11339 = mux_11339(v_11340);
  assign v_11340 = ~act_5401;
  assign v_11341 = v_11342 | v_11560;
  assign v_11342 = mux_11342(v_5402);
  assign v_11344 = v_11345 | v_11347;
  assign v_11345 = mux_11345(v_11346);
  assign v_11346 = ~act_5965;
  assign v_11347 = v_11348 | v_11454;
  assign v_11348 = mux_11348(v_5966);
  assign v_11350 = v_11351 | v_11353;
  assign v_11351 = mux_11351(v_11352);
  assign v_11352 = ~act_6241;
  assign v_11353 = v_11354 | v_11404;
  assign v_11354 = mux_11354(v_6242);
  assign v_11356 = v_11357 | v_11359;
  assign v_11357 = mux_11357(v_11358);
  assign v_11358 = ~act_6373;
  assign v_11359 = v_11360 | v_11382;
  assign v_11360 = mux_11360(v_6374);
  assign v_11362 = v_11363 | v_11365;
  assign v_11363 = mux_11363(v_11364);
  assign v_11364 = ~act_6433;
  assign v_11365 = v_11366 | v_11374;
  assign v_11366 = mux_11366(v_6434);
  assign v_11368 = v_11369 | v_11371;
  assign v_11369 = mux_11369(v_11370);
  assign v_11370 = ~act_6457;
  assign v_11371 = v_11372 | v_11373;
  assign v_11372 = mux_11372(v_666);
  assign v_11373 = mux_11373(v_660);
  assign v_11374 = mux_11374(v_6447);
  assign v_11376 = v_11377 | v_11379;
  assign v_11377 = mux_11377(v_11378);
  assign v_11378 = ~act_6440;
  assign v_11379 = v_11380 | v_11381;
  assign v_11380 = mux_11380(v_652);
  assign v_11381 = mux_11381(v_646);
  assign v_11382 = mux_11382(v_6423);
  assign v_11384 = v_11385 | v_11387;
  assign v_11385 = mux_11385(v_11386);
  assign v_11386 = ~act_6380;
  assign v_11387 = v_11388 | v_11396;
  assign v_11388 = mux_11388(v_6381);
  assign v_11390 = v_11391 | v_11393;
  assign v_11391 = mux_11391(v_11392);
  assign v_11392 = ~act_6404;
  assign v_11393 = v_11394 | v_11395;
  assign v_11394 = mux_11394(v_638);
  assign v_11395 = mux_11395(v_632);
  assign v_11396 = mux_11396(v_6394);
  assign v_11398 = v_11399 | v_11401;
  assign v_11399 = mux_11399(v_11400);
  assign v_11400 = ~act_6387;
  assign v_11401 = v_11402 | v_11403;
  assign v_11402 = mux_11402(v_624);
  assign v_11403 = mux_11403(v_618);
  assign v_11404 = mux_11404(v_6363);
  assign v_11406 = v_11407 | v_11409;
  assign v_11407 = mux_11407(v_11408);
  assign v_11408 = ~act_6248;
  assign v_11409 = v_11410 | v_11432;
  assign v_11410 = mux_11410(v_6249);
  assign v_11412 = v_11413 | v_11415;
  assign v_11413 = mux_11413(v_11414);
  assign v_11414 = ~act_6308;
  assign v_11415 = v_11416 | v_11424;
  assign v_11416 = mux_11416(v_6309);
  assign v_11418 = v_11419 | v_11421;
  assign v_11419 = mux_11419(v_11420);
  assign v_11420 = ~act_6332;
  assign v_11421 = v_11422 | v_11423;
  assign v_11422 = mux_11422(v_610);
  assign v_11423 = mux_11423(v_604);
  assign v_11424 = mux_11424(v_6322);
  assign v_11426 = v_11427 | v_11429;
  assign v_11427 = mux_11427(v_11428);
  assign v_11428 = ~act_6315;
  assign v_11429 = v_11430 | v_11431;
  assign v_11430 = mux_11430(v_596);
  assign v_11431 = mux_11431(v_590);
  assign v_11432 = mux_11432(v_6298);
  assign v_11434 = v_11435 | v_11437;
  assign v_11435 = mux_11435(v_11436);
  assign v_11436 = ~act_6255;
  assign v_11437 = v_11438 | v_11446;
  assign v_11438 = mux_11438(v_6256);
  assign v_11440 = v_11441 | v_11443;
  assign v_11441 = mux_11441(v_11442);
  assign v_11442 = ~act_6279;
  assign v_11443 = v_11444 | v_11445;
  assign v_11444 = mux_11444(v_582);
  assign v_11445 = mux_11445(v_576);
  assign v_11446 = mux_11446(v_6269);
  assign v_11448 = v_11449 | v_11451;
  assign v_11449 = mux_11449(v_11450);
  assign v_11450 = ~act_6262;
  assign v_11451 = v_11452 | v_11453;
  assign v_11452 = mux_11452(v_568);
  assign v_11453 = mux_11453(v_562);
  assign v_11454 = mux_11454(v_6231);
  assign v_11456 = v_11457 | v_11459;
  assign v_11457 = mux_11457(v_11458);
  assign v_11458 = ~act_5972;
  assign v_11459 = v_11460 | v_11510;
  assign v_11460 = mux_11460(v_5973);
  assign v_11462 = v_11463 | v_11465;
  assign v_11463 = mux_11463(v_11464);
  assign v_11464 = ~act_6104;
  assign v_11465 = v_11466 | v_11488;
  assign v_11466 = mux_11466(v_6105);
  assign v_11468 = v_11469 | v_11471;
  assign v_11469 = mux_11469(v_11470);
  assign v_11470 = ~act_6164;
  assign v_11471 = v_11472 | v_11480;
  assign v_11472 = mux_11472(v_6165);
  assign v_11474 = v_11475 | v_11477;
  assign v_11475 = mux_11475(v_11476);
  assign v_11476 = ~act_6188;
  assign v_11477 = v_11478 | v_11479;
  assign v_11478 = mux_11478(v_554);
  assign v_11479 = mux_11479(v_548);
  assign v_11480 = mux_11480(v_6178);
  assign v_11482 = v_11483 | v_11485;
  assign v_11483 = mux_11483(v_11484);
  assign v_11484 = ~act_6171;
  assign v_11485 = v_11486 | v_11487;
  assign v_11486 = mux_11486(v_540);
  assign v_11487 = mux_11487(v_534);
  assign v_11488 = mux_11488(v_6154);
  assign v_11490 = v_11491 | v_11493;
  assign v_11491 = mux_11491(v_11492);
  assign v_11492 = ~act_6111;
  assign v_11493 = v_11494 | v_11502;
  assign v_11494 = mux_11494(v_6112);
  assign v_11496 = v_11497 | v_11499;
  assign v_11497 = mux_11497(v_11498);
  assign v_11498 = ~act_6135;
  assign v_11499 = v_11500 | v_11501;
  assign v_11500 = mux_11500(v_526);
  assign v_11501 = mux_11501(v_520);
  assign v_11502 = mux_11502(v_6125);
  assign v_11504 = v_11505 | v_11507;
  assign v_11505 = mux_11505(v_11506);
  assign v_11506 = ~act_6118;
  assign v_11507 = v_11508 | v_11509;
  assign v_11508 = mux_11508(v_512);
  assign v_11509 = mux_11509(v_506);
  assign v_11510 = mux_11510(v_6094);
  assign v_11512 = v_11513 | v_11515;
  assign v_11513 = mux_11513(v_11514);
  assign v_11514 = ~act_5979;
  assign v_11515 = v_11516 | v_11538;
  assign v_11516 = mux_11516(v_5980);
  assign v_11518 = v_11519 | v_11521;
  assign v_11519 = mux_11519(v_11520);
  assign v_11520 = ~act_6039;
  assign v_11521 = v_11522 | v_11530;
  assign v_11522 = mux_11522(v_6040);
  assign v_11524 = v_11525 | v_11527;
  assign v_11525 = mux_11525(v_11526);
  assign v_11526 = ~act_6063;
  assign v_11527 = v_11528 | v_11529;
  assign v_11528 = mux_11528(v_498);
  assign v_11529 = mux_11529(v_492);
  assign v_11530 = mux_11530(v_6053);
  assign v_11532 = v_11533 | v_11535;
  assign v_11533 = mux_11533(v_11534);
  assign v_11534 = ~act_6046;
  assign v_11535 = v_11536 | v_11537;
  assign v_11536 = mux_11536(v_484);
  assign v_11537 = mux_11537(v_478);
  assign v_11538 = mux_11538(v_6029);
  assign v_11540 = v_11541 | v_11543;
  assign v_11541 = mux_11541(v_11542);
  assign v_11542 = ~act_5986;
  assign v_11543 = v_11544 | v_11552;
  assign v_11544 = mux_11544(v_5987);
  assign v_11546 = v_11547 | v_11549;
  assign v_11547 = mux_11547(v_11548);
  assign v_11548 = ~act_6010;
  assign v_11549 = v_11550 | v_11551;
  assign v_11550 = mux_11550(v_470);
  assign v_11551 = mux_11551(v_464);
  assign v_11552 = mux_11552(v_6000);
  assign v_11554 = v_11555 | v_11557;
  assign v_11555 = mux_11555(v_11556);
  assign v_11556 = ~act_5993;
  assign v_11557 = v_11558 | v_11559;
  assign v_11558 = mux_11558(v_456);
  assign v_11559 = mux_11559(v_450);
  assign v_11560 = mux_11560(v_5955);
  assign v_11562 = v_11563 | v_11565;
  assign v_11563 = mux_11563(v_11564);
  assign v_11564 = ~act_5408;
  assign v_11565 = v_11566 | v_11672;
  assign v_11566 = mux_11566(v_5409);
  assign v_11568 = v_11569 | v_11571;
  assign v_11569 = mux_11569(v_11570);
  assign v_11570 = ~act_5684;
  assign v_11571 = v_11572 | v_11622;
  assign v_11572 = mux_11572(v_5685);
  assign v_11574 = v_11575 | v_11577;
  assign v_11575 = mux_11575(v_11576);
  assign v_11576 = ~act_5816;
  assign v_11577 = v_11578 | v_11600;
  assign v_11578 = mux_11578(v_5817);
  assign v_11580 = v_11581 | v_11583;
  assign v_11581 = mux_11581(v_11582);
  assign v_11582 = ~act_5876;
  assign v_11583 = v_11584 | v_11592;
  assign v_11584 = mux_11584(v_5877);
  assign v_11586 = v_11587 | v_11589;
  assign v_11587 = mux_11587(v_11588);
  assign v_11588 = ~act_5900;
  assign v_11589 = v_11590 | v_11591;
  assign v_11590 = mux_11590(v_442);
  assign v_11591 = mux_11591(v_436);
  assign v_11592 = mux_11592(v_5890);
  assign v_11594 = v_11595 | v_11597;
  assign v_11595 = mux_11595(v_11596);
  assign v_11596 = ~act_5883;
  assign v_11597 = v_11598 | v_11599;
  assign v_11598 = mux_11598(v_428);
  assign v_11599 = mux_11599(v_422);
  assign v_11600 = mux_11600(v_5866);
  assign v_11602 = v_11603 | v_11605;
  assign v_11603 = mux_11603(v_11604);
  assign v_11604 = ~act_5823;
  assign v_11605 = v_11606 | v_11614;
  assign v_11606 = mux_11606(v_5824);
  assign v_11608 = v_11609 | v_11611;
  assign v_11609 = mux_11609(v_11610);
  assign v_11610 = ~act_5847;
  assign v_11611 = v_11612 | v_11613;
  assign v_11612 = mux_11612(v_414);
  assign v_11613 = mux_11613(v_408);
  assign v_11614 = mux_11614(v_5837);
  assign v_11616 = v_11617 | v_11619;
  assign v_11617 = mux_11617(v_11618);
  assign v_11618 = ~act_5830;
  assign v_11619 = v_11620 | v_11621;
  assign v_11620 = mux_11620(v_400);
  assign v_11621 = mux_11621(v_394);
  assign v_11622 = mux_11622(v_5806);
  assign v_11624 = v_11625 | v_11627;
  assign v_11625 = mux_11625(v_11626);
  assign v_11626 = ~act_5691;
  assign v_11627 = v_11628 | v_11650;
  assign v_11628 = mux_11628(v_5692);
  assign v_11630 = v_11631 | v_11633;
  assign v_11631 = mux_11631(v_11632);
  assign v_11632 = ~act_5751;
  assign v_11633 = v_11634 | v_11642;
  assign v_11634 = mux_11634(v_5752);
  assign v_11636 = v_11637 | v_11639;
  assign v_11637 = mux_11637(v_11638);
  assign v_11638 = ~act_5775;
  assign v_11639 = v_11640 | v_11641;
  assign v_11640 = mux_11640(v_386);
  assign v_11641 = mux_11641(v_380);
  assign v_11642 = mux_11642(v_5765);
  assign v_11644 = v_11645 | v_11647;
  assign v_11645 = mux_11645(v_11646);
  assign v_11646 = ~act_5758;
  assign v_11647 = v_11648 | v_11649;
  assign v_11648 = mux_11648(v_372);
  assign v_11649 = mux_11649(v_366);
  assign v_11650 = mux_11650(v_5741);
  assign v_11652 = v_11653 | v_11655;
  assign v_11653 = mux_11653(v_11654);
  assign v_11654 = ~act_5698;
  assign v_11655 = v_11656 | v_11664;
  assign v_11656 = mux_11656(v_5699);
  assign v_11658 = v_11659 | v_11661;
  assign v_11659 = mux_11659(v_11660);
  assign v_11660 = ~act_5722;
  assign v_11661 = v_11662 | v_11663;
  assign v_11662 = mux_11662(v_358);
  assign v_11663 = mux_11663(v_352);
  assign v_11664 = mux_11664(v_5712);
  assign v_11666 = v_11667 | v_11669;
  assign v_11667 = mux_11667(v_11668);
  assign v_11668 = ~act_5705;
  assign v_11669 = v_11670 | v_11671;
  assign v_11670 = mux_11670(v_344);
  assign v_11671 = mux_11671(v_338);
  assign v_11672 = mux_11672(v_5674);
  assign v_11674 = v_11675 | v_11677;
  assign v_11675 = mux_11675(v_11676);
  assign v_11676 = ~act_5415;
  assign v_11677 = v_11678 | v_11728;
  assign v_11678 = mux_11678(v_5416);
  assign v_11680 = v_11681 | v_11683;
  assign v_11681 = mux_11681(v_11682);
  assign v_11682 = ~act_5547;
  assign v_11683 = v_11684 | v_11706;
  assign v_11684 = mux_11684(v_5548);
  assign v_11686 = v_11687 | v_11689;
  assign v_11687 = mux_11687(v_11688);
  assign v_11688 = ~act_5607;
  assign v_11689 = v_11690 | v_11698;
  assign v_11690 = mux_11690(v_5608);
  assign v_11692 = v_11693 | v_11695;
  assign v_11693 = mux_11693(v_11694);
  assign v_11694 = ~act_5631;
  assign v_11695 = v_11696 | v_11697;
  assign v_11696 = mux_11696(v_330);
  assign v_11697 = mux_11697(v_324);
  assign v_11698 = mux_11698(v_5621);
  assign v_11700 = v_11701 | v_11703;
  assign v_11701 = mux_11701(v_11702);
  assign v_11702 = ~act_5614;
  assign v_11703 = v_11704 | v_11705;
  assign v_11704 = mux_11704(v_316);
  assign v_11705 = mux_11705(v_310);
  assign v_11706 = mux_11706(v_5597);
  assign v_11708 = v_11709 | v_11711;
  assign v_11709 = mux_11709(v_11710);
  assign v_11710 = ~act_5554;
  assign v_11711 = v_11712 | v_11720;
  assign v_11712 = mux_11712(v_5555);
  assign v_11714 = v_11715 | v_11717;
  assign v_11715 = mux_11715(v_11716);
  assign v_11716 = ~act_5578;
  assign v_11717 = v_11718 | v_11719;
  assign v_11718 = mux_11718(v_302);
  assign v_11719 = mux_11719(v_296);
  assign v_11720 = mux_11720(v_5568);
  assign v_11722 = v_11723 | v_11725;
  assign v_11723 = mux_11723(v_11724);
  assign v_11724 = ~act_5561;
  assign v_11725 = v_11726 | v_11727;
  assign v_11726 = mux_11726(v_288);
  assign v_11727 = mux_11727(v_282);
  assign v_11728 = mux_11728(v_5537);
  assign v_11730 = v_11731 | v_11733;
  assign v_11731 = mux_11731(v_11732);
  assign v_11732 = ~act_5422;
  assign v_11733 = v_11734 | v_11756;
  assign v_11734 = mux_11734(v_5423);
  assign v_11736 = v_11737 | v_11739;
  assign v_11737 = mux_11737(v_11738);
  assign v_11738 = ~act_5482;
  assign v_11739 = v_11740 | v_11748;
  assign v_11740 = mux_11740(v_5483);
  assign v_11742 = v_11743 | v_11745;
  assign v_11743 = mux_11743(v_11744);
  assign v_11744 = ~act_5506;
  assign v_11745 = v_11746 | v_11747;
  assign v_11746 = mux_11746(v_274);
  assign v_11747 = mux_11747(v_268);
  assign v_11748 = mux_11748(v_5496);
  assign v_11750 = v_11751 | v_11753;
  assign v_11751 = mux_11751(v_11752);
  assign v_11752 = ~act_5489;
  assign v_11753 = v_11754 | v_11755;
  assign v_11754 = mux_11754(v_260);
  assign v_11755 = mux_11755(v_254);
  assign v_11756 = mux_11756(v_5472);
  assign v_11758 = v_11759 | v_11761;
  assign v_11759 = mux_11759(v_11760);
  assign v_11760 = ~act_5429;
  assign v_11761 = v_11762 | v_11770;
  assign v_11762 = mux_11762(v_5430);
  assign v_11764 = v_11765 | v_11767;
  assign v_11765 = mux_11765(v_11766);
  assign v_11766 = ~act_5453;
  assign v_11767 = v_11768 | v_11769;
  assign v_11768 = mux_11768(v_246);
  assign v_11769 = mux_11769(v_240);
  assign v_11770 = mux_11770(v_5443);
  assign v_11772 = v_11773 | v_11775;
  assign v_11773 = mux_11773(v_11774);
  assign v_11774 = ~act_5436;
  assign v_11775 = v_11776 | v_11777;
  assign v_11776 = mux_11776(v_232);
  assign v_11777 = mux_11777(v_226);
  assign v_11778 = mux_11778(v_5377);
  assign v_11780 = v_11781 | v_11783;
  assign v_11781 = mux_11781(v_11782);
  assign v_11782 = ~act_2814;
  assign v_11783 = v_11784 | v_12338;
  assign v_11784 = mux_11784(v_2815);
  assign v_11786 = v_11787 | v_11789;
  assign v_11787 = mux_11787(v_11788);
  assign v_11788 = ~act_3954;
  assign v_11789 = v_11790 | v_12120;
  assign v_11790 = mux_11790(v_3955);
  assign v_11792 = v_11793 | v_11795;
  assign v_11793 = mux_11793(v_11794);
  assign v_11794 = ~act_4518;
  assign v_11795 = v_11796 | v_12014;
  assign v_11796 = mux_11796(v_4519);
  assign v_11798 = v_11799 | v_11801;
  assign v_11799 = mux_11799(v_11800);
  assign v_11800 = ~act_4794;
  assign v_11801 = v_11802 | v_11908;
  assign v_11802 = mux_11802(v_4795);
  assign v_11804 = v_11805 | v_11807;
  assign v_11805 = mux_11805(v_11806);
  assign v_11806 = ~act_5070;
  assign v_11807 = v_11808 | v_11858;
  assign v_11808 = mux_11808(v_5071);
  assign v_11810 = v_11811 | v_11813;
  assign v_11811 = mux_11811(v_11812);
  assign v_11812 = ~act_5202;
  assign v_11813 = v_11814 | v_11836;
  assign v_11814 = mux_11814(v_5203);
  assign v_11816 = v_11817 | v_11819;
  assign v_11817 = mux_11817(v_11818);
  assign v_11818 = ~act_5262;
  assign v_11819 = v_11820 | v_11828;
  assign v_11820 = mux_11820(v_5263);
  assign v_11822 = v_11823 | v_11825;
  assign v_11823 = mux_11823(v_11824);
  assign v_11824 = ~act_5286;
  assign v_11825 = v_11826 | v_11827;
  assign v_11826 = mux_11826(v_218);
  assign v_11827 = mux_11827(v_212);
  assign v_11828 = mux_11828(v_5276);
  assign v_11830 = v_11831 | v_11833;
  assign v_11831 = mux_11831(v_11832);
  assign v_11832 = ~act_5269;
  assign v_11833 = v_11834 | v_11835;
  assign v_11834 = mux_11834(v_204);
  assign v_11835 = mux_11835(v_198);
  assign v_11836 = mux_11836(v_5252);
  assign v_11838 = v_11839 | v_11841;
  assign v_11839 = mux_11839(v_11840);
  assign v_11840 = ~act_5209;
  assign v_11841 = v_11842 | v_11850;
  assign v_11842 = mux_11842(v_5210);
  assign v_11844 = v_11845 | v_11847;
  assign v_11845 = mux_11845(v_11846);
  assign v_11846 = ~act_5233;
  assign v_11847 = v_11848 | v_11849;
  assign v_11848 = mux_11848(v_190);
  assign v_11849 = mux_11849(v_184);
  assign v_11850 = mux_11850(v_5223);
  assign v_11852 = v_11853 | v_11855;
  assign v_11853 = mux_11853(v_11854);
  assign v_11854 = ~act_5216;
  assign v_11855 = v_11856 | v_11857;
  assign v_11856 = mux_11856(v_176);
  assign v_11857 = mux_11857(v_170);
  assign v_11858 = mux_11858(v_5192);
  assign v_11860 = v_11861 | v_11863;
  assign v_11861 = mux_11861(v_11862);
  assign v_11862 = ~act_5077;
  assign v_11863 = v_11864 | v_11886;
  assign v_11864 = mux_11864(v_5078);
  assign v_11866 = v_11867 | v_11869;
  assign v_11867 = mux_11867(v_11868);
  assign v_11868 = ~act_5137;
  assign v_11869 = v_11870 | v_11878;
  assign v_11870 = mux_11870(v_5138);
  assign v_11872 = v_11873 | v_11875;
  assign v_11873 = mux_11873(v_11874);
  assign v_11874 = ~act_5161;
  assign v_11875 = v_11876 | v_11877;
  assign v_11876 = mux_11876(v_162);
  assign v_11877 = mux_11877(v_156);
  assign v_11878 = mux_11878(v_5151);
  assign v_11880 = v_11881 | v_11883;
  assign v_11881 = mux_11881(v_11882);
  assign v_11882 = ~act_5144;
  assign v_11883 = v_11884 | v_11885;
  assign v_11884 = mux_11884(v_148);
  assign v_11885 = mux_11885(v_142);
  assign v_11886 = mux_11886(v_5127);
  assign v_11888 = v_11889 | v_11891;
  assign v_11889 = mux_11889(v_11890);
  assign v_11890 = ~act_5084;
  assign v_11891 = v_11892 | v_11900;
  assign v_11892 = mux_11892(v_5085);
  assign v_11894 = v_11895 | v_11897;
  assign v_11895 = mux_11895(v_11896);
  assign v_11896 = ~act_5108;
  assign v_11897 = v_11898 | v_11899;
  assign v_11898 = mux_11898(v_134);
  assign v_11899 = mux_11899(v_128);
  assign v_11900 = mux_11900(v_5098);
  assign v_11902 = v_11903 | v_11905;
  assign v_11903 = mux_11903(v_11904);
  assign v_11904 = ~act_5091;
  assign v_11905 = v_11906 | v_11907;
  assign v_11906 = mux_11906(v_120);
  assign v_11907 = mux_11907(v_114);
  assign v_11908 = mux_11908(v_5060);
  assign v_11910 = v_11911 | v_11913;
  assign v_11911 = mux_11911(v_11912);
  assign v_11912 = ~act_4801;
  assign v_11913 = v_11914 | v_11964;
  assign v_11914 = mux_11914(v_4802);
  assign v_11916 = v_11917 | v_11919;
  assign v_11917 = mux_11917(v_11918);
  assign v_11918 = ~act_4933;
  assign v_11919 = v_11920 | v_11942;
  assign v_11920 = mux_11920(v_4934);
  assign v_11922 = v_11923 | v_11925;
  assign v_11923 = mux_11923(v_11924);
  assign v_11924 = ~act_4993;
  assign v_11925 = v_11926 | v_11934;
  assign v_11926 = mux_11926(v_4994);
  assign v_11928 = v_11929 | v_11931;
  assign v_11929 = mux_11929(v_11930);
  assign v_11930 = ~act_5017;
  assign v_11931 = v_11932 | v_11933;
  assign v_11932 = mux_11932(v_106);
  assign v_11933 = mux_11933(v_100);
  assign v_11934 = mux_11934(v_5007);
  assign v_11936 = v_11937 | v_11939;
  assign v_11937 = mux_11937(v_11938);
  assign v_11938 = ~act_5000;
  assign v_11939 = v_11940 | v_11941;
  assign v_11940 = mux_11940(v_92);
  assign v_11941 = mux_11941(v_86);
  assign v_11942 = mux_11942(v_4983);
  assign v_11944 = v_11945 | v_11947;
  assign v_11945 = mux_11945(v_11946);
  assign v_11946 = ~act_4940;
  assign v_11947 = v_11948 | v_11956;
  assign v_11948 = mux_11948(v_4941);
  assign v_11950 = v_11951 | v_11953;
  assign v_11951 = mux_11951(v_11952);
  assign v_11952 = ~act_4964;
  assign v_11953 = v_11954 | v_11955;
  assign v_11954 = mux_11954(v_78);
  assign v_11955 = mux_11955(v_72);
  assign v_11956 = mux_11956(v_4954);
  assign v_11958 = v_11959 | v_11961;
  assign v_11959 = mux_11959(v_11960);
  assign v_11960 = ~act_4947;
  assign v_11961 = v_11962 | v_11963;
  assign v_11962 = mux_11962(v_64);
  assign v_11963 = mux_11963(v_58);
  assign v_11964 = mux_11964(v_4923);
  assign v_11966 = v_11967 | v_11969;
  assign v_11967 = mux_11967(v_11968);
  assign v_11968 = ~act_4808;
  assign v_11969 = v_11970 | v_11992;
  assign v_11970 = mux_11970(v_4809);
  assign v_11972 = v_11973 | v_11975;
  assign v_11973 = mux_11973(v_11974);
  assign v_11974 = ~act_4868;
  assign v_11975 = v_11976 | v_11984;
  assign v_11976 = mux_11976(v_4869);
  assign v_11978 = v_11979 | v_11981;
  assign v_11979 = mux_11979(v_11980);
  assign v_11980 = ~act_4892;
  assign v_11981 = v_11982 | v_11983;
  assign v_11982 = mux_11982(v_50);
  assign v_11983 = mux_11983(v_44);
  assign v_11984 = mux_11984(v_4882);
  assign v_11986 = v_11987 | v_11989;
  assign v_11987 = mux_11987(v_11988);
  assign v_11988 = ~act_4875;
  assign v_11989 = v_11990 | v_11991;
  assign v_11990 = mux_11990(v_36);
  assign v_11991 = mux_11991(v_30);
  assign v_11992 = mux_11992(v_4858);
  assign v_11994 = v_11995 | v_11997;
  assign v_11995 = mux_11995(v_11996);
  assign v_11996 = ~act_4815;
  assign v_11997 = v_11998 | v_12006;
  assign v_11998 = mux_11998(v_4816);
  assign v_12000 = v_12001 | v_12003;
  assign v_12001 = mux_12001(v_12002);
  assign v_12002 = ~act_4839;
  assign v_12003 = v_12004 | v_12005;
  assign v_12004 = mux_12004(v_22);
  assign v_12005 = mux_12005(v_16);
  assign v_12006 = mux_12006(v_4829);
  assign v_12008 = v_12009 | v_12011;
  assign v_12009 = mux_12009(v_12010);
  assign v_12010 = ~act_4822;
  assign v_12011 = v_12012 | v_12013;
  assign v_12012 = mux_12012(v_8);
  assign v_12013 = mux_12013(v_2);
  assign v_12014 = mux_12014(v_4784);
  assign v_12016 = v_12017 | v_12019;
  assign v_12017 = mux_12017(v_12018);
  assign v_12018 = ~act_4525;
  assign v_12019 = v_12020 | v_12070;
  assign v_12020 = mux_12020(v_4526);
  assign v_12022 = v_12023 | v_12025;
  assign v_12023 = mux_12023(v_12024);
  assign v_12024 = ~act_4657;
  assign v_12025 = v_12026 | v_12048;
  assign v_12026 = mux_12026(v_4658);
  assign v_12028 = v_12029 | v_12031;
  assign v_12029 = mux_12029(v_12030);
  assign v_12030 = ~act_4717;
  assign v_12031 = v_12032 | v_12040;
  assign v_12032 = mux_12032(v_4718);
  assign v_12034 = v_12035 | v_12037;
  assign v_12035 = mux_12035(v_12036);
  assign v_12036 = ~act_4741;
  assign v_12037 = v_12038 | v_12039;
  assign v_12038 = mux_12038(v_2794);
  assign v_12039 = mux_12039(v_2788);
  assign v_12040 = mux_12040(v_4731);
  assign v_12042 = v_12043 | v_12045;
  assign v_12043 = mux_12043(v_12044);
  assign v_12044 = ~act_4724;
  assign v_12045 = v_12046 | v_12047;
  assign v_12046 = mux_12046(v_2780);
  assign v_12047 = mux_12047(v_2774);
  assign v_12048 = mux_12048(v_4707);
  assign v_12050 = v_12051 | v_12053;
  assign v_12051 = mux_12051(v_12052);
  assign v_12052 = ~act_4664;
  assign v_12053 = v_12054 | v_12062;
  assign v_12054 = mux_12054(v_4665);
  assign v_12056 = v_12057 | v_12059;
  assign v_12057 = mux_12057(v_12058);
  assign v_12058 = ~act_4688;
  assign v_12059 = v_12060 | v_12061;
  assign v_12060 = mux_12060(v_2766);
  assign v_12061 = mux_12061(v_2760);
  assign v_12062 = mux_12062(v_4678);
  assign v_12064 = v_12065 | v_12067;
  assign v_12065 = mux_12065(v_12066);
  assign v_12066 = ~act_4671;
  assign v_12067 = v_12068 | v_12069;
  assign v_12068 = mux_12068(v_2752);
  assign v_12069 = mux_12069(v_2746);
  assign v_12070 = mux_12070(v_4647);
  assign v_12072 = v_12073 | v_12075;
  assign v_12073 = mux_12073(v_12074);
  assign v_12074 = ~act_4532;
  assign v_12075 = v_12076 | v_12098;
  assign v_12076 = mux_12076(v_4533);
  assign v_12078 = v_12079 | v_12081;
  assign v_12079 = mux_12079(v_12080);
  assign v_12080 = ~act_4592;
  assign v_12081 = v_12082 | v_12090;
  assign v_12082 = mux_12082(v_4593);
  assign v_12084 = v_12085 | v_12087;
  assign v_12085 = mux_12085(v_12086);
  assign v_12086 = ~act_4616;
  assign v_12087 = v_12088 | v_12089;
  assign v_12088 = mux_12088(v_2738);
  assign v_12089 = mux_12089(v_2732);
  assign v_12090 = mux_12090(v_4606);
  assign v_12092 = v_12093 | v_12095;
  assign v_12093 = mux_12093(v_12094);
  assign v_12094 = ~act_4599;
  assign v_12095 = v_12096 | v_12097;
  assign v_12096 = mux_12096(v_2724);
  assign v_12097 = mux_12097(v_2718);
  assign v_12098 = mux_12098(v_4582);
  assign v_12100 = v_12101 | v_12103;
  assign v_12101 = mux_12101(v_12102);
  assign v_12102 = ~act_4539;
  assign v_12103 = v_12104 | v_12112;
  assign v_12104 = mux_12104(v_4540);
  assign v_12106 = v_12107 | v_12109;
  assign v_12107 = mux_12107(v_12108);
  assign v_12108 = ~act_4563;
  assign v_12109 = v_12110 | v_12111;
  assign v_12110 = mux_12110(v_2710);
  assign v_12111 = mux_12111(v_2704);
  assign v_12112 = mux_12112(v_4553);
  assign v_12114 = v_12115 | v_12117;
  assign v_12115 = mux_12115(v_12116);
  assign v_12116 = ~act_4546;
  assign v_12117 = v_12118 | v_12119;
  assign v_12118 = mux_12118(v_2696);
  assign v_12119 = mux_12119(v_2690);
  assign v_12120 = mux_12120(v_4508);
  assign v_12122 = v_12123 | v_12125;
  assign v_12123 = mux_12123(v_12124);
  assign v_12124 = ~act_3961;
  assign v_12125 = v_12126 | v_12232;
  assign v_12126 = mux_12126(v_3962);
  assign v_12128 = v_12129 | v_12131;
  assign v_12129 = mux_12129(v_12130);
  assign v_12130 = ~act_4237;
  assign v_12131 = v_12132 | v_12182;
  assign v_12132 = mux_12132(v_4238);
  assign v_12134 = v_12135 | v_12137;
  assign v_12135 = mux_12135(v_12136);
  assign v_12136 = ~act_4369;
  assign v_12137 = v_12138 | v_12160;
  assign v_12138 = mux_12138(v_4370);
  assign v_12140 = v_12141 | v_12143;
  assign v_12141 = mux_12141(v_12142);
  assign v_12142 = ~act_4429;
  assign v_12143 = v_12144 | v_12152;
  assign v_12144 = mux_12144(v_4430);
  assign v_12146 = v_12147 | v_12149;
  assign v_12147 = mux_12147(v_12148);
  assign v_12148 = ~act_4453;
  assign v_12149 = v_12150 | v_12151;
  assign v_12150 = mux_12150(v_2682);
  assign v_12151 = mux_12151(v_2676);
  assign v_12152 = mux_12152(v_4443);
  assign v_12154 = v_12155 | v_12157;
  assign v_12155 = mux_12155(v_12156);
  assign v_12156 = ~act_4436;
  assign v_12157 = v_12158 | v_12159;
  assign v_12158 = mux_12158(v_2668);
  assign v_12159 = mux_12159(v_2662);
  assign v_12160 = mux_12160(v_4419);
  assign v_12162 = v_12163 | v_12165;
  assign v_12163 = mux_12163(v_12164);
  assign v_12164 = ~act_4376;
  assign v_12165 = v_12166 | v_12174;
  assign v_12166 = mux_12166(v_4377);
  assign v_12168 = v_12169 | v_12171;
  assign v_12169 = mux_12169(v_12170);
  assign v_12170 = ~act_4400;
  assign v_12171 = v_12172 | v_12173;
  assign v_12172 = mux_12172(v_2654);
  assign v_12173 = mux_12173(v_2648);
  assign v_12174 = mux_12174(v_4390);
  assign v_12176 = v_12177 | v_12179;
  assign v_12177 = mux_12177(v_12178);
  assign v_12178 = ~act_4383;
  assign v_12179 = v_12180 | v_12181;
  assign v_12180 = mux_12180(v_2640);
  assign v_12181 = mux_12181(v_2634);
  assign v_12182 = mux_12182(v_4359);
  assign v_12184 = v_12185 | v_12187;
  assign v_12185 = mux_12185(v_12186);
  assign v_12186 = ~act_4244;
  assign v_12187 = v_12188 | v_12210;
  assign v_12188 = mux_12188(v_4245);
  assign v_12190 = v_12191 | v_12193;
  assign v_12191 = mux_12191(v_12192);
  assign v_12192 = ~act_4304;
  assign v_12193 = v_12194 | v_12202;
  assign v_12194 = mux_12194(v_4305);
  assign v_12196 = v_12197 | v_12199;
  assign v_12197 = mux_12197(v_12198);
  assign v_12198 = ~act_4328;
  assign v_12199 = v_12200 | v_12201;
  assign v_12200 = mux_12200(v_2626);
  assign v_12201 = mux_12201(v_2620);
  assign v_12202 = mux_12202(v_4318);
  assign v_12204 = v_12205 | v_12207;
  assign v_12205 = mux_12205(v_12206);
  assign v_12206 = ~act_4311;
  assign v_12207 = v_12208 | v_12209;
  assign v_12208 = mux_12208(v_2612);
  assign v_12209 = mux_12209(v_2606);
  assign v_12210 = mux_12210(v_4294);
  assign v_12212 = v_12213 | v_12215;
  assign v_12213 = mux_12213(v_12214);
  assign v_12214 = ~act_4251;
  assign v_12215 = v_12216 | v_12224;
  assign v_12216 = mux_12216(v_4252);
  assign v_12218 = v_12219 | v_12221;
  assign v_12219 = mux_12219(v_12220);
  assign v_12220 = ~act_4275;
  assign v_12221 = v_12222 | v_12223;
  assign v_12222 = mux_12222(v_2598);
  assign v_12223 = mux_12223(v_2592);
  assign v_12224 = mux_12224(v_4265);
  assign v_12226 = v_12227 | v_12229;
  assign v_12227 = mux_12227(v_12228);
  assign v_12228 = ~act_4258;
  assign v_12229 = v_12230 | v_12231;
  assign v_12230 = mux_12230(v_2584);
  assign v_12231 = mux_12231(v_2578);
  assign v_12232 = mux_12232(v_4227);
  assign v_12234 = v_12235 | v_12237;
  assign v_12235 = mux_12235(v_12236);
  assign v_12236 = ~act_3968;
  assign v_12237 = v_12238 | v_12288;
  assign v_12238 = mux_12238(v_3969);
  assign v_12240 = v_12241 | v_12243;
  assign v_12241 = mux_12241(v_12242);
  assign v_12242 = ~act_4100;
  assign v_12243 = v_12244 | v_12266;
  assign v_12244 = mux_12244(v_4101);
  assign v_12246 = v_12247 | v_12249;
  assign v_12247 = mux_12247(v_12248);
  assign v_12248 = ~act_4160;
  assign v_12249 = v_12250 | v_12258;
  assign v_12250 = mux_12250(v_4161);
  assign v_12252 = v_12253 | v_12255;
  assign v_12253 = mux_12253(v_12254);
  assign v_12254 = ~act_4184;
  assign v_12255 = v_12256 | v_12257;
  assign v_12256 = mux_12256(v_2570);
  assign v_12257 = mux_12257(v_2564);
  assign v_12258 = mux_12258(v_4174);
  assign v_12260 = v_12261 | v_12263;
  assign v_12261 = mux_12261(v_12262);
  assign v_12262 = ~act_4167;
  assign v_12263 = v_12264 | v_12265;
  assign v_12264 = mux_12264(v_2556);
  assign v_12265 = mux_12265(v_2550);
  assign v_12266 = mux_12266(v_4150);
  assign v_12268 = v_12269 | v_12271;
  assign v_12269 = mux_12269(v_12270);
  assign v_12270 = ~act_4107;
  assign v_12271 = v_12272 | v_12280;
  assign v_12272 = mux_12272(v_4108);
  assign v_12274 = v_12275 | v_12277;
  assign v_12275 = mux_12275(v_12276);
  assign v_12276 = ~act_4131;
  assign v_12277 = v_12278 | v_12279;
  assign v_12278 = mux_12278(v_2542);
  assign v_12279 = mux_12279(v_2536);
  assign v_12280 = mux_12280(v_4121);
  assign v_12282 = v_12283 | v_12285;
  assign v_12283 = mux_12283(v_12284);
  assign v_12284 = ~act_4114;
  assign v_12285 = v_12286 | v_12287;
  assign v_12286 = mux_12286(v_2528);
  assign v_12287 = mux_12287(v_2522);
  assign v_12288 = mux_12288(v_4090);
  assign v_12290 = v_12291 | v_12293;
  assign v_12291 = mux_12291(v_12292);
  assign v_12292 = ~act_3975;
  assign v_12293 = v_12294 | v_12316;
  assign v_12294 = mux_12294(v_3976);
  assign v_12296 = v_12297 | v_12299;
  assign v_12297 = mux_12297(v_12298);
  assign v_12298 = ~act_4035;
  assign v_12299 = v_12300 | v_12308;
  assign v_12300 = mux_12300(v_4036);
  assign v_12302 = v_12303 | v_12305;
  assign v_12303 = mux_12303(v_12304);
  assign v_12304 = ~act_4059;
  assign v_12305 = v_12306 | v_12307;
  assign v_12306 = mux_12306(v_2514);
  assign v_12307 = mux_12307(v_2508);
  assign v_12308 = mux_12308(v_4049);
  assign v_12310 = v_12311 | v_12313;
  assign v_12311 = mux_12311(v_12312);
  assign v_12312 = ~act_4042;
  assign v_12313 = v_12314 | v_12315;
  assign v_12314 = mux_12314(v_2500);
  assign v_12315 = mux_12315(v_2494);
  assign v_12316 = mux_12316(v_4025);
  assign v_12318 = v_12319 | v_12321;
  assign v_12319 = mux_12319(v_12320);
  assign v_12320 = ~act_3982;
  assign v_12321 = v_12322 | v_12330;
  assign v_12322 = mux_12322(v_3983);
  assign v_12324 = v_12325 | v_12327;
  assign v_12325 = mux_12325(v_12326);
  assign v_12326 = ~act_4006;
  assign v_12327 = v_12328 | v_12329;
  assign v_12328 = mux_12328(v_2486);
  assign v_12329 = mux_12329(v_2480);
  assign v_12330 = mux_12330(v_3996);
  assign v_12332 = v_12333 | v_12335;
  assign v_12333 = mux_12333(v_12334);
  assign v_12334 = ~act_3989;
  assign v_12335 = v_12336 | v_12337;
  assign v_12336 = mux_12336(v_2472);
  assign v_12337 = mux_12337(v_2466);
  assign v_12338 = mux_12338(v_3944);
  assign v_12340 = v_12341 | v_12343;
  assign v_12341 = mux_12341(v_12342);
  assign v_12342 = ~act_2821;
  assign v_12343 = v_12344 | v_12562;
  assign v_12344 = mux_12344(v_2822);
  assign v_12346 = v_12347 | v_12349;
  assign v_12347 = mux_12347(v_12348);
  assign v_12348 = ~act_3385;
  assign v_12349 = v_12350 | v_12456;
  assign v_12350 = mux_12350(v_3386);
  assign v_12352 = v_12353 | v_12355;
  assign v_12353 = mux_12353(v_12354);
  assign v_12354 = ~act_3661;
  assign v_12355 = v_12356 | v_12406;
  assign v_12356 = mux_12356(v_3662);
  assign v_12358 = v_12359 | v_12361;
  assign v_12359 = mux_12359(v_12360);
  assign v_12360 = ~act_3793;
  assign v_12361 = v_12362 | v_12384;
  assign v_12362 = mux_12362(v_3794);
  assign v_12364 = v_12365 | v_12367;
  assign v_12365 = mux_12365(v_12366);
  assign v_12366 = ~act_3853;
  assign v_12367 = v_12368 | v_12376;
  assign v_12368 = mux_12368(v_3854);
  assign v_12370 = v_12371 | v_12373;
  assign v_12371 = mux_12371(v_12372);
  assign v_12372 = ~act_3877;
  assign v_12373 = v_12374 | v_12375;
  assign v_12374 = mux_12374(v_2458);
  assign v_12375 = mux_12375(v_2452);
  assign v_12376 = mux_12376(v_3867);
  assign v_12378 = v_12379 | v_12381;
  assign v_12379 = mux_12379(v_12380);
  assign v_12380 = ~act_3860;
  assign v_12381 = v_12382 | v_12383;
  assign v_12382 = mux_12382(v_2444);
  assign v_12383 = mux_12383(v_2438);
  assign v_12384 = mux_12384(v_3843);
  assign v_12386 = v_12387 | v_12389;
  assign v_12387 = mux_12387(v_12388);
  assign v_12388 = ~act_3800;
  assign v_12389 = v_12390 | v_12398;
  assign v_12390 = mux_12390(v_3801);
  assign v_12392 = v_12393 | v_12395;
  assign v_12393 = mux_12393(v_12394);
  assign v_12394 = ~act_3824;
  assign v_12395 = v_12396 | v_12397;
  assign v_12396 = mux_12396(v_2430);
  assign v_12397 = mux_12397(v_2424);
  assign v_12398 = mux_12398(v_3814);
  assign v_12400 = v_12401 | v_12403;
  assign v_12401 = mux_12401(v_12402);
  assign v_12402 = ~act_3807;
  assign v_12403 = v_12404 | v_12405;
  assign v_12404 = mux_12404(v_2416);
  assign v_12405 = mux_12405(v_2410);
  assign v_12406 = mux_12406(v_3783);
  assign v_12408 = v_12409 | v_12411;
  assign v_12409 = mux_12409(v_12410);
  assign v_12410 = ~act_3668;
  assign v_12411 = v_12412 | v_12434;
  assign v_12412 = mux_12412(v_3669);
  assign v_12414 = v_12415 | v_12417;
  assign v_12415 = mux_12415(v_12416);
  assign v_12416 = ~act_3728;
  assign v_12417 = v_12418 | v_12426;
  assign v_12418 = mux_12418(v_3729);
  assign v_12420 = v_12421 | v_12423;
  assign v_12421 = mux_12421(v_12422);
  assign v_12422 = ~act_3752;
  assign v_12423 = v_12424 | v_12425;
  assign v_12424 = mux_12424(v_2402);
  assign v_12425 = mux_12425(v_2396);
  assign v_12426 = mux_12426(v_3742);
  assign v_12428 = v_12429 | v_12431;
  assign v_12429 = mux_12429(v_12430);
  assign v_12430 = ~act_3735;
  assign v_12431 = v_12432 | v_12433;
  assign v_12432 = mux_12432(v_2388);
  assign v_12433 = mux_12433(v_2382);
  assign v_12434 = mux_12434(v_3718);
  assign v_12436 = v_12437 | v_12439;
  assign v_12437 = mux_12437(v_12438);
  assign v_12438 = ~act_3675;
  assign v_12439 = v_12440 | v_12448;
  assign v_12440 = mux_12440(v_3676);
  assign v_12442 = v_12443 | v_12445;
  assign v_12443 = mux_12443(v_12444);
  assign v_12444 = ~act_3699;
  assign v_12445 = v_12446 | v_12447;
  assign v_12446 = mux_12446(v_2374);
  assign v_12447 = mux_12447(v_2368);
  assign v_12448 = mux_12448(v_3689);
  assign v_12450 = v_12451 | v_12453;
  assign v_12451 = mux_12451(v_12452);
  assign v_12452 = ~act_3682;
  assign v_12453 = v_12454 | v_12455;
  assign v_12454 = mux_12454(v_2360);
  assign v_12455 = mux_12455(v_2354);
  assign v_12456 = mux_12456(v_3651);
  assign v_12458 = v_12459 | v_12461;
  assign v_12459 = mux_12459(v_12460);
  assign v_12460 = ~act_3392;
  assign v_12461 = v_12462 | v_12512;
  assign v_12462 = mux_12462(v_3393);
  assign v_12464 = v_12465 | v_12467;
  assign v_12465 = mux_12465(v_12466);
  assign v_12466 = ~act_3524;
  assign v_12467 = v_12468 | v_12490;
  assign v_12468 = mux_12468(v_3525);
  assign v_12470 = v_12471 | v_12473;
  assign v_12471 = mux_12471(v_12472);
  assign v_12472 = ~act_3584;
  assign v_12473 = v_12474 | v_12482;
  assign v_12474 = mux_12474(v_3585);
  assign v_12476 = v_12477 | v_12479;
  assign v_12477 = mux_12477(v_12478);
  assign v_12478 = ~act_3608;
  assign v_12479 = v_12480 | v_12481;
  assign v_12480 = mux_12480(v_2346);
  assign v_12481 = mux_12481(v_2340);
  assign v_12482 = mux_12482(v_3598);
  assign v_12484 = v_12485 | v_12487;
  assign v_12485 = mux_12485(v_12486);
  assign v_12486 = ~act_3591;
  assign v_12487 = v_12488 | v_12489;
  assign v_12488 = mux_12488(v_2332);
  assign v_12489 = mux_12489(v_2326);
  assign v_12490 = mux_12490(v_3574);
  assign v_12492 = v_12493 | v_12495;
  assign v_12493 = mux_12493(v_12494);
  assign v_12494 = ~act_3531;
  assign v_12495 = v_12496 | v_12504;
  assign v_12496 = mux_12496(v_3532);
  assign v_12498 = v_12499 | v_12501;
  assign v_12499 = mux_12499(v_12500);
  assign v_12500 = ~act_3555;
  assign v_12501 = v_12502 | v_12503;
  assign v_12502 = mux_12502(v_2318);
  assign v_12503 = mux_12503(v_2312);
  assign v_12504 = mux_12504(v_3545);
  assign v_12506 = v_12507 | v_12509;
  assign v_12507 = mux_12507(v_12508);
  assign v_12508 = ~act_3538;
  assign v_12509 = v_12510 | v_12511;
  assign v_12510 = mux_12510(v_2304);
  assign v_12511 = mux_12511(v_2298);
  assign v_12512 = mux_12512(v_3514);
  assign v_12514 = v_12515 | v_12517;
  assign v_12515 = mux_12515(v_12516);
  assign v_12516 = ~act_3399;
  assign v_12517 = v_12518 | v_12540;
  assign v_12518 = mux_12518(v_3400);
  assign v_12520 = v_12521 | v_12523;
  assign v_12521 = mux_12521(v_12522);
  assign v_12522 = ~act_3459;
  assign v_12523 = v_12524 | v_12532;
  assign v_12524 = mux_12524(v_3460);
  assign v_12526 = v_12527 | v_12529;
  assign v_12527 = mux_12527(v_12528);
  assign v_12528 = ~act_3483;
  assign v_12529 = v_12530 | v_12531;
  assign v_12530 = mux_12530(v_2290);
  assign v_12531 = mux_12531(v_2284);
  assign v_12532 = mux_12532(v_3473);
  assign v_12534 = v_12535 | v_12537;
  assign v_12535 = mux_12535(v_12536);
  assign v_12536 = ~act_3466;
  assign v_12537 = v_12538 | v_12539;
  assign v_12538 = mux_12538(v_2276);
  assign v_12539 = mux_12539(v_2270);
  assign v_12540 = mux_12540(v_3449);
  assign v_12542 = v_12543 | v_12545;
  assign v_12543 = mux_12543(v_12544);
  assign v_12544 = ~act_3406;
  assign v_12545 = v_12546 | v_12554;
  assign v_12546 = mux_12546(v_3407);
  assign v_12548 = v_12549 | v_12551;
  assign v_12549 = mux_12549(v_12550);
  assign v_12550 = ~act_3430;
  assign v_12551 = v_12552 | v_12553;
  assign v_12552 = mux_12552(v_2262);
  assign v_12553 = mux_12553(v_2256);
  assign v_12554 = mux_12554(v_3420);
  assign v_12556 = v_12557 | v_12559;
  assign v_12557 = mux_12557(v_12558);
  assign v_12558 = ~act_3413;
  assign v_12559 = v_12560 | v_12561;
  assign v_12560 = mux_12560(v_2248);
  assign v_12561 = mux_12561(v_2242);
  assign v_12562 = mux_12562(v_3375);
  assign v_12564 = v_12565 | v_12567;
  assign v_12565 = mux_12565(v_12566);
  assign v_12566 = ~act_2828;
  assign v_12567 = v_12568 | v_12674;
  assign v_12568 = mux_12568(v_2829);
  assign v_12570 = v_12571 | v_12573;
  assign v_12571 = mux_12571(v_12572);
  assign v_12572 = ~act_3104;
  assign v_12573 = v_12574 | v_12624;
  assign v_12574 = mux_12574(v_3105);
  assign v_12576 = v_12577 | v_12579;
  assign v_12577 = mux_12577(v_12578);
  assign v_12578 = ~act_3236;
  assign v_12579 = v_12580 | v_12602;
  assign v_12580 = mux_12580(v_3237);
  assign v_12582 = v_12583 | v_12585;
  assign v_12583 = mux_12583(v_12584);
  assign v_12584 = ~act_3296;
  assign v_12585 = v_12586 | v_12594;
  assign v_12586 = mux_12586(v_3297);
  assign v_12588 = v_12589 | v_12591;
  assign v_12589 = mux_12589(v_12590);
  assign v_12590 = ~act_3320;
  assign v_12591 = v_12592 | v_12593;
  assign v_12592 = mux_12592(v_2234);
  assign v_12593 = mux_12593(v_2228);
  assign v_12594 = mux_12594(v_3310);
  assign v_12596 = v_12597 | v_12599;
  assign v_12597 = mux_12597(v_12598);
  assign v_12598 = ~act_3303;
  assign v_12599 = v_12600 | v_12601;
  assign v_12600 = mux_12600(v_2220);
  assign v_12601 = mux_12601(v_2214);
  assign v_12602 = mux_12602(v_3286);
  assign v_12604 = v_12605 | v_12607;
  assign v_12605 = mux_12605(v_12606);
  assign v_12606 = ~act_3243;
  assign v_12607 = v_12608 | v_12616;
  assign v_12608 = mux_12608(v_3244);
  assign v_12610 = v_12611 | v_12613;
  assign v_12611 = mux_12611(v_12612);
  assign v_12612 = ~act_3267;
  assign v_12613 = v_12614 | v_12615;
  assign v_12614 = mux_12614(v_2206);
  assign v_12615 = mux_12615(v_2200);
  assign v_12616 = mux_12616(v_3257);
  assign v_12618 = v_12619 | v_12621;
  assign v_12619 = mux_12619(v_12620);
  assign v_12620 = ~act_3250;
  assign v_12621 = v_12622 | v_12623;
  assign v_12622 = mux_12622(v_2192);
  assign v_12623 = mux_12623(v_2186);
  assign v_12624 = mux_12624(v_3226);
  assign v_12626 = v_12627 | v_12629;
  assign v_12627 = mux_12627(v_12628);
  assign v_12628 = ~act_3111;
  assign v_12629 = v_12630 | v_12652;
  assign v_12630 = mux_12630(v_3112);
  assign v_12632 = v_12633 | v_12635;
  assign v_12633 = mux_12633(v_12634);
  assign v_12634 = ~act_3171;
  assign v_12635 = v_12636 | v_12644;
  assign v_12636 = mux_12636(v_3172);
  assign v_12638 = v_12639 | v_12641;
  assign v_12639 = mux_12639(v_12640);
  assign v_12640 = ~act_3195;
  assign v_12641 = v_12642 | v_12643;
  assign v_12642 = mux_12642(v_2178);
  assign v_12643 = mux_12643(v_2172);
  assign v_12644 = mux_12644(v_3185);
  assign v_12646 = v_12647 | v_12649;
  assign v_12647 = mux_12647(v_12648);
  assign v_12648 = ~act_3178;
  assign v_12649 = v_12650 | v_12651;
  assign v_12650 = mux_12650(v_2164);
  assign v_12651 = mux_12651(v_2158);
  assign v_12652 = mux_12652(v_3161);
  assign v_12654 = v_12655 | v_12657;
  assign v_12655 = mux_12655(v_12656);
  assign v_12656 = ~act_3118;
  assign v_12657 = v_12658 | v_12666;
  assign v_12658 = mux_12658(v_3119);
  assign v_12660 = v_12661 | v_12663;
  assign v_12661 = mux_12661(v_12662);
  assign v_12662 = ~act_3142;
  assign v_12663 = v_12664 | v_12665;
  assign v_12664 = mux_12664(v_2150);
  assign v_12665 = mux_12665(v_2144);
  assign v_12666 = mux_12666(v_3132);
  assign v_12668 = v_12669 | v_12671;
  assign v_12669 = mux_12669(v_12670);
  assign v_12670 = ~act_3125;
  assign v_12671 = v_12672 | v_12673;
  assign v_12672 = mux_12672(v_2136);
  assign v_12673 = mux_12673(v_2130);
  assign v_12674 = mux_12674(v_3094);
  assign v_12676 = v_12677 | v_12679;
  assign v_12677 = mux_12677(v_12678);
  assign v_12678 = ~act_2835;
  assign v_12679 = v_12680 | v_12730;
  assign v_12680 = mux_12680(v_2836);
  assign v_12682 = v_12683 | v_12685;
  assign v_12683 = mux_12683(v_12684);
  assign v_12684 = ~act_2967;
  assign v_12685 = v_12686 | v_12708;
  assign v_12686 = mux_12686(v_2968);
  assign v_12688 = v_12689 | v_12691;
  assign v_12689 = mux_12689(v_12690);
  assign v_12690 = ~act_3027;
  assign v_12691 = v_12692 | v_12700;
  assign v_12692 = mux_12692(v_3028);
  assign v_12694 = v_12695 | v_12697;
  assign v_12695 = mux_12695(v_12696);
  assign v_12696 = ~act_3051;
  assign v_12697 = v_12698 | v_12699;
  assign v_12698 = mux_12698(v_2122);
  assign v_12699 = mux_12699(v_2116);
  assign v_12700 = mux_12700(v_3041);
  assign v_12702 = v_12703 | v_12705;
  assign v_12703 = mux_12703(v_12704);
  assign v_12704 = ~act_3034;
  assign v_12705 = v_12706 | v_12707;
  assign v_12706 = mux_12706(v_2108);
  assign v_12707 = mux_12707(v_2102);
  assign v_12708 = mux_12708(v_3017);
  assign v_12710 = v_12711 | v_12713;
  assign v_12711 = mux_12711(v_12712);
  assign v_12712 = ~act_2974;
  assign v_12713 = v_12714 | v_12722;
  assign v_12714 = mux_12714(v_2975);
  assign v_12716 = v_12717 | v_12719;
  assign v_12717 = mux_12717(v_12718);
  assign v_12718 = ~act_2998;
  assign v_12719 = v_12720 | v_12721;
  assign v_12720 = mux_12720(v_2094);
  assign v_12721 = mux_12721(v_2088);
  assign v_12722 = mux_12722(v_2988);
  assign v_12724 = v_12725 | v_12727;
  assign v_12725 = mux_12725(v_12726);
  assign v_12726 = ~act_2981;
  assign v_12727 = v_12728 | v_12729;
  assign v_12728 = mux_12728(v_2080);
  assign v_12729 = mux_12729(v_2074);
  assign v_12730 = mux_12730(v_2957);
  assign v_12732 = v_12733 | v_12735;
  assign v_12733 = mux_12733(v_12734);
  assign v_12734 = ~act_2842;
  assign v_12735 = v_12736 | v_12758;
  assign v_12736 = mux_12736(v_2843);
  assign v_12738 = v_12739 | v_12741;
  assign v_12739 = mux_12739(v_12740);
  assign v_12740 = ~act_2902;
  assign v_12741 = v_12742 | v_12750;
  assign v_12742 = mux_12742(v_2903);
  assign v_12744 = v_12745 | v_12747;
  assign v_12745 = mux_12745(v_12746);
  assign v_12746 = ~act_2926;
  assign v_12747 = v_12748 | v_12749;
  assign v_12748 = mux_12748(v_2066);
  assign v_12749 = mux_12749(v_2060);
  assign v_12750 = mux_12750(v_2916);
  assign v_12752 = v_12753 | v_12755;
  assign v_12753 = mux_12753(v_12754);
  assign v_12754 = ~act_2909;
  assign v_12755 = v_12756 | v_12757;
  assign v_12756 = mux_12756(v_2052);
  assign v_12757 = mux_12757(v_2046);
  assign v_12758 = mux_12758(v_2892);
  assign v_12760 = v_12761 | v_12763;
  assign v_12761 = mux_12761(v_12762);
  assign v_12762 = ~act_2849;
  assign v_12763 = v_12764 | v_12772;
  assign v_12764 = mux_12764(v_2850);
  assign v_12766 = v_12767 | v_12769;
  assign v_12767 = mux_12767(v_12768);
  assign v_12768 = ~act_2873;
  assign v_12769 = v_12770 | v_12771;
  assign v_12770 = mux_12770(v_2038);
  assign v_12771 = mux_12771(v_2032);
  assign v_12772 = mux_12772(v_2863);
  assign v_12774 = v_12775 | v_12777;
  assign v_12775 = mux_12775(v_12776);
  assign v_12776 = ~act_2856;
  assign v_12777 = v_12778 | v_12779;
  assign v_12778 = mux_12778(v_2024);
  assign v_12779 = mux_12779(v_2018);
  assign v_12780 = in0_canPeek;
  assign v_12781 = in0_peek;
  // Always block
  //////////////////////////////////////////////////////////////////////////////
  always @(posedge clock) begin
    if (reset) begin
      v_2804 <= 1'h0;
      v_2811 <= 1'h0;
      v_2818 <= 1'h0;
      v_2825 <= 1'h0;
      v_2832 <= 1'h0;
      v_2839 <= 1'h0;
      v_2846 <= 1'h0;
      v_2853 <= 1'h0;
      v_2870 <= 1'h0;
      v_2899 <= 1'h0;
      v_2906 <= 1'h0;
      v_2923 <= 1'h0;
      v_2964 <= 1'h0;
      v_2971 <= 1'h0;
      v_2978 <= 1'h0;
      v_2995 <= 1'h0;
      v_3024 <= 1'h0;
      v_3031 <= 1'h0;
      v_3048 <= 1'h0;
      v_3101 <= 1'h0;
      v_3108 <= 1'h0;
      v_3115 <= 1'h0;
      v_3122 <= 1'h0;
      v_3139 <= 1'h0;
      v_3168 <= 1'h0;
      v_3175 <= 1'h0;
      v_3192 <= 1'h0;
      v_3233 <= 1'h0;
      v_3240 <= 1'h0;
      v_3247 <= 1'h0;
      v_3264 <= 1'h0;
      v_3293 <= 1'h0;
      v_3300 <= 1'h0;
      v_3317 <= 1'h0;
      v_3382 <= 1'h0;
      v_3389 <= 1'h0;
      v_3396 <= 1'h0;
      v_3403 <= 1'h0;
      v_3410 <= 1'h0;
      v_3427 <= 1'h0;
      v_3456 <= 1'h0;
      v_3463 <= 1'h0;
      v_3480 <= 1'h0;
      v_3521 <= 1'h0;
      v_3528 <= 1'h0;
      v_3535 <= 1'h0;
      v_3552 <= 1'h0;
      v_3581 <= 1'h0;
      v_3588 <= 1'h0;
      v_3605 <= 1'h0;
      v_3658 <= 1'h0;
      v_3665 <= 1'h0;
      v_3672 <= 1'h0;
      v_3679 <= 1'h0;
      v_3696 <= 1'h0;
      v_3725 <= 1'h0;
      v_3732 <= 1'h0;
      v_3749 <= 1'h0;
      v_3790 <= 1'h0;
      v_3797 <= 1'h0;
      v_3804 <= 1'h0;
      v_3821 <= 1'h0;
      v_3850 <= 1'h0;
      v_3857 <= 1'h0;
      v_3874 <= 1'h0;
      v_3951 <= 1'h0;
      v_3958 <= 1'h0;
      v_3965 <= 1'h0;
      v_3972 <= 1'h0;
      v_3979 <= 1'h0;
      v_3986 <= 1'h0;
      v_4003 <= 1'h0;
      v_4032 <= 1'h0;
      v_4039 <= 1'h0;
      v_4056 <= 1'h0;
      v_4097 <= 1'h0;
      v_4104 <= 1'h0;
      v_4111 <= 1'h0;
      v_4128 <= 1'h0;
      v_4157 <= 1'h0;
      v_4164 <= 1'h0;
      v_4181 <= 1'h0;
      v_4234 <= 1'h0;
      v_4241 <= 1'h0;
      v_4248 <= 1'h0;
      v_4255 <= 1'h0;
      v_4272 <= 1'h0;
      v_4301 <= 1'h0;
      v_4308 <= 1'h0;
      v_4325 <= 1'h0;
      v_4366 <= 1'h0;
      v_4373 <= 1'h0;
      v_4380 <= 1'h0;
      v_4397 <= 1'h0;
      v_4426 <= 1'h0;
      v_4433 <= 1'h0;
      v_4450 <= 1'h0;
      v_4515 <= 1'h0;
      v_4522 <= 1'h0;
      v_4529 <= 1'h0;
      v_4536 <= 1'h0;
      v_4543 <= 1'h0;
      v_4560 <= 1'h0;
      v_4589 <= 1'h0;
      v_4596 <= 1'h0;
      v_4613 <= 1'h0;
      v_4654 <= 1'h0;
      v_4661 <= 1'h0;
      v_4668 <= 1'h0;
      v_4685 <= 1'h0;
      v_4714 <= 1'h0;
      v_4721 <= 1'h0;
      v_4738 <= 1'h0;
      v_4791 <= 1'h0;
      v_4798 <= 1'h0;
      v_4805 <= 1'h0;
      v_4812 <= 1'h0;
      v_4819 <= 1'h0;
      v_4836 <= 1'h0;
      v_4865 <= 1'h0;
      v_4872 <= 1'h0;
      v_4889 <= 1'h0;
      v_4930 <= 1'h0;
      v_4937 <= 1'h0;
      v_4944 <= 1'h0;
      v_4961 <= 1'h0;
      v_4990 <= 1'h0;
      v_4997 <= 1'h0;
      v_5014 <= 1'h0;
      v_5067 <= 1'h0;
      v_5074 <= 1'h0;
      v_5081 <= 1'h0;
      v_5088 <= 1'h0;
      v_5105 <= 1'h0;
      v_5134 <= 1'h0;
      v_5141 <= 1'h0;
      v_5158 <= 1'h0;
      v_5199 <= 1'h0;
      v_5206 <= 1'h0;
      v_5213 <= 1'h0;
      v_5230 <= 1'h0;
      v_5259 <= 1'h0;
      v_5266 <= 1'h0;
      v_5283 <= 1'h0;
      v_5384 <= 1'h0;
      v_5391 <= 1'h0;
      v_5398 <= 1'h0;
      v_5405 <= 1'h0;
      v_5412 <= 1'h0;
      v_5419 <= 1'h0;
      v_5426 <= 1'h0;
      v_5433 <= 1'h0;
      v_5450 <= 1'h0;
      v_5479 <= 1'h0;
      v_5486 <= 1'h0;
      v_5503 <= 1'h0;
      v_5544 <= 1'h0;
      v_5551 <= 1'h0;
      v_5558 <= 1'h0;
      v_5575 <= 1'h0;
      v_5604 <= 1'h0;
      v_5611 <= 1'h0;
      v_5628 <= 1'h0;
      v_5681 <= 1'h0;
      v_5688 <= 1'h0;
      v_5695 <= 1'h0;
      v_5702 <= 1'h0;
      v_5719 <= 1'h0;
      v_5748 <= 1'h0;
      v_5755 <= 1'h0;
      v_5772 <= 1'h0;
      v_5813 <= 1'h0;
      v_5820 <= 1'h0;
      v_5827 <= 1'h0;
      v_5844 <= 1'h0;
      v_5873 <= 1'h0;
      v_5880 <= 1'h0;
      v_5897 <= 1'h0;
      v_5962 <= 1'h0;
      v_5969 <= 1'h0;
      v_5976 <= 1'h0;
      v_5983 <= 1'h0;
      v_5990 <= 1'h0;
      v_6007 <= 1'h0;
      v_6036 <= 1'h0;
      v_6043 <= 1'h0;
      v_6060 <= 1'h0;
      v_6101 <= 1'h0;
      v_6108 <= 1'h0;
      v_6115 <= 1'h0;
      v_6132 <= 1'h0;
      v_6161 <= 1'h0;
      v_6168 <= 1'h0;
      v_6185 <= 1'h0;
      v_6238 <= 1'h0;
      v_6245 <= 1'h0;
      v_6252 <= 1'h0;
      v_6259 <= 1'h0;
      v_6276 <= 1'h0;
      v_6305 <= 1'h0;
      v_6312 <= 1'h0;
      v_6329 <= 1'h0;
      v_6370 <= 1'h0;
      v_6377 <= 1'h0;
      v_6384 <= 1'h0;
      v_6401 <= 1'h0;
      v_6430 <= 1'h0;
      v_6437 <= 1'h0;
      v_6454 <= 1'h0;
      v_6531 <= 1'h0;
      v_6538 <= 1'h0;
      v_6545 <= 1'h0;
      v_6552 <= 1'h0;
      v_6559 <= 1'h0;
      v_6566 <= 1'h0;
      v_6583 <= 1'h0;
      v_6612 <= 1'h0;
      v_6619 <= 1'h0;
      v_6636 <= 1'h0;
      v_6677 <= 1'h0;
      v_6684 <= 1'h0;
      v_6691 <= 1'h0;
      v_6708 <= 1'h0;
      v_6737 <= 1'h0;
      v_6744 <= 1'h0;
      v_6761 <= 1'h0;
      v_6814 <= 1'h0;
      v_6821 <= 1'h0;
      v_6828 <= 1'h0;
      v_6835 <= 1'h0;
      v_6852 <= 1'h0;
      v_6881 <= 1'h0;
      v_6888 <= 1'h0;
      v_6905 <= 1'h0;
      v_6946 <= 1'h0;
      v_6953 <= 1'h0;
      v_6960 <= 1'h0;
      v_6977 <= 1'h0;
      v_7006 <= 1'h0;
      v_7013 <= 1'h0;
      v_7030 <= 1'h0;
      v_7095 <= 1'h0;
      v_7102 <= 1'h0;
      v_7109 <= 1'h0;
      v_7116 <= 1'h0;
      v_7123 <= 1'h0;
      v_7140 <= 1'h0;
      v_7169 <= 1'h0;
      v_7176 <= 1'h0;
      v_7193 <= 1'h0;
      v_7234 <= 1'h0;
      v_7241 <= 1'h0;
      v_7248 <= 1'h0;
      v_7265 <= 1'h0;
      v_7294 <= 1'h0;
      v_7301 <= 1'h0;
      v_7318 <= 1'h0;
      v_7371 <= 1'h0;
      v_7378 <= 1'h0;
      v_7385 <= 1'h0;
      v_7392 <= 1'h0;
      v_7409 <= 1'h0;
      v_7438 <= 1'h0;
      v_7445 <= 1'h0;
      v_7462 <= 1'h0;
      v_7503 <= 1'h0;
      v_7510 <= 1'h0;
      v_7517 <= 1'h0;
      v_7534 <= 1'h0;
      v_7563 <= 1'h0;
      v_7570 <= 1'h0;
      v_7587 <= 1'h0;
      v_7676 <= 1'h0;
      v_7683 <= 1'h0;
      v_7690 <= 1'h0;
      v_7697 <= 1'h0;
      v_7704 <= 1'h0;
      v_7711 <= 1'h0;
      v_7718 <= 1'h0;
      v_7735 <= 1'h0;
      v_7764 <= 1'h0;
      v_7771 <= 1'h0;
      v_7788 <= 1'h0;
      v_7829 <= 1'h0;
      v_7836 <= 1'h0;
      v_7843 <= 1'h0;
      v_7860 <= 1'h0;
      v_7889 <= 1'h0;
      v_7896 <= 1'h0;
      v_7913 <= 1'h0;
      v_7966 <= 1'h0;
      v_7973 <= 1'h0;
      v_7980 <= 1'h0;
      v_7987 <= 1'h0;
      v_8004 <= 1'h0;
      v_8033 <= 1'h0;
      v_8040 <= 1'h0;
      v_8057 <= 1'h0;
      v_8098 <= 1'h0;
      v_8105 <= 1'h0;
      v_8112 <= 1'h0;
      v_8129 <= 1'h0;
      v_8158 <= 1'h0;
      v_8165 <= 1'h0;
      v_8182 <= 1'h0;
      v_8247 <= 1'h0;
      v_8254 <= 1'h0;
      v_8261 <= 1'h0;
      v_8268 <= 1'h0;
      v_8275 <= 1'h0;
      v_8292 <= 1'h0;
      v_8321 <= 1'h0;
      v_8328 <= 1'h0;
      v_8345 <= 1'h0;
      v_8386 <= 1'h0;
      v_8393 <= 1'h0;
      v_8400 <= 1'h0;
      v_8417 <= 1'h0;
      v_8446 <= 1'h0;
      v_8453 <= 1'h0;
      v_8470 <= 1'h0;
      v_8523 <= 1'h0;
      v_8530 <= 1'h0;
      v_8537 <= 1'h0;
      v_8544 <= 1'h0;
      v_8561 <= 1'h0;
      v_8590 <= 1'h0;
      v_8597 <= 1'h0;
      v_8614 <= 1'h0;
      v_8655 <= 1'h0;
      v_8662 <= 1'h0;
      v_8669 <= 1'h0;
      v_8686 <= 1'h0;
      v_8715 <= 1'h0;
      v_8722 <= 1'h0;
      v_8739 <= 1'h0;
      v_8816 <= 1'h0;
      v_8823 <= 1'h0;
      v_8830 <= 1'h0;
      v_8837 <= 1'h0;
      v_8844 <= 1'h0;
      v_8851 <= 1'h0;
      v_8868 <= 1'h0;
      v_8897 <= 1'h0;
      v_8904 <= 1'h0;
      v_8921 <= 1'h0;
      v_8962 <= 1'h0;
      v_8969 <= 1'h0;
      v_8976 <= 1'h0;
      v_8993 <= 1'h0;
      v_9022 <= 1'h0;
      v_9029 <= 1'h0;
      v_9046 <= 1'h0;
      v_9099 <= 1'h0;
      v_9106 <= 1'h0;
      v_9113 <= 1'h0;
      v_9120 <= 1'h0;
      v_9137 <= 1'h0;
      v_9166 <= 1'h0;
      v_9173 <= 1'h0;
      v_9190 <= 1'h0;
      v_9231 <= 1'h0;
      v_9238 <= 1'h0;
      v_9245 <= 1'h0;
      v_9262 <= 1'h0;
      v_9291 <= 1'h0;
      v_9298 <= 1'h0;
      v_9315 <= 1'h0;
      v_9380 <= 1'h0;
      v_9387 <= 1'h0;
      v_9394 <= 1'h0;
      v_9401 <= 1'h0;
      v_9408 <= 1'h0;
      v_9425 <= 1'h0;
      v_9454 <= 1'h0;
      v_9461 <= 1'h0;
      v_9478 <= 1'h0;
      v_9519 <= 1'h0;
      v_9526 <= 1'h0;
      v_9533 <= 1'h0;
      v_9550 <= 1'h0;
      v_9579 <= 1'h0;
      v_9586 <= 1'h0;
      v_9603 <= 1'h0;
      v_9656 <= 1'h0;
      v_9663 <= 1'h0;
      v_9670 <= 1'h0;
      v_9677 <= 1'h0;
      v_9694 <= 1'h0;
      v_9723 <= 1'h0;
      v_9730 <= 1'h0;
      v_9747 <= 1'h0;
      v_9788 <= 1'h0;
      v_9795 <= 1'h0;
      v_9802 <= 1'h0;
      v_9819 <= 1'h0;
      v_9848 <= 1'h0;
      v_9855 <= 1'h0;
      v_9872 <= 1'h0;
      v_9987 <= 8'h0;
      v_9993 <= 8'h0;
      v_9999 <= 8'h0;
      v_10005 <= 8'h0;
      v_10011 <= 8'h0;
      v_10017 <= 8'h0;
      v_10023 <= 8'h0;
      v_10029 <= 8'h0;
      v_10035 <= 8'h0;
      v_10043 <= 8'h0;
      v_10051 <= 8'h0;
      v_10057 <= 8'h0;
      v_10065 <= 8'h0;
      v_10073 <= 8'h0;
      v_10079 <= 8'h0;
      v_10085 <= 8'h0;
      v_10093 <= 8'h0;
      v_10101 <= 8'h0;
      v_10107 <= 8'h0;
      v_10115 <= 8'h0;
      v_10123 <= 8'h0;
      v_10129 <= 8'h0;
      v_10135 <= 8'h0;
      v_10141 <= 8'h0;
      v_10149 <= 8'h0;
      v_10157 <= 8'h0;
      v_10163 <= 8'h0;
      v_10171 <= 8'h0;
      v_10179 <= 8'h0;
      v_10185 <= 8'h0;
      v_10191 <= 8'h0;
      v_10199 <= 8'h0;
      v_10207 <= 8'h0;
      v_10213 <= 8'h0;
      v_10221 <= 8'h0;
      v_10229 <= 8'h0;
      v_10235 <= 8'h0;
      v_10241 <= 8'h0;
      v_10247 <= 8'h0;
      v_10253 <= 8'h0;
      v_10261 <= 8'h0;
      v_10269 <= 8'h0;
      v_10275 <= 8'h0;
      v_10283 <= 8'h0;
      v_10291 <= 8'h0;
      v_10297 <= 8'h0;
      v_10303 <= 8'h0;
      v_10311 <= 8'h0;
      v_10319 <= 8'h0;
      v_10325 <= 8'h0;
      v_10333 <= 8'h0;
      v_10341 <= 8'h0;
      v_10347 <= 8'h0;
      v_10353 <= 8'h0;
      v_10359 <= 8'h0;
      v_10367 <= 8'h0;
      v_10375 <= 8'h0;
      v_10381 <= 8'h0;
      v_10389 <= 8'h0;
      v_10397 <= 8'h0;
      v_10403 <= 8'h0;
      v_10409 <= 8'h0;
      v_10417 <= 8'h0;
      v_10425 <= 8'h0;
      v_10431 <= 8'h0;
      v_10439 <= 8'h0;
      v_10447 <= 8'h0;
      v_10453 <= 8'h0;
      v_10459 <= 8'h0;
      v_10465 <= 8'h0;
      v_10471 <= 8'h0;
      v_10477 <= 8'h0;
      v_10485 <= 8'h0;
      v_10493 <= 8'h0;
      v_10499 <= 8'h0;
      v_10507 <= 8'h0;
      v_10515 <= 8'h0;
      v_10521 <= 8'h0;
      v_10527 <= 8'h0;
      v_10535 <= 8'h0;
      v_10543 <= 8'h0;
      v_10549 <= 8'h0;
      v_10557 <= 8'h0;
      v_10565 <= 8'h0;
      v_10571 <= 8'h0;
      v_10577 <= 8'h0;
      v_10583 <= 8'h0;
      v_10591 <= 8'h0;
      v_10599 <= 8'h0;
      v_10605 <= 8'h0;
      v_10613 <= 8'h0;
      v_10621 <= 8'h0;
      v_10627 <= 8'h0;
      v_10633 <= 8'h0;
      v_10641 <= 8'h0;
      v_10649 <= 8'h0;
      v_10655 <= 8'h0;
      v_10663 <= 8'h0;
      v_10671 <= 8'h0;
      v_10677 <= 8'h0;
      v_10683 <= 8'h0;
      v_10689 <= 8'h0;
      v_10695 <= 8'h0;
      v_10703 <= 8'h0;
      v_10711 <= 8'h0;
      v_10717 <= 8'h0;
      v_10725 <= 8'h0;
      v_10733 <= 8'h0;
      v_10739 <= 8'h0;
      v_10745 <= 8'h0;
      v_10753 <= 8'h0;
      v_10761 <= 8'h0;
      v_10767 <= 8'h0;
      v_10775 <= 8'h0;
      v_10783 <= 8'h0;
      v_10789 <= 8'h0;
      v_10795 <= 8'h0;
      v_10801 <= 8'h0;
      v_10809 <= 8'h0;
      v_10817 <= 8'h0;
      v_10823 <= 8'h0;
      v_10831 <= 8'h0;
      v_10839 <= 8'h0;
      v_10845 <= 8'h0;
      v_10851 <= 8'h0;
      v_10859 <= 8'h0;
      v_10867 <= 8'h0;
      v_10873 <= 8'h0;
      v_10881 <= 8'h0;
      v_10889 <= 8'h0;
      v_10895 <= 8'h0;
      v_10901 <= 8'h0;
      v_10907 <= 8'h0;
      v_10913 <= 8'h0;
      v_10919 <= 8'h0;
      v_10925 <= 8'h0;
      v_10933 <= 8'h0;
      v_10941 <= 8'h0;
      v_10947 <= 8'h0;
      v_10955 <= 8'h0;
      v_10963 <= 8'h0;
      v_10969 <= 8'h0;
      v_10975 <= 8'h0;
      v_10983 <= 8'h0;
      v_10991 <= 8'h0;
      v_10997 <= 8'h0;
      v_11005 <= 8'h0;
      v_11013 <= 8'h0;
      v_11019 <= 8'h0;
      v_11025 <= 8'h0;
      v_11031 <= 8'h0;
      v_11039 <= 8'h0;
      v_11047 <= 8'h0;
      v_11053 <= 8'h0;
      v_11061 <= 8'h0;
      v_11069 <= 8'h0;
      v_11075 <= 8'h0;
      v_11081 <= 8'h0;
      v_11089 <= 8'h0;
      v_11097 <= 8'h0;
      v_11103 <= 8'h0;
      v_11111 <= 8'h0;
      v_11119 <= 8'h0;
      v_11125 <= 8'h0;
      v_11131 <= 8'h0;
      v_11137 <= 8'h0;
      v_11143 <= 8'h0;
      v_11151 <= 8'h0;
      v_11159 <= 8'h0;
      v_11165 <= 8'h0;
      v_11173 <= 8'h0;
      v_11181 <= 8'h0;
      v_11187 <= 8'h0;
      v_11193 <= 8'h0;
      v_11201 <= 8'h0;
      v_11209 <= 8'h0;
      v_11215 <= 8'h0;
      v_11223 <= 8'h0;
      v_11231 <= 8'h0;
      v_11237 <= 8'h0;
      v_11243 <= 8'h0;
      v_11249 <= 8'h0;
      v_11257 <= 8'h0;
      v_11265 <= 8'h0;
      v_11271 <= 8'h0;
      v_11279 <= 8'h0;
      v_11287 <= 8'h0;
      v_11293 <= 8'h0;
      v_11299 <= 8'h0;
      v_11307 <= 8'h0;
      v_11315 <= 8'h0;
      v_11321 <= 8'h0;
      v_11329 <= 8'h0;
      v_11337 <= 8'h0;
      v_11343 <= 8'h0;
      v_11349 <= 8'h0;
      v_11355 <= 8'h0;
      v_11361 <= 8'h0;
      v_11367 <= 8'h0;
      v_11375 <= 8'h0;
      v_11383 <= 8'h0;
      v_11389 <= 8'h0;
      v_11397 <= 8'h0;
      v_11405 <= 8'h0;
      v_11411 <= 8'h0;
      v_11417 <= 8'h0;
      v_11425 <= 8'h0;
      v_11433 <= 8'h0;
      v_11439 <= 8'h0;
      v_11447 <= 8'h0;
      v_11455 <= 8'h0;
      v_11461 <= 8'h0;
      v_11467 <= 8'h0;
      v_11473 <= 8'h0;
      v_11481 <= 8'h0;
      v_11489 <= 8'h0;
      v_11495 <= 8'h0;
      v_11503 <= 8'h0;
      v_11511 <= 8'h0;
      v_11517 <= 8'h0;
      v_11523 <= 8'h0;
      v_11531 <= 8'h0;
      v_11539 <= 8'h0;
      v_11545 <= 8'h0;
      v_11553 <= 8'h0;
      v_11561 <= 8'h0;
      v_11567 <= 8'h0;
      v_11573 <= 8'h0;
      v_11579 <= 8'h0;
      v_11585 <= 8'h0;
      v_11593 <= 8'h0;
      v_11601 <= 8'h0;
      v_11607 <= 8'h0;
      v_11615 <= 8'h0;
      v_11623 <= 8'h0;
      v_11629 <= 8'h0;
      v_11635 <= 8'h0;
      v_11643 <= 8'h0;
      v_11651 <= 8'h0;
      v_11657 <= 8'h0;
      v_11665 <= 8'h0;
      v_11673 <= 8'h0;
      v_11679 <= 8'h0;
      v_11685 <= 8'h0;
      v_11691 <= 8'h0;
      v_11699 <= 8'h0;
      v_11707 <= 8'h0;
      v_11713 <= 8'h0;
      v_11721 <= 8'h0;
      v_11729 <= 8'h0;
      v_11735 <= 8'h0;
      v_11741 <= 8'h0;
      v_11749 <= 8'h0;
      v_11757 <= 8'h0;
      v_11763 <= 8'h0;
      v_11771 <= 8'h0;
      v_11779 <= 8'h0;
      v_11785 <= 8'h0;
      v_11791 <= 8'h0;
      v_11797 <= 8'h0;
      v_11803 <= 8'h0;
      v_11809 <= 8'h0;
      v_11815 <= 8'h0;
      v_11821 <= 8'h0;
      v_11829 <= 8'h0;
      v_11837 <= 8'h0;
      v_11843 <= 8'h0;
      v_11851 <= 8'h0;
      v_11859 <= 8'h0;
      v_11865 <= 8'h0;
      v_11871 <= 8'h0;
      v_11879 <= 8'h0;
      v_11887 <= 8'h0;
      v_11893 <= 8'h0;
      v_11901 <= 8'h0;
      v_11909 <= 8'h0;
      v_11915 <= 8'h0;
      v_11921 <= 8'h0;
      v_11927 <= 8'h0;
      v_11935 <= 8'h0;
      v_11943 <= 8'h0;
      v_11949 <= 8'h0;
      v_11957 <= 8'h0;
      v_11965 <= 8'h0;
      v_11971 <= 8'h0;
      v_11977 <= 8'h0;
      v_11985 <= 8'h0;
      v_11993 <= 8'h0;
      v_11999 <= 8'h0;
      v_12007 <= 8'h0;
      v_12015 <= 8'h0;
      v_12021 <= 8'h0;
      v_12027 <= 8'h0;
      v_12033 <= 8'h0;
      v_12041 <= 8'h0;
      v_12049 <= 8'h0;
      v_12055 <= 8'h0;
      v_12063 <= 8'h0;
      v_12071 <= 8'h0;
      v_12077 <= 8'h0;
      v_12083 <= 8'h0;
      v_12091 <= 8'h0;
      v_12099 <= 8'h0;
      v_12105 <= 8'h0;
      v_12113 <= 8'h0;
      v_12121 <= 8'h0;
      v_12127 <= 8'h0;
      v_12133 <= 8'h0;
      v_12139 <= 8'h0;
      v_12145 <= 8'h0;
      v_12153 <= 8'h0;
      v_12161 <= 8'h0;
      v_12167 <= 8'h0;
      v_12175 <= 8'h0;
      v_12183 <= 8'h0;
      v_12189 <= 8'h0;
      v_12195 <= 8'h0;
      v_12203 <= 8'h0;
      v_12211 <= 8'h0;
      v_12217 <= 8'h0;
      v_12225 <= 8'h0;
      v_12233 <= 8'h0;
      v_12239 <= 8'h0;
      v_12245 <= 8'h0;
      v_12251 <= 8'h0;
      v_12259 <= 8'h0;
      v_12267 <= 8'h0;
      v_12273 <= 8'h0;
      v_12281 <= 8'h0;
      v_12289 <= 8'h0;
      v_12295 <= 8'h0;
      v_12301 <= 8'h0;
      v_12309 <= 8'h0;
      v_12317 <= 8'h0;
      v_12323 <= 8'h0;
      v_12331 <= 8'h0;
      v_12339 <= 8'h0;
      v_12345 <= 8'h0;
      v_12351 <= 8'h0;
      v_12357 <= 8'h0;
      v_12363 <= 8'h0;
      v_12369 <= 8'h0;
      v_12377 <= 8'h0;
      v_12385 <= 8'h0;
      v_12391 <= 8'h0;
      v_12399 <= 8'h0;
      v_12407 <= 8'h0;
      v_12413 <= 8'h0;
      v_12419 <= 8'h0;
      v_12427 <= 8'h0;
      v_12435 <= 8'h0;
      v_12441 <= 8'h0;
      v_12449 <= 8'h0;
      v_12457 <= 8'h0;
      v_12463 <= 8'h0;
      v_12469 <= 8'h0;
      v_12475 <= 8'h0;
      v_12483 <= 8'h0;
      v_12491 <= 8'h0;
      v_12497 <= 8'h0;
      v_12505 <= 8'h0;
      v_12513 <= 8'h0;
      v_12519 <= 8'h0;
      v_12525 <= 8'h0;
      v_12533 <= 8'h0;
      v_12541 <= 8'h0;
      v_12547 <= 8'h0;
      v_12555 <= 8'h0;
      v_12563 <= 8'h0;
      v_12569 <= 8'h0;
      v_12575 <= 8'h0;
      v_12581 <= 8'h0;
      v_12587 <= 8'h0;
      v_12595 <= 8'h0;
      v_12603 <= 8'h0;
      v_12609 <= 8'h0;
      v_12617 <= 8'h0;
      v_12625 <= 8'h0;
      v_12631 <= 8'h0;
      v_12637 <= 8'h0;
      v_12645 <= 8'h0;
      v_12653 <= 8'h0;
      v_12659 <= 8'h0;
      v_12667 <= 8'h0;
      v_12675 <= 8'h0;
      v_12681 <= 8'h0;
      v_12687 <= 8'h0;
      v_12693 <= 8'h0;
      v_12701 <= 8'h0;
      v_12709 <= 8'h0;
      v_12715 <= 8'h0;
      v_12723 <= 8'h0;
      v_12731 <= 8'h0;
      v_12737 <= 8'h0;
      v_12743 <= 8'h0;
      v_12751 <= 8'h0;
      v_12759 <= 8'h0;
      v_12765 <= 8'h0;
      v_12773 <= 8'h0;
    end else begin
      if (v_2805 == 1) v_2804 <= v_9983;
      if (v_2812 == 1) v_2811 <= v_5381;
      if (v_2819 == 1) v_2818 <= v_3948;
      if (v_2826 == 1) v_2825 <= v_3379;
      if (v_2833 == 1) v_2832 <= v_3098;
      if (v_2840 == 1) v_2839 <= v_2961;
      if (v_2847 == 1) v_2846 <= v_2896;
      if (v_2854 == 1) v_2853 <= v_2867;
      if (v_2871 == 1) v_2870 <= v_2883;
      if (v_2900 == 1) v_2899 <= v_2948;
      if (v_2907 == 1) v_2906 <= v_2920;
      if (v_2924 == 1) v_2923 <= v_2936;
      if (v_2965 == 1) v_2964 <= v_3085;
      if (v_2972 == 1) v_2971 <= v_3021;
      if (v_2979 == 1) v_2978 <= v_2992;
      if (v_2996 == 1) v_2995 <= v_3008;
      if (v_3025 == 1) v_3024 <= v_3073;
      if (v_3032 == 1) v_3031 <= v_3045;
      if (v_3049 == 1) v_3048 <= v_3061;
      if (v_3102 == 1) v_3101 <= v_3366;
      if (v_3109 == 1) v_3108 <= v_3230;
      if (v_3116 == 1) v_3115 <= v_3165;
      if (v_3123 == 1) v_3122 <= v_3136;
      if (v_3140 == 1) v_3139 <= v_3152;
      if (v_3169 == 1) v_3168 <= v_3217;
      if (v_3176 == 1) v_3175 <= v_3189;
      if (v_3193 == 1) v_3192 <= v_3205;
      if (v_3234 == 1) v_3233 <= v_3354;
      if (v_3241 == 1) v_3240 <= v_3290;
      if (v_3248 == 1) v_3247 <= v_3261;
      if (v_3265 == 1) v_3264 <= v_3277;
      if (v_3294 == 1) v_3293 <= v_3342;
      if (v_3301 == 1) v_3300 <= v_3314;
      if (v_3318 == 1) v_3317 <= v_3330;
      if (v_3383 == 1) v_3382 <= v_3935;
      if (v_3390 == 1) v_3389 <= v_3655;
      if (v_3397 == 1) v_3396 <= v_3518;
      if (v_3404 == 1) v_3403 <= v_3453;
      if (v_3411 == 1) v_3410 <= v_3424;
      if (v_3428 == 1) v_3427 <= v_3440;
      if (v_3457 == 1) v_3456 <= v_3505;
      if (v_3464 == 1) v_3463 <= v_3477;
      if (v_3481 == 1) v_3480 <= v_3493;
      if (v_3522 == 1) v_3521 <= v_3642;
      if (v_3529 == 1) v_3528 <= v_3578;
      if (v_3536 == 1) v_3535 <= v_3549;
      if (v_3553 == 1) v_3552 <= v_3565;
      if (v_3582 == 1) v_3581 <= v_3630;
      if (v_3589 == 1) v_3588 <= v_3602;
      if (v_3606 == 1) v_3605 <= v_3618;
      if (v_3659 == 1) v_3658 <= v_3923;
      if (v_3666 == 1) v_3665 <= v_3787;
      if (v_3673 == 1) v_3672 <= v_3722;
      if (v_3680 == 1) v_3679 <= v_3693;
      if (v_3697 == 1) v_3696 <= v_3709;
      if (v_3726 == 1) v_3725 <= v_3774;
      if (v_3733 == 1) v_3732 <= v_3746;
      if (v_3750 == 1) v_3749 <= v_3762;
      if (v_3791 == 1) v_3790 <= v_3911;
      if (v_3798 == 1) v_3797 <= v_3847;
      if (v_3805 == 1) v_3804 <= v_3818;
      if (v_3822 == 1) v_3821 <= v_3834;
      if (v_3851 == 1) v_3850 <= v_3899;
      if (v_3858 == 1) v_3857 <= v_3871;
      if (v_3875 == 1) v_3874 <= v_3887;
      if (v_3952 == 1) v_3951 <= v_5368;
      if (v_3959 == 1) v_3958 <= v_4512;
      if (v_3966 == 1) v_3965 <= v_4231;
      if (v_3973 == 1) v_3972 <= v_4094;
      if (v_3980 == 1) v_3979 <= v_4029;
      if (v_3987 == 1) v_3986 <= v_4000;
      if (v_4004 == 1) v_4003 <= v_4016;
      if (v_4033 == 1) v_4032 <= v_4081;
      if (v_4040 == 1) v_4039 <= v_4053;
      if (v_4057 == 1) v_4056 <= v_4069;
      if (v_4098 == 1) v_4097 <= v_4218;
      if (v_4105 == 1) v_4104 <= v_4154;
      if (v_4112 == 1) v_4111 <= v_4125;
      if (v_4129 == 1) v_4128 <= v_4141;
      if (v_4158 == 1) v_4157 <= v_4206;
      if (v_4165 == 1) v_4164 <= v_4178;
      if (v_4182 == 1) v_4181 <= v_4194;
      if (v_4235 == 1) v_4234 <= v_4499;
      if (v_4242 == 1) v_4241 <= v_4363;
      if (v_4249 == 1) v_4248 <= v_4298;
      if (v_4256 == 1) v_4255 <= v_4269;
      if (v_4273 == 1) v_4272 <= v_4285;
      if (v_4302 == 1) v_4301 <= v_4350;
      if (v_4309 == 1) v_4308 <= v_4322;
      if (v_4326 == 1) v_4325 <= v_4338;
      if (v_4367 == 1) v_4366 <= v_4487;
      if (v_4374 == 1) v_4373 <= v_4423;
      if (v_4381 == 1) v_4380 <= v_4394;
      if (v_4398 == 1) v_4397 <= v_4410;
      if (v_4427 == 1) v_4426 <= v_4475;
      if (v_4434 == 1) v_4433 <= v_4447;
      if (v_4451 == 1) v_4450 <= v_4463;
      if (v_4516 == 1) v_4515 <= v_5356;
      if (v_4523 == 1) v_4522 <= v_4788;
      if (v_4530 == 1) v_4529 <= v_4651;
      if (v_4537 == 1) v_4536 <= v_4586;
      if (v_4544 == 1) v_4543 <= v_4557;
      if (v_4561 == 1) v_4560 <= v_4573;
      if (v_4590 == 1) v_4589 <= v_4638;
      if (v_4597 == 1) v_4596 <= v_4610;
      if (v_4614 == 1) v_4613 <= v_4626;
      if (v_4655 == 1) v_4654 <= v_4775;
      if (v_4662 == 1) v_4661 <= v_4711;
      if (v_4669 == 1) v_4668 <= v_4682;
      if (v_4686 == 1) v_4685 <= v_4698;
      if (v_4715 == 1) v_4714 <= v_4763;
      if (v_4722 == 1) v_4721 <= v_4735;
      if (v_4739 == 1) v_4738 <= v_4751;
      if (v_4792 == 1) v_4791 <= v_5344;
      if (v_4799 == 1) v_4798 <= v_5064;
      if (v_4806 == 1) v_4805 <= v_4927;
      if (v_4813 == 1) v_4812 <= v_4862;
      if (v_4820 == 1) v_4819 <= v_4833;
      if (v_4837 == 1) v_4836 <= v_4849;
      if (v_4866 == 1) v_4865 <= v_4914;
      if (v_4873 == 1) v_4872 <= v_4886;
      if (v_4890 == 1) v_4889 <= v_4902;
      if (v_4931 == 1) v_4930 <= v_5051;
      if (v_4938 == 1) v_4937 <= v_4987;
      if (v_4945 == 1) v_4944 <= v_4958;
      if (v_4962 == 1) v_4961 <= v_4974;
      if (v_4991 == 1) v_4990 <= v_5039;
      if (v_4998 == 1) v_4997 <= v_5011;
      if (v_5015 == 1) v_5014 <= v_5027;
      if (v_5068 == 1) v_5067 <= v_5332;
      if (v_5075 == 1) v_5074 <= v_5196;
      if (v_5082 == 1) v_5081 <= v_5131;
      if (v_5089 == 1) v_5088 <= v_5102;
      if (v_5106 == 1) v_5105 <= v_5118;
      if (v_5135 == 1) v_5134 <= v_5183;
      if (v_5142 == 1) v_5141 <= v_5155;
      if (v_5159 == 1) v_5158 <= v_5171;
      if (v_5200 == 1) v_5199 <= v_5320;
      if (v_5207 == 1) v_5206 <= v_5256;
      if (v_5214 == 1) v_5213 <= v_5227;
      if (v_5231 == 1) v_5230 <= v_5243;
      if (v_5260 == 1) v_5259 <= v_5308;
      if (v_5267 == 1) v_5266 <= v_5280;
      if (v_5284 == 1) v_5283 <= v_5296;
      if (v_5385 == 1) v_5384 <= v_9969;
      if (v_5392 == 1) v_5391 <= v_7673;
      if (v_5399 == 1) v_5398 <= v_6528;
      if (v_5406 == 1) v_5405 <= v_5959;
      if (v_5413 == 1) v_5412 <= v_5678;
      if (v_5420 == 1) v_5419 <= v_5541;
      if (v_5427 == 1) v_5426 <= v_5476;
      if (v_5434 == 1) v_5433 <= v_5447;
      if (v_5451 == 1) v_5450 <= v_5463;
      if (v_5480 == 1) v_5479 <= v_5528;
      if (v_5487 == 1) v_5486 <= v_5500;
      if (v_5504 == 1) v_5503 <= v_5516;
      if (v_5545 == 1) v_5544 <= v_5665;
      if (v_5552 == 1) v_5551 <= v_5601;
      if (v_5559 == 1) v_5558 <= v_5572;
      if (v_5576 == 1) v_5575 <= v_5588;
      if (v_5605 == 1) v_5604 <= v_5653;
      if (v_5612 == 1) v_5611 <= v_5625;
      if (v_5629 == 1) v_5628 <= v_5641;
      if (v_5682 == 1) v_5681 <= v_5946;
      if (v_5689 == 1) v_5688 <= v_5810;
      if (v_5696 == 1) v_5695 <= v_5745;
      if (v_5703 == 1) v_5702 <= v_5716;
      if (v_5720 == 1) v_5719 <= v_5732;
      if (v_5749 == 1) v_5748 <= v_5797;
      if (v_5756 == 1) v_5755 <= v_5769;
      if (v_5773 == 1) v_5772 <= v_5785;
      if (v_5814 == 1) v_5813 <= v_5934;
      if (v_5821 == 1) v_5820 <= v_5870;
      if (v_5828 == 1) v_5827 <= v_5841;
      if (v_5845 == 1) v_5844 <= v_5857;
      if (v_5874 == 1) v_5873 <= v_5922;
      if (v_5881 == 1) v_5880 <= v_5894;
      if (v_5898 == 1) v_5897 <= v_5910;
      if (v_5963 == 1) v_5962 <= v_6515;
      if (v_5970 == 1) v_5969 <= v_6235;
      if (v_5977 == 1) v_5976 <= v_6098;
      if (v_5984 == 1) v_5983 <= v_6033;
      if (v_5991 == 1) v_5990 <= v_6004;
      if (v_6008 == 1) v_6007 <= v_6020;
      if (v_6037 == 1) v_6036 <= v_6085;
      if (v_6044 == 1) v_6043 <= v_6057;
      if (v_6061 == 1) v_6060 <= v_6073;
      if (v_6102 == 1) v_6101 <= v_6222;
      if (v_6109 == 1) v_6108 <= v_6158;
      if (v_6116 == 1) v_6115 <= v_6129;
      if (v_6133 == 1) v_6132 <= v_6145;
      if (v_6162 == 1) v_6161 <= v_6210;
      if (v_6169 == 1) v_6168 <= v_6182;
      if (v_6186 == 1) v_6185 <= v_6198;
      if (v_6239 == 1) v_6238 <= v_6503;
      if (v_6246 == 1) v_6245 <= v_6367;
      if (v_6253 == 1) v_6252 <= v_6302;
      if (v_6260 == 1) v_6259 <= v_6273;
      if (v_6277 == 1) v_6276 <= v_6289;
      if (v_6306 == 1) v_6305 <= v_6354;
      if (v_6313 == 1) v_6312 <= v_6326;
      if (v_6330 == 1) v_6329 <= v_6342;
      if (v_6371 == 1) v_6370 <= v_6491;
      if (v_6378 == 1) v_6377 <= v_6427;
      if (v_6385 == 1) v_6384 <= v_6398;
      if (v_6402 == 1) v_6401 <= v_6414;
      if (v_6431 == 1) v_6430 <= v_6479;
      if (v_6438 == 1) v_6437 <= v_6451;
      if (v_6455 == 1) v_6454 <= v_6467;
      if (v_6532 == 1) v_6531 <= v_7660;
      if (v_6539 == 1) v_6538 <= v_7092;
      if (v_6546 == 1) v_6545 <= v_6811;
      if (v_6553 == 1) v_6552 <= v_6674;
      if (v_6560 == 1) v_6559 <= v_6609;
      if (v_6567 == 1) v_6566 <= v_6580;
      if (v_6584 == 1) v_6583 <= v_6596;
      if (v_6613 == 1) v_6612 <= v_6661;
      if (v_6620 == 1) v_6619 <= v_6633;
      if (v_6637 == 1) v_6636 <= v_6649;
      if (v_6678 == 1) v_6677 <= v_6798;
      if (v_6685 == 1) v_6684 <= v_6734;
      if (v_6692 == 1) v_6691 <= v_6705;
      if (v_6709 == 1) v_6708 <= v_6721;
      if (v_6738 == 1) v_6737 <= v_6786;
      if (v_6745 == 1) v_6744 <= v_6758;
      if (v_6762 == 1) v_6761 <= v_6774;
      if (v_6815 == 1) v_6814 <= v_7079;
      if (v_6822 == 1) v_6821 <= v_6943;
      if (v_6829 == 1) v_6828 <= v_6878;
      if (v_6836 == 1) v_6835 <= v_6849;
      if (v_6853 == 1) v_6852 <= v_6865;
      if (v_6882 == 1) v_6881 <= v_6930;
      if (v_6889 == 1) v_6888 <= v_6902;
      if (v_6906 == 1) v_6905 <= v_6918;
      if (v_6947 == 1) v_6946 <= v_7067;
      if (v_6954 == 1) v_6953 <= v_7003;
      if (v_6961 == 1) v_6960 <= v_6974;
      if (v_6978 == 1) v_6977 <= v_6990;
      if (v_7007 == 1) v_7006 <= v_7055;
      if (v_7014 == 1) v_7013 <= v_7027;
      if (v_7031 == 1) v_7030 <= v_7043;
      if (v_7096 == 1) v_7095 <= v_7648;
      if (v_7103 == 1) v_7102 <= v_7368;
      if (v_7110 == 1) v_7109 <= v_7231;
      if (v_7117 == 1) v_7116 <= v_7166;
      if (v_7124 == 1) v_7123 <= v_7137;
      if (v_7141 == 1) v_7140 <= v_7153;
      if (v_7170 == 1) v_7169 <= v_7218;
      if (v_7177 == 1) v_7176 <= v_7190;
      if (v_7194 == 1) v_7193 <= v_7206;
      if (v_7235 == 1) v_7234 <= v_7355;
      if (v_7242 == 1) v_7241 <= v_7291;
      if (v_7249 == 1) v_7248 <= v_7262;
      if (v_7266 == 1) v_7265 <= v_7278;
      if (v_7295 == 1) v_7294 <= v_7343;
      if (v_7302 == 1) v_7301 <= v_7315;
      if (v_7319 == 1) v_7318 <= v_7331;
      if (v_7372 == 1) v_7371 <= v_7636;
      if (v_7379 == 1) v_7378 <= v_7500;
      if (v_7386 == 1) v_7385 <= v_7435;
      if (v_7393 == 1) v_7392 <= v_7406;
      if (v_7410 == 1) v_7409 <= v_7422;
      if (v_7439 == 1) v_7438 <= v_7487;
      if (v_7446 == 1) v_7445 <= v_7459;
      if (v_7463 == 1) v_7462 <= v_7475;
      if (v_7504 == 1) v_7503 <= v_7624;
      if (v_7511 == 1) v_7510 <= v_7560;
      if (v_7518 == 1) v_7517 <= v_7531;
      if (v_7535 == 1) v_7534 <= v_7547;
      if (v_7564 == 1) v_7563 <= v_7612;
      if (v_7571 == 1) v_7570 <= v_7584;
      if (v_7588 == 1) v_7587 <= v_7600;
      if (v_7677 == 1) v_7676 <= v_9957;
      if (v_7684 == 1) v_7683 <= v_8813;
      if (v_7691 == 1) v_7690 <= v_8244;
      if (v_7698 == 1) v_7697 <= v_7963;
      if (v_7705 == 1) v_7704 <= v_7826;
      if (v_7712 == 1) v_7711 <= v_7761;
      if (v_7719 == 1) v_7718 <= v_7732;
      if (v_7736 == 1) v_7735 <= v_7748;
      if (v_7765 == 1) v_7764 <= v_7813;
      if (v_7772 == 1) v_7771 <= v_7785;
      if (v_7789 == 1) v_7788 <= v_7801;
      if (v_7830 == 1) v_7829 <= v_7950;
      if (v_7837 == 1) v_7836 <= v_7886;
      if (v_7844 == 1) v_7843 <= v_7857;
      if (v_7861 == 1) v_7860 <= v_7873;
      if (v_7890 == 1) v_7889 <= v_7938;
      if (v_7897 == 1) v_7896 <= v_7910;
      if (v_7914 == 1) v_7913 <= v_7926;
      if (v_7967 == 1) v_7966 <= v_8231;
      if (v_7974 == 1) v_7973 <= v_8095;
      if (v_7981 == 1) v_7980 <= v_8030;
      if (v_7988 == 1) v_7987 <= v_8001;
      if (v_8005 == 1) v_8004 <= v_8017;
      if (v_8034 == 1) v_8033 <= v_8082;
      if (v_8041 == 1) v_8040 <= v_8054;
      if (v_8058 == 1) v_8057 <= v_8070;
      if (v_8099 == 1) v_8098 <= v_8219;
      if (v_8106 == 1) v_8105 <= v_8155;
      if (v_8113 == 1) v_8112 <= v_8126;
      if (v_8130 == 1) v_8129 <= v_8142;
      if (v_8159 == 1) v_8158 <= v_8207;
      if (v_8166 == 1) v_8165 <= v_8179;
      if (v_8183 == 1) v_8182 <= v_8195;
      if (v_8248 == 1) v_8247 <= v_8800;
      if (v_8255 == 1) v_8254 <= v_8520;
      if (v_8262 == 1) v_8261 <= v_8383;
      if (v_8269 == 1) v_8268 <= v_8318;
      if (v_8276 == 1) v_8275 <= v_8289;
      if (v_8293 == 1) v_8292 <= v_8305;
      if (v_8322 == 1) v_8321 <= v_8370;
      if (v_8329 == 1) v_8328 <= v_8342;
      if (v_8346 == 1) v_8345 <= v_8358;
      if (v_8387 == 1) v_8386 <= v_8507;
      if (v_8394 == 1) v_8393 <= v_8443;
      if (v_8401 == 1) v_8400 <= v_8414;
      if (v_8418 == 1) v_8417 <= v_8430;
      if (v_8447 == 1) v_8446 <= v_8495;
      if (v_8454 == 1) v_8453 <= v_8467;
      if (v_8471 == 1) v_8470 <= v_8483;
      if (v_8524 == 1) v_8523 <= v_8788;
      if (v_8531 == 1) v_8530 <= v_8652;
      if (v_8538 == 1) v_8537 <= v_8587;
      if (v_8545 == 1) v_8544 <= v_8558;
      if (v_8562 == 1) v_8561 <= v_8574;
      if (v_8591 == 1) v_8590 <= v_8639;
      if (v_8598 == 1) v_8597 <= v_8611;
      if (v_8615 == 1) v_8614 <= v_8627;
      if (v_8656 == 1) v_8655 <= v_8776;
      if (v_8663 == 1) v_8662 <= v_8712;
      if (v_8670 == 1) v_8669 <= v_8683;
      if (v_8687 == 1) v_8686 <= v_8699;
      if (v_8716 == 1) v_8715 <= v_8764;
      if (v_8723 == 1) v_8722 <= v_8736;
      if (v_8740 == 1) v_8739 <= v_8752;
      if (v_8817 == 1) v_8816 <= v_9945;
      if (v_8824 == 1) v_8823 <= v_9377;
      if (v_8831 == 1) v_8830 <= v_9096;
      if (v_8838 == 1) v_8837 <= v_8959;
      if (v_8845 == 1) v_8844 <= v_8894;
      if (v_8852 == 1) v_8851 <= v_8865;
      if (v_8869 == 1) v_8868 <= v_8881;
      if (v_8898 == 1) v_8897 <= v_8946;
      if (v_8905 == 1) v_8904 <= v_8918;
      if (v_8922 == 1) v_8921 <= v_8934;
      if (v_8963 == 1) v_8962 <= v_9083;
      if (v_8970 == 1) v_8969 <= v_9019;
      if (v_8977 == 1) v_8976 <= v_8990;
      if (v_8994 == 1) v_8993 <= v_9006;
      if (v_9023 == 1) v_9022 <= v_9071;
      if (v_9030 == 1) v_9029 <= v_9043;
      if (v_9047 == 1) v_9046 <= v_9059;
      if (v_9100 == 1) v_9099 <= v_9364;
      if (v_9107 == 1) v_9106 <= v_9228;
      if (v_9114 == 1) v_9113 <= v_9163;
      if (v_9121 == 1) v_9120 <= v_9134;
      if (v_9138 == 1) v_9137 <= v_9150;
      if (v_9167 == 1) v_9166 <= v_9215;
      if (v_9174 == 1) v_9173 <= v_9187;
      if (v_9191 == 1) v_9190 <= v_9203;
      if (v_9232 == 1) v_9231 <= v_9352;
      if (v_9239 == 1) v_9238 <= v_9288;
      if (v_9246 == 1) v_9245 <= v_9259;
      if (v_9263 == 1) v_9262 <= v_9275;
      if (v_9292 == 1) v_9291 <= v_9340;
      if (v_9299 == 1) v_9298 <= v_9312;
      if (v_9316 == 1) v_9315 <= v_9328;
      if (v_9381 == 1) v_9380 <= v_9933;
      if (v_9388 == 1) v_9387 <= v_9653;
      if (v_9395 == 1) v_9394 <= v_9516;
      if (v_9402 == 1) v_9401 <= v_9451;
      if (v_9409 == 1) v_9408 <= v_9422;
      if (v_9426 == 1) v_9425 <= v_9438;
      if (v_9455 == 1) v_9454 <= v_9503;
      if (v_9462 == 1) v_9461 <= v_9475;
      if (v_9479 == 1) v_9478 <= v_9491;
      if (v_9520 == 1) v_9519 <= v_9640;
      if (v_9527 == 1) v_9526 <= v_9576;
      if (v_9534 == 1) v_9533 <= v_9547;
      if (v_9551 == 1) v_9550 <= v_9563;
      if (v_9580 == 1) v_9579 <= v_9628;
      if (v_9587 == 1) v_9586 <= v_9600;
      if (v_9604 == 1) v_9603 <= v_9616;
      if (v_9657 == 1) v_9656 <= v_9921;
      if (v_9664 == 1) v_9663 <= v_9785;
      if (v_9671 == 1) v_9670 <= v_9720;
      if (v_9678 == 1) v_9677 <= v_9691;
      if (v_9695 == 1) v_9694 <= v_9707;
      if (v_9724 == 1) v_9723 <= v_9772;
      if (v_9731 == 1) v_9730 <= v_9744;
      if (v_9748 == 1) v_9747 <= v_9760;
      if (v_9789 == 1) v_9788 <= v_9909;
      if (v_9796 == 1) v_9795 <= v_9845;
      if (v_9803 == 1) v_9802 <= v_9816;
      if (v_9820 == 1) v_9819 <= v_9832;
      if (v_9849 == 1) v_9848 <= v_9897;
      if (v_9856 == 1) v_9855 <= v_9869;
      if (v_9873 == 1) v_9872 <= v_9885;
      if (v_2806 == 1) v_9987 <= v_9988;
      if (v_5386 == 1) v_9993 <= v_9994;
      if (v_7678 == 1) v_9999 <= v_10000;
      if (v_8818 == 1) v_10005 <= v_10006;
      if (v_9382 == 1) v_10011 <= v_10012;
      if (v_9658 == 1) v_10017 <= v_10018;
      if (v_9790 == 1) v_10023 <= v_10024;
      if (v_9850 == 1) v_10029 <= v_10030;
      if (v_9874 == 1) v_10035 <= v_10036;
      if (v_9857 == 1) v_10043 <= v_10044;
      if (v_9797 == 1) v_10051 <= v_10052;
      if (v_9821 == 1) v_10057 <= v_10058;
      if (v_9804 == 1) v_10065 <= v_10066;
      if (v_9665 == 1) v_10073 <= v_10074;
      if (v_9725 == 1) v_10079 <= v_10080;
      if (v_9749 == 1) v_10085 <= v_10086;
      if (v_9732 == 1) v_10093 <= v_10094;
      if (v_9672 == 1) v_10101 <= v_10102;
      if (v_9696 == 1) v_10107 <= v_10108;
      if (v_9679 == 1) v_10115 <= v_10116;
      if (v_9389 == 1) v_10123 <= v_10124;
      if (v_9521 == 1) v_10129 <= v_10130;
      if (v_9581 == 1) v_10135 <= v_10136;
      if (v_9605 == 1) v_10141 <= v_10142;
      if (v_9588 == 1) v_10149 <= v_10150;
      if (v_9528 == 1) v_10157 <= v_10158;
      if (v_9552 == 1) v_10163 <= v_10164;
      if (v_9535 == 1) v_10171 <= v_10172;
      if (v_9396 == 1) v_10179 <= v_10180;
      if (v_9456 == 1) v_10185 <= v_10186;
      if (v_9480 == 1) v_10191 <= v_10192;
      if (v_9463 == 1) v_10199 <= v_10200;
      if (v_9403 == 1) v_10207 <= v_10208;
      if (v_9427 == 1) v_10213 <= v_10214;
      if (v_9410 == 1) v_10221 <= v_10222;
      if (v_8825 == 1) v_10229 <= v_10230;
      if (v_9101 == 1) v_10235 <= v_10236;
      if (v_9233 == 1) v_10241 <= v_10242;
      if (v_9293 == 1) v_10247 <= v_10248;
      if (v_9317 == 1) v_10253 <= v_10254;
      if (v_9300 == 1) v_10261 <= v_10262;
      if (v_9240 == 1) v_10269 <= v_10270;
      if (v_9264 == 1) v_10275 <= v_10276;
      if (v_9247 == 1) v_10283 <= v_10284;
      if (v_9108 == 1) v_10291 <= v_10292;
      if (v_9168 == 1) v_10297 <= v_10298;
      if (v_9192 == 1) v_10303 <= v_10304;
      if (v_9175 == 1) v_10311 <= v_10312;
      if (v_9115 == 1) v_10319 <= v_10320;
      if (v_9139 == 1) v_10325 <= v_10326;
      if (v_9122 == 1) v_10333 <= v_10334;
      if (v_8832 == 1) v_10341 <= v_10342;
      if (v_8964 == 1) v_10347 <= v_10348;
      if (v_9024 == 1) v_10353 <= v_10354;
      if (v_9048 == 1) v_10359 <= v_10360;
      if (v_9031 == 1) v_10367 <= v_10368;
      if (v_8971 == 1) v_10375 <= v_10376;
      if (v_8995 == 1) v_10381 <= v_10382;
      if (v_8978 == 1) v_10389 <= v_10390;
      if (v_8839 == 1) v_10397 <= v_10398;
      if (v_8899 == 1) v_10403 <= v_10404;
      if (v_8923 == 1) v_10409 <= v_10410;
      if (v_8906 == 1) v_10417 <= v_10418;
      if (v_8846 == 1) v_10425 <= v_10426;
      if (v_8870 == 1) v_10431 <= v_10432;
      if (v_8853 == 1) v_10439 <= v_10440;
      if (v_7685 == 1) v_10447 <= v_10448;
      if (v_8249 == 1) v_10453 <= v_10454;
      if (v_8525 == 1) v_10459 <= v_10460;
      if (v_8657 == 1) v_10465 <= v_10466;
      if (v_8717 == 1) v_10471 <= v_10472;
      if (v_8741 == 1) v_10477 <= v_10478;
      if (v_8724 == 1) v_10485 <= v_10486;
      if (v_8664 == 1) v_10493 <= v_10494;
      if (v_8688 == 1) v_10499 <= v_10500;
      if (v_8671 == 1) v_10507 <= v_10508;
      if (v_8532 == 1) v_10515 <= v_10516;
      if (v_8592 == 1) v_10521 <= v_10522;
      if (v_8616 == 1) v_10527 <= v_10528;
      if (v_8599 == 1) v_10535 <= v_10536;
      if (v_8539 == 1) v_10543 <= v_10544;
      if (v_8563 == 1) v_10549 <= v_10550;
      if (v_8546 == 1) v_10557 <= v_10558;
      if (v_8256 == 1) v_10565 <= v_10566;
      if (v_8388 == 1) v_10571 <= v_10572;
      if (v_8448 == 1) v_10577 <= v_10578;
      if (v_8472 == 1) v_10583 <= v_10584;
      if (v_8455 == 1) v_10591 <= v_10592;
      if (v_8395 == 1) v_10599 <= v_10600;
      if (v_8419 == 1) v_10605 <= v_10606;
      if (v_8402 == 1) v_10613 <= v_10614;
      if (v_8263 == 1) v_10621 <= v_10622;
      if (v_8323 == 1) v_10627 <= v_10628;
      if (v_8347 == 1) v_10633 <= v_10634;
      if (v_8330 == 1) v_10641 <= v_10642;
      if (v_8270 == 1) v_10649 <= v_10650;
      if (v_8294 == 1) v_10655 <= v_10656;
      if (v_8277 == 1) v_10663 <= v_10664;
      if (v_7692 == 1) v_10671 <= v_10672;
      if (v_7968 == 1) v_10677 <= v_10678;
      if (v_8100 == 1) v_10683 <= v_10684;
      if (v_8160 == 1) v_10689 <= v_10690;
      if (v_8184 == 1) v_10695 <= v_10696;
      if (v_8167 == 1) v_10703 <= v_10704;
      if (v_8107 == 1) v_10711 <= v_10712;
      if (v_8131 == 1) v_10717 <= v_10718;
      if (v_8114 == 1) v_10725 <= v_10726;
      if (v_7975 == 1) v_10733 <= v_10734;
      if (v_8035 == 1) v_10739 <= v_10740;
      if (v_8059 == 1) v_10745 <= v_10746;
      if (v_8042 == 1) v_10753 <= v_10754;
      if (v_7982 == 1) v_10761 <= v_10762;
      if (v_8006 == 1) v_10767 <= v_10768;
      if (v_7989 == 1) v_10775 <= v_10776;
      if (v_7699 == 1) v_10783 <= v_10784;
      if (v_7831 == 1) v_10789 <= v_10790;
      if (v_7891 == 1) v_10795 <= v_10796;
      if (v_7915 == 1) v_10801 <= v_10802;
      if (v_7898 == 1) v_10809 <= v_10810;
      if (v_7838 == 1) v_10817 <= v_10818;
      if (v_7862 == 1) v_10823 <= v_10824;
      if (v_7845 == 1) v_10831 <= v_10832;
      if (v_7706 == 1) v_10839 <= v_10840;
      if (v_7766 == 1) v_10845 <= v_10846;
      if (v_7790 == 1) v_10851 <= v_10852;
      if (v_7773 == 1) v_10859 <= v_10860;
      if (v_7713 == 1) v_10867 <= v_10868;
      if (v_7737 == 1) v_10873 <= v_10874;
      if (v_7720 == 1) v_10881 <= v_10882;
      if (v_5393 == 1) v_10889 <= v_10890;
      if (v_6533 == 1) v_10895 <= v_10896;
      if (v_7097 == 1) v_10901 <= v_10902;
      if (v_7373 == 1) v_10907 <= v_10908;
      if (v_7505 == 1) v_10913 <= v_10914;
      if (v_7565 == 1) v_10919 <= v_10920;
      if (v_7589 == 1) v_10925 <= v_10926;
      if (v_7572 == 1) v_10933 <= v_10934;
      if (v_7512 == 1) v_10941 <= v_10942;
      if (v_7536 == 1) v_10947 <= v_10948;
      if (v_7519 == 1) v_10955 <= v_10956;
      if (v_7380 == 1) v_10963 <= v_10964;
      if (v_7440 == 1) v_10969 <= v_10970;
      if (v_7464 == 1) v_10975 <= v_10976;
      if (v_7447 == 1) v_10983 <= v_10984;
      if (v_7387 == 1) v_10991 <= v_10992;
      if (v_7411 == 1) v_10997 <= v_10998;
      if (v_7394 == 1) v_11005 <= v_11006;
      if (v_7104 == 1) v_11013 <= v_11014;
      if (v_7236 == 1) v_11019 <= v_11020;
      if (v_7296 == 1) v_11025 <= v_11026;
      if (v_7320 == 1) v_11031 <= v_11032;
      if (v_7303 == 1) v_11039 <= v_11040;
      if (v_7243 == 1) v_11047 <= v_11048;
      if (v_7267 == 1) v_11053 <= v_11054;
      if (v_7250 == 1) v_11061 <= v_11062;
      if (v_7111 == 1) v_11069 <= v_11070;
      if (v_7171 == 1) v_11075 <= v_11076;
      if (v_7195 == 1) v_11081 <= v_11082;
      if (v_7178 == 1) v_11089 <= v_11090;
      if (v_7118 == 1) v_11097 <= v_11098;
      if (v_7142 == 1) v_11103 <= v_11104;
      if (v_7125 == 1) v_11111 <= v_11112;
      if (v_6540 == 1) v_11119 <= v_11120;
      if (v_6816 == 1) v_11125 <= v_11126;
      if (v_6948 == 1) v_11131 <= v_11132;
      if (v_7008 == 1) v_11137 <= v_11138;
      if (v_7032 == 1) v_11143 <= v_11144;
      if (v_7015 == 1) v_11151 <= v_11152;
      if (v_6955 == 1) v_11159 <= v_11160;
      if (v_6979 == 1) v_11165 <= v_11166;
      if (v_6962 == 1) v_11173 <= v_11174;
      if (v_6823 == 1) v_11181 <= v_11182;
      if (v_6883 == 1) v_11187 <= v_11188;
      if (v_6907 == 1) v_11193 <= v_11194;
      if (v_6890 == 1) v_11201 <= v_11202;
      if (v_6830 == 1) v_11209 <= v_11210;
      if (v_6854 == 1) v_11215 <= v_11216;
      if (v_6837 == 1) v_11223 <= v_11224;
      if (v_6547 == 1) v_11231 <= v_11232;
      if (v_6679 == 1) v_11237 <= v_11238;
      if (v_6739 == 1) v_11243 <= v_11244;
      if (v_6763 == 1) v_11249 <= v_11250;
      if (v_6746 == 1) v_11257 <= v_11258;
      if (v_6686 == 1) v_11265 <= v_11266;
      if (v_6710 == 1) v_11271 <= v_11272;
      if (v_6693 == 1) v_11279 <= v_11280;
      if (v_6554 == 1) v_11287 <= v_11288;
      if (v_6614 == 1) v_11293 <= v_11294;
      if (v_6638 == 1) v_11299 <= v_11300;
      if (v_6621 == 1) v_11307 <= v_11308;
      if (v_6561 == 1) v_11315 <= v_11316;
      if (v_6585 == 1) v_11321 <= v_11322;
      if (v_6568 == 1) v_11329 <= v_11330;
      if (v_5400 == 1) v_11337 <= v_11338;
      if (v_5964 == 1) v_11343 <= v_11344;
      if (v_6240 == 1) v_11349 <= v_11350;
      if (v_6372 == 1) v_11355 <= v_11356;
      if (v_6432 == 1) v_11361 <= v_11362;
      if (v_6456 == 1) v_11367 <= v_11368;
      if (v_6439 == 1) v_11375 <= v_11376;
      if (v_6379 == 1) v_11383 <= v_11384;
      if (v_6403 == 1) v_11389 <= v_11390;
      if (v_6386 == 1) v_11397 <= v_11398;
      if (v_6247 == 1) v_11405 <= v_11406;
      if (v_6307 == 1) v_11411 <= v_11412;
      if (v_6331 == 1) v_11417 <= v_11418;
      if (v_6314 == 1) v_11425 <= v_11426;
      if (v_6254 == 1) v_11433 <= v_11434;
      if (v_6278 == 1) v_11439 <= v_11440;
      if (v_6261 == 1) v_11447 <= v_11448;
      if (v_5971 == 1) v_11455 <= v_11456;
      if (v_6103 == 1) v_11461 <= v_11462;
      if (v_6163 == 1) v_11467 <= v_11468;
      if (v_6187 == 1) v_11473 <= v_11474;
      if (v_6170 == 1) v_11481 <= v_11482;
      if (v_6110 == 1) v_11489 <= v_11490;
      if (v_6134 == 1) v_11495 <= v_11496;
      if (v_6117 == 1) v_11503 <= v_11504;
      if (v_5978 == 1) v_11511 <= v_11512;
      if (v_6038 == 1) v_11517 <= v_11518;
      if (v_6062 == 1) v_11523 <= v_11524;
      if (v_6045 == 1) v_11531 <= v_11532;
      if (v_5985 == 1) v_11539 <= v_11540;
      if (v_6009 == 1) v_11545 <= v_11546;
      if (v_5992 == 1) v_11553 <= v_11554;
      if (v_5407 == 1) v_11561 <= v_11562;
      if (v_5683 == 1) v_11567 <= v_11568;
      if (v_5815 == 1) v_11573 <= v_11574;
      if (v_5875 == 1) v_11579 <= v_11580;
      if (v_5899 == 1) v_11585 <= v_11586;
      if (v_5882 == 1) v_11593 <= v_11594;
      if (v_5822 == 1) v_11601 <= v_11602;
      if (v_5846 == 1) v_11607 <= v_11608;
      if (v_5829 == 1) v_11615 <= v_11616;
      if (v_5690 == 1) v_11623 <= v_11624;
      if (v_5750 == 1) v_11629 <= v_11630;
      if (v_5774 == 1) v_11635 <= v_11636;
      if (v_5757 == 1) v_11643 <= v_11644;
      if (v_5697 == 1) v_11651 <= v_11652;
      if (v_5721 == 1) v_11657 <= v_11658;
      if (v_5704 == 1) v_11665 <= v_11666;
      if (v_5414 == 1) v_11673 <= v_11674;
      if (v_5546 == 1) v_11679 <= v_11680;
      if (v_5606 == 1) v_11685 <= v_11686;
      if (v_5630 == 1) v_11691 <= v_11692;
      if (v_5613 == 1) v_11699 <= v_11700;
      if (v_5553 == 1) v_11707 <= v_11708;
      if (v_5577 == 1) v_11713 <= v_11714;
      if (v_5560 == 1) v_11721 <= v_11722;
      if (v_5421 == 1) v_11729 <= v_11730;
      if (v_5481 == 1) v_11735 <= v_11736;
      if (v_5505 == 1) v_11741 <= v_11742;
      if (v_5488 == 1) v_11749 <= v_11750;
      if (v_5428 == 1) v_11757 <= v_11758;
      if (v_5452 == 1) v_11763 <= v_11764;
      if (v_5435 == 1) v_11771 <= v_11772;
      if (v_2813 == 1) v_11779 <= v_11780;
      if (v_3953 == 1) v_11785 <= v_11786;
      if (v_4517 == 1) v_11791 <= v_11792;
      if (v_4793 == 1) v_11797 <= v_11798;
      if (v_5069 == 1) v_11803 <= v_11804;
      if (v_5201 == 1) v_11809 <= v_11810;
      if (v_5261 == 1) v_11815 <= v_11816;
      if (v_5285 == 1) v_11821 <= v_11822;
      if (v_5268 == 1) v_11829 <= v_11830;
      if (v_5208 == 1) v_11837 <= v_11838;
      if (v_5232 == 1) v_11843 <= v_11844;
      if (v_5215 == 1) v_11851 <= v_11852;
      if (v_5076 == 1) v_11859 <= v_11860;
      if (v_5136 == 1) v_11865 <= v_11866;
      if (v_5160 == 1) v_11871 <= v_11872;
      if (v_5143 == 1) v_11879 <= v_11880;
      if (v_5083 == 1) v_11887 <= v_11888;
      if (v_5107 == 1) v_11893 <= v_11894;
      if (v_5090 == 1) v_11901 <= v_11902;
      if (v_4800 == 1) v_11909 <= v_11910;
      if (v_4932 == 1) v_11915 <= v_11916;
      if (v_4992 == 1) v_11921 <= v_11922;
      if (v_5016 == 1) v_11927 <= v_11928;
      if (v_4999 == 1) v_11935 <= v_11936;
      if (v_4939 == 1) v_11943 <= v_11944;
      if (v_4963 == 1) v_11949 <= v_11950;
      if (v_4946 == 1) v_11957 <= v_11958;
      if (v_4807 == 1) v_11965 <= v_11966;
      if (v_4867 == 1) v_11971 <= v_11972;
      if (v_4891 == 1) v_11977 <= v_11978;
      if (v_4874 == 1) v_11985 <= v_11986;
      if (v_4814 == 1) v_11993 <= v_11994;
      if (v_4838 == 1) v_11999 <= v_12000;
      if (v_4821 == 1) v_12007 <= v_12008;
      if (v_4524 == 1) v_12015 <= v_12016;
      if (v_4656 == 1) v_12021 <= v_12022;
      if (v_4716 == 1) v_12027 <= v_12028;
      if (v_4740 == 1) v_12033 <= v_12034;
      if (v_4723 == 1) v_12041 <= v_12042;
      if (v_4663 == 1) v_12049 <= v_12050;
      if (v_4687 == 1) v_12055 <= v_12056;
      if (v_4670 == 1) v_12063 <= v_12064;
      if (v_4531 == 1) v_12071 <= v_12072;
      if (v_4591 == 1) v_12077 <= v_12078;
      if (v_4615 == 1) v_12083 <= v_12084;
      if (v_4598 == 1) v_12091 <= v_12092;
      if (v_4538 == 1) v_12099 <= v_12100;
      if (v_4562 == 1) v_12105 <= v_12106;
      if (v_4545 == 1) v_12113 <= v_12114;
      if (v_3960 == 1) v_12121 <= v_12122;
      if (v_4236 == 1) v_12127 <= v_12128;
      if (v_4368 == 1) v_12133 <= v_12134;
      if (v_4428 == 1) v_12139 <= v_12140;
      if (v_4452 == 1) v_12145 <= v_12146;
      if (v_4435 == 1) v_12153 <= v_12154;
      if (v_4375 == 1) v_12161 <= v_12162;
      if (v_4399 == 1) v_12167 <= v_12168;
      if (v_4382 == 1) v_12175 <= v_12176;
      if (v_4243 == 1) v_12183 <= v_12184;
      if (v_4303 == 1) v_12189 <= v_12190;
      if (v_4327 == 1) v_12195 <= v_12196;
      if (v_4310 == 1) v_12203 <= v_12204;
      if (v_4250 == 1) v_12211 <= v_12212;
      if (v_4274 == 1) v_12217 <= v_12218;
      if (v_4257 == 1) v_12225 <= v_12226;
      if (v_3967 == 1) v_12233 <= v_12234;
      if (v_4099 == 1) v_12239 <= v_12240;
      if (v_4159 == 1) v_12245 <= v_12246;
      if (v_4183 == 1) v_12251 <= v_12252;
      if (v_4166 == 1) v_12259 <= v_12260;
      if (v_4106 == 1) v_12267 <= v_12268;
      if (v_4130 == 1) v_12273 <= v_12274;
      if (v_4113 == 1) v_12281 <= v_12282;
      if (v_3974 == 1) v_12289 <= v_12290;
      if (v_4034 == 1) v_12295 <= v_12296;
      if (v_4058 == 1) v_12301 <= v_12302;
      if (v_4041 == 1) v_12309 <= v_12310;
      if (v_3981 == 1) v_12317 <= v_12318;
      if (v_4005 == 1) v_12323 <= v_12324;
      if (v_3988 == 1) v_12331 <= v_12332;
      if (v_2820 == 1) v_12339 <= v_12340;
      if (v_3384 == 1) v_12345 <= v_12346;
      if (v_3660 == 1) v_12351 <= v_12352;
      if (v_3792 == 1) v_12357 <= v_12358;
      if (v_3852 == 1) v_12363 <= v_12364;
      if (v_3876 == 1) v_12369 <= v_12370;
      if (v_3859 == 1) v_12377 <= v_12378;
      if (v_3799 == 1) v_12385 <= v_12386;
      if (v_3823 == 1) v_12391 <= v_12392;
      if (v_3806 == 1) v_12399 <= v_12400;
      if (v_3667 == 1) v_12407 <= v_12408;
      if (v_3727 == 1) v_12413 <= v_12414;
      if (v_3751 == 1) v_12419 <= v_12420;
      if (v_3734 == 1) v_12427 <= v_12428;
      if (v_3674 == 1) v_12435 <= v_12436;
      if (v_3698 == 1) v_12441 <= v_12442;
      if (v_3681 == 1) v_12449 <= v_12450;
      if (v_3391 == 1) v_12457 <= v_12458;
      if (v_3523 == 1) v_12463 <= v_12464;
      if (v_3583 == 1) v_12469 <= v_12470;
      if (v_3607 == 1) v_12475 <= v_12476;
      if (v_3590 == 1) v_12483 <= v_12484;
      if (v_3530 == 1) v_12491 <= v_12492;
      if (v_3554 == 1) v_12497 <= v_12498;
      if (v_3537 == 1) v_12505 <= v_12506;
      if (v_3398 == 1) v_12513 <= v_12514;
      if (v_3458 == 1) v_12519 <= v_12520;
      if (v_3482 == 1) v_12525 <= v_12526;
      if (v_3465 == 1) v_12533 <= v_12534;
      if (v_3405 == 1) v_12541 <= v_12542;
      if (v_3429 == 1) v_12547 <= v_12548;
      if (v_3412 == 1) v_12555 <= v_12556;
      if (v_2827 == 1) v_12563 <= v_12564;
      if (v_3103 == 1) v_12569 <= v_12570;
      if (v_3235 == 1) v_12575 <= v_12576;
      if (v_3295 == 1) v_12581 <= v_12582;
      if (v_3319 == 1) v_12587 <= v_12588;
      if (v_3302 == 1) v_12595 <= v_12596;
      if (v_3242 == 1) v_12603 <= v_12604;
      if (v_3266 == 1) v_12609 <= v_12610;
      if (v_3249 == 1) v_12617 <= v_12618;
      if (v_3110 == 1) v_12625 <= v_12626;
      if (v_3170 == 1) v_12631 <= v_12632;
      if (v_3194 == 1) v_12637 <= v_12638;
      if (v_3177 == 1) v_12645 <= v_12646;
      if (v_3117 == 1) v_12653 <= v_12654;
      if (v_3141 == 1) v_12659 <= v_12660;
      if (v_3124 == 1) v_12667 <= v_12668;
      if (v_2834 == 1) v_12675 <= v_12676;
      if (v_2966 == 1) v_12681 <= v_12682;
      if (v_3026 == 1) v_12687 <= v_12688;
      if (v_3050 == 1) v_12693 <= v_12694;
      if (v_3033 == 1) v_12701 <= v_12702;
      if (v_2973 == 1) v_12709 <= v_12710;
      if (v_2997 == 1) v_12715 <= v_12716;
      if (v_2980 == 1) v_12723 <= v_12724;
      if (v_2841 == 1) v_12731 <= v_12732;
      if (v_2901 == 1) v_12737 <= v_12738;
      if (v_2925 == 1) v_12743 <= v_12744;
      if (v_2908 == 1) v_12751 <= v_12752;
      if (v_2848 == 1) v_12759 <= v_12760;
      if (v_2872 == 1) v_12765 <= v_12766;
      if (v_2855 == 1) v_12773 <= v_12774;
    end
  end
endmodule